magic
tech sky130A
magscale 1 2
timestamp 1653512069
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118720
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9678 119200 9734 120000
rect 11150 119200 11206 120000
rect 12622 119200 12678 120000
rect 14094 119200 14150 120000
rect 15566 119200 15622 120000
rect 17038 119200 17094 120000
rect 18602 119200 18658 120000
rect 20074 119200 20130 120000
rect 21546 119200 21602 120000
rect 23018 119200 23074 120000
rect 24490 119200 24546 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30470 119200 30526 120000
rect 31942 119200 31998 120000
rect 33414 119200 33470 120000
rect 34886 119200 34942 120000
rect 36450 119200 36506 120000
rect 37922 119200 37978 120000
rect 39394 119200 39450 120000
rect 40866 119200 40922 120000
rect 42338 119200 42394 120000
rect 43902 119200 43958 120000
rect 45374 119200 45430 120000
rect 46846 119200 46902 120000
rect 48318 119200 48374 120000
rect 49790 119200 49846 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54298 119200 54354 120000
rect 55770 119200 55826 120000
rect 57242 119200 57298 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63222 119200 63278 120000
rect 64694 119200 64750 120000
rect 66166 119200 66222 120000
rect 67638 119200 67694 120000
rect 69110 119200 69166 120000
rect 70674 119200 70730 120000
rect 72146 119200 72202 120000
rect 73618 119200 73674 120000
rect 75090 119200 75146 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79598 119200 79654 120000
rect 81070 119200 81126 120000
rect 82542 119200 82598 120000
rect 84014 119200 84070 120000
rect 85486 119200 85542 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89994 119200 90050 120000
rect 91466 119200 91522 120000
rect 92938 119200 92994 120000
rect 94410 119200 94466 120000
rect 95974 119200 96030 120000
rect 97446 119200 97502 120000
rect 98918 119200 98974 120000
rect 100390 119200 100446 120000
rect 101862 119200 101918 120000
rect 103334 119200 103390 120000
rect 104898 119200 104954 120000
rect 106370 119200 106426 120000
rect 107842 119200 107898 120000
rect 109314 119200 109370 120000
rect 110786 119200 110842 120000
rect 112350 119200 112406 120000
rect 113822 119200 113878 120000
rect 115294 119200 115350 120000
rect 116766 119200 116822 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122746 119200 122802 120000
rect 124218 119200 124274 120000
rect 125690 119200 125746 120000
rect 127162 119200 127218 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131670 119200 131726 120000
rect 133142 119200 133198 120000
rect 134614 119200 134670 120000
rect 136086 119200 136142 120000
rect 137558 119200 137614 120000
rect 139122 119200 139178 120000
rect 140594 119200 140650 120000
rect 142066 119200 142122 120000
rect 143538 119200 143594 120000
rect 145010 119200 145066 120000
rect 146574 119200 146630 120000
rect 148046 119200 148102 120000
rect 149518 119200 149574 120000
rect 150990 119200 151046 120000
rect 152462 119200 152518 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 156970 119200 157026 120000
rect 158442 119200 158498 120000
rect 159914 119200 159970 120000
rect 161386 119200 161442 120000
rect 162858 119200 162914 120000
rect 164422 119200 164478 120000
rect 165894 119200 165950 120000
rect 167366 119200 167422 120000
rect 168838 119200 168894 120000
rect 170310 119200 170366 120000
rect 171782 119200 171838 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39854 0 39910 800
rect 40222 0 40278 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61842 0 61898 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65154 0 65210 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69110 0 69166 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70214 0 70270 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140318 0 140374 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141422 0 141478 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159822 0 159878 800
rect 160190 0 160246 800
rect 160558 0 160614 800
rect 160926 0 160982 800
rect 161294 0 161350 800
rect 161662 0 161718 800
rect 162030 0 162086 800
rect 162398 0 162454 800
rect 162766 0 162822 800
rect 163134 0 163190 800
rect 163502 0 163558 800
rect 163870 0 163926 800
rect 164238 0 164294 800
rect 164606 0 164662 800
rect 164882 0 164938 800
rect 165250 0 165306 800
rect 165618 0 165674 800
rect 165986 0 166042 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 167090 0 167146 800
rect 167458 0 167514 800
rect 167826 0 167882 800
rect 168194 0 168250 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6586 119354
rect 6754 119144 8058 119354
rect 8226 119144 9622 119354
rect 9790 119144 11094 119354
rect 11262 119144 12566 119354
rect 12734 119144 14038 119354
rect 14206 119144 15510 119354
rect 15678 119144 16982 119354
rect 17150 119144 18546 119354
rect 18714 119144 20018 119354
rect 20186 119144 21490 119354
rect 21658 119144 22962 119354
rect 23130 119144 24434 119354
rect 24602 119144 25906 119354
rect 26074 119144 27470 119354
rect 27638 119144 28942 119354
rect 29110 119144 30414 119354
rect 30582 119144 31886 119354
rect 32054 119144 33358 119354
rect 33526 119144 34830 119354
rect 34998 119144 36394 119354
rect 36562 119144 37866 119354
rect 38034 119144 39338 119354
rect 39506 119144 40810 119354
rect 40978 119144 42282 119354
rect 42450 119144 43846 119354
rect 44014 119144 45318 119354
rect 45486 119144 46790 119354
rect 46958 119144 48262 119354
rect 48430 119144 49734 119354
rect 49902 119144 51206 119354
rect 51374 119144 52770 119354
rect 52938 119144 54242 119354
rect 54410 119144 55714 119354
rect 55882 119144 57186 119354
rect 57354 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61694 119354
rect 61862 119144 63166 119354
rect 63334 119144 64638 119354
rect 64806 119144 66110 119354
rect 66278 119144 67582 119354
rect 67750 119144 69054 119354
rect 69222 119144 70618 119354
rect 70786 119144 72090 119354
rect 72258 119144 73562 119354
rect 73730 119144 75034 119354
rect 75202 119144 76506 119354
rect 76674 119144 78070 119354
rect 78238 119144 79542 119354
rect 79710 119144 81014 119354
rect 81182 119144 82486 119354
rect 82654 119144 83958 119354
rect 84126 119144 85430 119354
rect 85598 119144 86994 119354
rect 87162 119144 88466 119354
rect 88634 119144 89938 119354
rect 90106 119144 91410 119354
rect 91578 119144 92882 119354
rect 93050 119144 94354 119354
rect 94522 119144 95918 119354
rect 96086 119144 97390 119354
rect 97558 119144 98862 119354
rect 99030 119144 100334 119354
rect 100502 119144 101806 119354
rect 101974 119144 103278 119354
rect 103446 119144 104842 119354
rect 105010 119144 106314 119354
rect 106482 119144 107786 119354
rect 107954 119144 109258 119354
rect 109426 119144 110730 119354
rect 110898 119144 112294 119354
rect 112462 119144 113766 119354
rect 113934 119144 115238 119354
rect 115406 119144 116710 119354
rect 116878 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121218 119354
rect 121386 119144 122690 119354
rect 122858 119144 124162 119354
rect 124330 119144 125634 119354
rect 125802 119144 127106 119354
rect 127274 119144 128578 119354
rect 128746 119144 130142 119354
rect 130310 119144 131614 119354
rect 131782 119144 133086 119354
rect 133254 119144 134558 119354
rect 134726 119144 136030 119354
rect 136198 119144 137502 119354
rect 137670 119144 139066 119354
rect 139234 119144 140538 119354
rect 140706 119144 142010 119354
rect 142178 119144 143482 119354
rect 143650 119144 144954 119354
rect 145122 119144 146518 119354
rect 146686 119144 147990 119354
rect 148158 119144 149462 119354
rect 149630 119144 150934 119354
rect 151102 119144 152406 119354
rect 152574 119144 153878 119354
rect 154046 119144 155442 119354
rect 155610 119144 156914 119354
rect 157082 119144 158386 119354
rect 158554 119144 159858 119354
rect 160026 119144 161330 119354
rect 161498 119144 162802 119354
rect 162970 119144 164366 119354
rect 164534 119144 165838 119354
rect 166006 119144 167310 119354
rect 167478 119144 168782 119354
rect 168950 119144 170254 119354
rect 170422 119144 171726 119354
rect 171894 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4378 856
rect 4546 800 4746 856
rect 4914 800 5114 856
rect 5282 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6862 856
rect 7030 800 7230 856
rect 7398 800 7598 856
rect 7766 800 7966 856
rect 8134 800 8334 856
rect 8502 800 8702 856
rect 8870 800 9070 856
rect 9238 800 9438 856
rect 9606 800 9806 856
rect 9974 800 10174 856
rect 10342 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 13026 856
rect 13194 800 13394 856
rect 13562 800 13762 856
rect 13930 800 14130 856
rect 14298 800 14498 856
rect 14666 800 14866 856
rect 15034 800 15234 856
rect 15402 800 15510 856
rect 15678 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16614 856
rect 16782 800 16982 856
rect 17150 800 17350 856
rect 17518 800 17718 856
rect 17886 800 18086 856
rect 18254 800 18454 856
rect 18622 800 18822 856
rect 18990 800 19190 856
rect 19358 800 19558 856
rect 19726 800 19926 856
rect 20094 800 20294 856
rect 20462 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23146 856
rect 23314 800 23514 856
rect 23682 800 23882 856
rect 24050 800 24250 856
rect 24418 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26734 856
rect 26902 800 27102 856
rect 27270 800 27470 856
rect 27638 800 27838 856
rect 28006 800 28206 856
rect 28374 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29310 856
rect 29478 800 29678 856
rect 29846 800 30046 856
rect 30214 800 30414 856
rect 30582 800 30782 856
rect 30950 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33634 856
rect 33802 800 34002 856
rect 34170 800 34370 856
rect 34538 800 34738 856
rect 34906 800 35106 856
rect 35274 800 35474 856
rect 35642 800 35842 856
rect 36010 800 36118 856
rect 36286 800 36486 856
rect 36654 800 36854 856
rect 37022 800 37222 856
rect 37390 800 37590 856
rect 37758 800 37958 856
rect 38126 800 38326 856
rect 38494 800 38694 856
rect 38862 800 39062 856
rect 39230 800 39430 856
rect 39598 800 39798 856
rect 39966 800 40166 856
rect 40334 800 40534 856
rect 40702 800 40902 856
rect 41070 800 41178 856
rect 41346 800 41546 856
rect 41714 800 41914 856
rect 42082 800 42282 856
rect 42450 800 42650 856
rect 42818 800 43018 856
rect 43186 800 43386 856
rect 43554 800 43754 856
rect 43922 800 44122 856
rect 44290 800 44490 856
rect 44658 800 44858 856
rect 45026 800 45226 856
rect 45394 800 45594 856
rect 45762 800 45962 856
rect 46130 800 46330 856
rect 46498 800 46606 856
rect 46774 800 46974 856
rect 47142 800 47342 856
rect 47510 800 47710 856
rect 47878 800 48078 856
rect 48246 800 48446 856
rect 48614 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49550 856
rect 49718 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50654 856
rect 50822 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51666 856
rect 51834 800 52034 856
rect 52202 800 52402 856
rect 52570 800 52770 856
rect 52938 800 53138 856
rect 53306 800 53506 856
rect 53674 800 53874 856
rect 54042 800 54242 856
rect 54410 800 54610 856
rect 54778 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55714 856
rect 55882 800 56082 856
rect 56250 800 56450 856
rect 56618 800 56726 856
rect 56894 800 57094 856
rect 57262 800 57462 856
rect 57630 800 57830 856
rect 57998 800 58198 856
rect 58366 800 58566 856
rect 58734 800 58934 856
rect 59102 800 59302 856
rect 59470 800 59670 856
rect 59838 800 60038 856
rect 60206 800 60406 856
rect 60574 800 60774 856
rect 60942 800 61142 856
rect 61310 800 61510 856
rect 61678 800 61786 856
rect 61954 800 62154 856
rect 62322 800 62522 856
rect 62690 800 62890 856
rect 63058 800 63258 856
rect 63426 800 63626 856
rect 63794 800 63994 856
rect 64162 800 64362 856
rect 64530 800 64730 856
rect 64898 800 65098 856
rect 65266 800 65466 856
rect 65634 800 65834 856
rect 66002 800 66202 856
rect 66370 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68318 856
rect 68486 800 68686 856
rect 68854 800 69054 856
rect 69222 800 69422 856
rect 69590 800 69790 856
rect 69958 800 70158 856
rect 70326 800 70526 856
rect 70694 800 70894 856
rect 71062 800 71262 856
rect 71430 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72274 856
rect 72442 800 72642 856
rect 72810 800 73010 856
rect 73178 800 73378 856
rect 73546 800 73746 856
rect 73914 800 74114 856
rect 74282 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75218 856
rect 75386 800 75586 856
rect 75754 800 75954 856
rect 76122 800 76322 856
rect 76490 800 76690 856
rect 76858 800 77058 856
rect 77226 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78806 856
rect 78974 800 79174 856
rect 79342 800 79542 856
rect 79710 800 79910 856
rect 80078 800 80278 856
rect 80446 800 80646 856
rect 80814 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81750 856
rect 81918 800 82118 856
rect 82286 800 82394 856
rect 82562 800 82762 856
rect 82930 800 83130 856
rect 83298 800 83498 856
rect 83666 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85338 856
rect 85506 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87454 856
rect 87622 800 87822 856
rect 87990 800 88190 856
rect 88358 800 88558 856
rect 88726 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90398 856
rect 90566 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93250 856
rect 93418 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96194 856
rect 96362 800 96562 856
rect 96730 800 96930 856
rect 97098 800 97298 856
rect 97466 800 97666 856
rect 97834 800 97942 856
rect 98110 800 98310 856
rect 98478 800 98678 856
rect 98846 800 99046 856
rect 99214 800 99414 856
rect 99582 800 99782 856
rect 99950 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101254 856
rect 101422 800 101622 856
rect 101790 800 101990 856
rect 102158 800 102358 856
rect 102526 800 102726 856
rect 102894 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104842 856
rect 105010 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105946 856
rect 106114 800 106314 856
rect 106482 800 106682 856
rect 106850 800 107050 856
rect 107218 800 107418 856
rect 107586 800 107786 856
rect 107954 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108798 856
rect 108966 800 109166 856
rect 109334 800 109534 856
rect 109702 800 109902 856
rect 110070 800 110270 856
rect 110438 800 110638 856
rect 110806 800 111006 856
rect 111174 800 111374 856
rect 111542 800 111742 856
rect 111910 800 112110 856
rect 112278 800 112478 856
rect 112646 800 112846 856
rect 113014 800 113214 856
rect 113382 800 113490 856
rect 113658 800 113858 856
rect 114026 800 114226 856
rect 114394 800 114594 856
rect 114762 800 114962 856
rect 115130 800 115330 856
rect 115498 800 115698 856
rect 115866 800 116066 856
rect 116234 800 116434 856
rect 116602 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117538 856
rect 117706 800 117906 856
rect 118074 800 118274 856
rect 118442 800 118550 856
rect 118718 800 118918 856
rect 119086 800 119286 856
rect 119454 800 119654 856
rect 119822 800 120022 856
rect 120190 800 120390 856
rect 120558 800 120758 856
rect 120926 800 121126 856
rect 121294 800 121494 856
rect 121662 800 121862 856
rect 122030 800 122230 856
rect 122398 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123610 856
rect 123778 800 123978 856
rect 124146 800 124346 856
rect 124514 800 124714 856
rect 124882 800 125082 856
rect 125250 800 125450 856
rect 125618 800 125818 856
rect 125986 800 126186 856
rect 126354 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127290 856
rect 127458 800 127658 856
rect 127826 800 128026 856
rect 128194 800 128394 856
rect 128562 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130510 856
rect 130678 800 130878 856
rect 131046 800 131246 856
rect 131414 800 131614 856
rect 131782 800 131982 856
rect 132150 800 132350 856
rect 132518 800 132718 856
rect 132886 800 133086 856
rect 133254 800 133454 856
rect 133622 800 133730 856
rect 133898 800 134098 856
rect 134266 800 134466 856
rect 134634 800 134834 856
rect 135002 800 135202 856
rect 135370 800 135570 856
rect 135738 800 135938 856
rect 136106 800 136306 856
rect 136474 800 136674 856
rect 136842 800 137042 856
rect 137210 800 137410 856
rect 137578 800 137778 856
rect 137946 800 138146 856
rect 138314 800 138514 856
rect 138682 800 138882 856
rect 139050 800 139158 856
rect 139326 800 139526 856
rect 139694 800 139894 856
rect 140062 800 140262 856
rect 140430 800 140630 856
rect 140798 800 140998 856
rect 141166 800 141366 856
rect 141534 800 141734 856
rect 141902 800 142102 856
rect 142270 800 142470 856
rect 142638 800 142838 856
rect 143006 800 143206 856
rect 143374 800 143574 856
rect 143742 800 143942 856
rect 144110 800 144218 856
rect 144386 800 144586 856
rect 144754 800 144954 856
rect 145122 800 145322 856
rect 145490 800 145690 856
rect 145858 800 146058 856
rect 146226 800 146426 856
rect 146594 800 146794 856
rect 146962 800 147162 856
rect 147330 800 147530 856
rect 147698 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 149002 856
rect 149170 800 149278 856
rect 149446 800 149646 856
rect 149814 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150750 856
rect 150918 800 151118 856
rect 151286 800 151486 856
rect 151654 800 151854 856
rect 152022 800 152222 856
rect 152390 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153326 856
rect 153494 800 153694 856
rect 153862 800 154062 856
rect 154230 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159766 856
rect 159934 800 160134 856
rect 160302 800 160502 856
rect 160670 800 160870 856
rect 161038 800 161238 856
rect 161406 800 161606 856
rect 161774 800 161974 856
rect 162142 800 162342 856
rect 162510 800 162710 856
rect 162878 800 163078 856
rect 163246 800 163446 856
rect 163614 800 163814 856
rect 163982 800 164182 856
rect 164350 800 164550 856
rect 164718 800 164826 856
rect 164994 800 165194 856
rect 165362 800 165562 856
rect 165730 800 165930 856
rect 166098 800 166298 856
rect 166466 800 166666 856
rect 166834 800 167034 856
rect 167202 800 167402 856
rect 167570 800 167770 856
rect 167938 800 168138 856
rect 168306 800 168506 856
rect 168674 800 168874 856
rect 169042 800 169242 856
rect 169410 800 169610 856
rect 169778 800 169886 856
rect 170054 800 170254 856
rect 170422 800 170622 856
rect 170790 800 170990 856
rect 171158 800 171358 856
rect 171526 800 171726 856
rect 171894 800 172094 856
rect 172262 800 172462 856
rect 172630 800 172830 856
rect 172998 800 173198 856
rect 173366 800 173566 856
rect 173734 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 174946 856
rect 175114 800 175314 856
rect 175482 800 175682 856
rect 175850 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178186 856
<< metal3 >>
rect 0 114384 800 114504
rect 179200 112344 180000 112464
rect 0 103504 800 103624
rect 179200 97384 180000 97504
rect 0 92624 800 92744
rect 179200 82424 180000 82544
rect 0 81744 800 81864
rect 0 70864 800 70984
rect 179200 67464 180000 67584
rect 0 59848 800 59968
rect 179200 52368 180000 52488
rect 0 48968 800 49088
rect 0 38088 800 38208
rect 179200 37408 180000 37528
rect 0 27208 800 27328
rect 179200 22448 180000 22568
rect 0 16328 800 16448
rect 179200 7488 180000 7608
rect 0 5448 800 5568
<< obsm3 >>
rect 800 114584 179200 118149
rect 880 114304 179200 114584
rect 800 112544 179200 114304
rect 800 112264 179120 112544
rect 800 103704 179200 112264
rect 880 103424 179200 103704
rect 800 97584 179200 103424
rect 800 97304 179120 97584
rect 800 92824 179200 97304
rect 880 92544 179200 92824
rect 800 82624 179200 92544
rect 800 82344 179120 82624
rect 800 81944 179200 82344
rect 880 81664 179200 81944
rect 800 71064 179200 81664
rect 880 70784 179200 71064
rect 800 67664 179200 70784
rect 800 67384 179120 67664
rect 800 60048 179200 67384
rect 880 59768 179200 60048
rect 800 52568 179200 59768
rect 800 52288 179120 52568
rect 800 49168 179200 52288
rect 880 48888 179200 49168
rect 800 38288 179200 48888
rect 880 38008 179200 38288
rect 800 37608 179200 38008
rect 800 37328 179120 37608
rect 800 27408 179200 37328
rect 880 27128 179200 27408
rect 800 22648 179200 27128
rect 800 22368 179120 22648
rect 800 16528 179200 22368
rect 880 16248 179200 16528
rect 800 7688 179200 16248
rect 800 7408 179120 7688
rect 800 5648 179200 7408
rect 880 5368 179200 5648
rect 800 2143 179200 5368
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 65011 117632 98013 118149
rect 65011 109787 65568 117632
rect 66048 109787 80928 117632
rect 81408 109787 96288 117632
rect 96768 109787 98013 117632
<< labels >>
rlabel metal3 s 0 5448 800 5568 6 active
port 1 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal3 s 179200 52368 180000 52488 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 179200 67464 180000 67584 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal3 s 0 70864 800 70984 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal3 s 0 81744 800 81864 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 0 27208 800 27328 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal3 s 0 92624 800 92744 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 179200 82424 180000 82544 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal3 s 0 103504 800 103624 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal3 s 0 114384 800 114504 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal3 s 179200 97384 180000 97504 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 179200 112344 180000 112464 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 0 38088 800 38208 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 0 48968 800 49088 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal2 s 170310 119200 170366 120000 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 0 59848 800 59968 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal2 s 171782 119200 171838 120000 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 45374 119200 45430 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 49790 119200 49846 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 54298 119200 54354 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 58714 119200 58770 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 63222 119200 63278 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 67638 119200 67694 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 81070 119200 81126 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 85486 119200 85542 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 89994 119200 90050 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 94410 119200 94466 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 98918 119200 98974 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 103334 119200 103390 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 107842 119200 107898 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 116766 119200 116822 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 121274 119200 121330 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 125690 119200 125746 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 130198 119200 130254 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 148046 119200 148102 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 152462 119200 152518 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 156970 119200 157026 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 161386 119200 161442 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 165894 119200 165950 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 14094 119200 14150 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18602 119200 18658 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 23018 119200 23074 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 27526 119200 27582 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31942 119200 31998 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 36450 119200 36506 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 40866 119200 40922 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 46846 119200 46902 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 69110 119200 69166 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 73618 119200 73674 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 95974 119200 96030 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 100390 119200 100446 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 104898 119200 104954 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 109314 119200 109370 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 113822 119200 113878 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 122746 119200 122802 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 127162 119200 127218 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 131670 119200 131726 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 11150 119200 11206 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 140594 119200 140650 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 145010 119200 145066 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 149518 119200 149574 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 158442 119200 158498 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 162858 119200 162914 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15566 119200 15622 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 33414 119200 33470 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 37922 119200 37978 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 42338 119200 42394 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 48318 119200 48374 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 57242 119200 57298 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 61750 119200 61806 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 66166 119200 66222 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 84014 119200 84070 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 92938 119200 92994 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 101862 119200 101918 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 128634 119200 128690 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 133142 119200 133198 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12622 119200 12678 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 137558 119200 137614 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 142066 119200 142122 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 146574 119200 146630 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 150990 119200 151046 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 159914 119200 159970 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 164422 119200 164478 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 168838 119200 168894 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 17038 119200 17094 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21546 119200 21602 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 43902 119200 43958 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 163502 0 163558 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72330 0 72386 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 98366 0 98422 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 118974 0 119030 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 179200 7488 180000 7608 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 user_irq[0]
port 530 nsew signal output
rlabel metal3 s 179200 22448 180000 22568 6 user_irq[1]
port 531 nsew signal output
rlabel metal3 s 179200 37408 180000 37528 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6680776
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_10.magic.gds
string GDS_START 295056
<< end >>

