magic
tech sky130A
magscale 1 2
timestamp 1654261361
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 117972
<< metal2 >>
rect 662 119200 718 120000
rect 2042 119200 2098 120000
rect 3514 119200 3570 120000
rect 4986 119200 5042 120000
rect 6458 119200 6514 120000
rect 7838 119200 7894 120000
rect 9310 119200 9366 120000
rect 10782 119200 10838 120000
rect 12254 119200 12310 120000
rect 13726 119200 13782 120000
rect 15106 119200 15162 120000
rect 16578 119200 16634 120000
rect 18050 119200 18106 120000
rect 19522 119200 19578 120000
rect 20902 119200 20958 120000
rect 22374 119200 22430 120000
rect 23846 119200 23902 120000
rect 25318 119200 25374 120000
rect 26790 119200 26846 120000
rect 28170 119200 28226 120000
rect 29642 119200 29698 120000
rect 31114 119200 31170 120000
rect 32586 119200 32642 120000
rect 33966 119200 34022 120000
rect 35438 119200 35494 120000
rect 36910 119200 36966 120000
rect 38382 119200 38438 120000
rect 39854 119200 39910 120000
rect 41234 119200 41290 120000
rect 42706 119200 42762 120000
rect 44178 119200 44234 120000
rect 45650 119200 45706 120000
rect 47122 119200 47178 120000
rect 48502 119200 48558 120000
rect 49974 119200 50030 120000
rect 51446 119200 51502 120000
rect 52918 119200 52974 120000
rect 54298 119200 54354 120000
rect 55770 119200 55826 120000
rect 57242 119200 57298 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61566 119200 61622 120000
rect 63038 119200 63094 120000
rect 64510 119200 64566 120000
rect 65982 119200 66038 120000
rect 67362 119200 67418 120000
rect 68834 119200 68890 120000
rect 70306 119200 70362 120000
rect 71778 119200 71834 120000
rect 73250 119200 73306 120000
rect 74630 119200 74686 120000
rect 76102 119200 76158 120000
rect 77574 119200 77630 120000
rect 79046 119200 79102 120000
rect 80518 119200 80574 120000
rect 81898 119200 81954 120000
rect 83370 119200 83426 120000
rect 84842 119200 84898 120000
rect 86314 119200 86370 120000
rect 87694 119200 87750 120000
rect 89166 119200 89222 120000
rect 90638 119200 90694 120000
rect 92110 119200 92166 120000
rect 93582 119200 93638 120000
rect 94962 119200 95018 120000
rect 96434 119200 96490 120000
rect 97906 119200 97962 120000
rect 99378 119200 99434 120000
rect 100758 119200 100814 120000
rect 102230 119200 102286 120000
rect 103702 119200 103758 120000
rect 105174 119200 105230 120000
rect 106646 119200 106702 120000
rect 108026 119200 108082 120000
rect 109498 119200 109554 120000
rect 110970 119200 111026 120000
rect 112442 119200 112498 120000
rect 113914 119200 113970 120000
rect 115294 119200 115350 120000
rect 116766 119200 116822 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121090 119200 121146 120000
rect 122562 119200 122618 120000
rect 124034 119200 124090 120000
rect 125506 119200 125562 120000
rect 126978 119200 127034 120000
rect 128358 119200 128414 120000
rect 129830 119200 129886 120000
rect 131302 119200 131358 120000
rect 132774 119200 132830 120000
rect 134154 119200 134210 120000
rect 135626 119200 135682 120000
rect 137098 119200 137154 120000
rect 138570 119200 138626 120000
rect 140042 119200 140098 120000
rect 141422 119200 141478 120000
rect 142894 119200 142950 120000
rect 144366 119200 144422 120000
rect 145838 119200 145894 120000
rect 147310 119200 147366 120000
rect 148690 119200 148746 120000
rect 150162 119200 150218 120000
rect 151634 119200 151690 120000
rect 153106 119200 153162 120000
rect 154486 119200 154542 120000
rect 155958 119200 156014 120000
rect 157430 119200 157486 120000
rect 158902 119200 158958 120000
rect 160374 119200 160430 120000
rect 161754 119200 161810 120000
rect 163226 119200 163282 120000
rect 164698 119200 164754 120000
rect 166170 119200 166226 120000
rect 167550 119200 167606 120000
rect 169022 119200 169078 120000
rect 170494 119200 170550 120000
rect 171966 119200 172022 120000
rect 173438 119200 173494 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37002 0 37058 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38106 0 38162 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54758 0 54814 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95330 0 95386 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106922 0 106978 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 108026 0 108082 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122838 0 122894 800
rect 123206 0 123262 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138110 0 138166 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 142066 0 142122 800
rect 142434 0 142490 800
rect 142802 0 142858 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143906 0 143962 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145010 0 145066 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147862 0 147918 800
rect 148230 0 148286 800
rect 148598 0 148654 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156878 0 156934 800
rect 157246 0 157302 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160190 0 160246 800
rect 160558 0 160614 800
rect 160926 0 160982 800
rect 161294 0 161350 800
rect 161662 0 161718 800
rect 162030 0 162086 800
rect 162398 0 162454 800
rect 162674 0 162730 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163778 0 163834 800
rect 164146 0 164202 800
rect 164514 0 164570 800
rect 164882 0 164938 800
rect 165250 0 165306 800
rect 165618 0 165674 800
rect 165986 0 166042 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 167090 0 167146 800
rect 167458 0 167514 800
rect 167826 0 167882 800
rect 168194 0 168250 800
rect 168470 0 168526 800
rect 168838 0 168894 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 774 119144 1986 119354
rect 2154 119144 3458 119354
rect 3626 119144 4930 119354
rect 5098 119144 6402 119354
rect 6570 119144 7782 119354
rect 7950 119144 9254 119354
rect 9422 119144 10726 119354
rect 10894 119144 12198 119354
rect 12366 119144 13670 119354
rect 13838 119144 15050 119354
rect 15218 119144 16522 119354
rect 16690 119144 17994 119354
rect 18162 119144 19466 119354
rect 19634 119144 20846 119354
rect 21014 119144 22318 119354
rect 22486 119144 23790 119354
rect 23958 119144 25262 119354
rect 25430 119144 26734 119354
rect 26902 119144 28114 119354
rect 28282 119144 29586 119354
rect 29754 119144 31058 119354
rect 31226 119144 32530 119354
rect 32698 119144 33910 119354
rect 34078 119144 35382 119354
rect 35550 119144 36854 119354
rect 37022 119144 38326 119354
rect 38494 119144 39798 119354
rect 39966 119144 41178 119354
rect 41346 119144 42650 119354
rect 42818 119144 44122 119354
rect 44290 119144 45594 119354
rect 45762 119144 47066 119354
rect 47234 119144 48446 119354
rect 48614 119144 49918 119354
rect 50086 119144 51390 119354
rect 51558 119144 52862 119354
rect 53030 119144 54242 119354
rect 54410 119144 55714 119354
rect 55882 119144 57186 119354
rect 57354 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61510 119354
rect 61678 119144 62982 119354
rect 63150 119144 64454 119354
rect 64622 119144 65926 119354
rect 66094 119144 67306 119354
rect 67474 119144 68778 119354
rect 68946 119144 70250 119354
rect 70418 119144 71722 119354
rect 71890 119144 73194 119354
rect 73362 119144 74574 119354
rect 74742 119144 76046 119354
rect 76214 119144 77518 119354
rect 77686 119144 78990 119354
rect 79158 119144 80462 119354
rect 80630 119144 81842 119354
rect 82010 119144 83314 119354
rect 83482 119144 84786 119354
rect 84954 119144 86258 119354
rect 86426 119144 87638 119354
rect 87806 119144 89110 119354
rect 89278 119144 90582 119354
rect 90750 119144 92054 119354
rect 92222 119144 93526 119354
rect 93694 119144 94906 119354
rect 95074 119144 96378 119354
rect 96546 119144 97850 119354
rect 98018 119144 99322 119354
rect 99490 119144 100702 119354
rect 100870 119144 102174 119354
rect 102342 119144 103646 119354
rect 103814 119144 105118 119354
rect 105286 119144 106590 119354
rect 106758 119144 107970 119354
rect 108138 119144 109442 119354
rect 109610 119144 110914 119354
rect 111082 119144 112386 119354
rect 112554 119144 113858 119354
rect 114026 119144 115238 119354
rect 115406 119144 116710 119354
rect 116878 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121034 119354
rect 121202 119144 122506 119354
rect 122674 119144 123978 119354
rect 124146 119144 125450 119354
rect 125618 119144 126922 119354
rect 127090 119144 128302 119354
rect 128470 119144 129774 119354
rect 129942 119144 131246 119354
rect 131414 119144 132718 119354
rect 132886 119144 134098 119354
rect 134266 119144 135570 119354
rect 135738 119144 137042 119354
rect 137210 119144 138514 119354
rect 138682 119144 139986 119354
rect 140154 119144 141366 119354
rect 141534 119144 142838 119354
rect 143006 119144 144310 119354
rect 144478 119144 145782 119354
rect 145950 119144 147254 119354
rect 147422 119144 148634 119354
rect 148802 119144 150106 119354
rect 150274 119144 151578 119354
rect 151746 119144 153050 119354
rect 153218 119144 154430 119354
rect 154598 119144 155902 119354
rect 156070 119144 157374 119354
rect 157542 119144 158846 119354
rect 159014 119144 160318 119354
rect 160486 119144 161698 119354
rect 161866 119144 163170 119354
rect 163338 119144 164642 119354
rect 164810 119144 166114 119354
rect 166282 119144 167494 119354
rect 167662 119144 168966 119354
rect 169134 119144 170438 119354
rect 170606 119144 171910 119354
rect 172078 119144 173382 119354
rect 173550 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6126 856
rect 6294 734 6494 856
rect 6662 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7966 856
rect 8134 734 8334 856
rect 8502 734 8702 856
rect 8870 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9806 856
rect 9974 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 11922 856
rect 12090 734 12290 856
rect 12458 734 12658 856
rect 12826 734 13026 856
rect 13194 734 13394 856
rect 13562 734 13762 856
rect 13930 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14866 856
rect 15034 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15970 856
rect 16138 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17718 856
rect 17886 734 18086 856
rect 18254 734 18454 856
rect 18622 734 18822 856
rect 18990 734 19190 856
rect 19358 734 19558 856
rect 19726 734 19926 856
rect 20094 734 20294 856
rect 20462 734 20662 856
rect 20830 734 21030 856
rect 21198 734 21398 856
rect 21566 734 21766 856
rect 21934 734 22134 856
rect 22302 734 22502 856
rect 22670 734 22870 856
rect 23038 734 23238 856
rect 23406 734 23514 856
rect 23682 734 23882 856
rect 24050 734 24250 856
rect 24418 734 24618 856
rect 24786 734 24986 856
rect 25154 734 25354 856
rect 25522 734 25722 856
rect 25890 734 26090 856
rect 26258 734 26458 856
rect 26626 734 26826 856
rect 26994 734 27194 856
rect 27362 734 27562 856
rect 27730 734 27930 856
rect 28098 734 28298 856
rect 28466 734 28666 856
rect 28834 734 29034 856
rect 29202 734 29310 856
rect 29478 734 29678 856
rect 29846 734 30046 856
rect 30214 734 30414 856
rect 30582 734 30782 856
rect 30950 734 31150 856
rect 31318 734 31518 856
rect 31686 734 31886 856
rect 32054 734 32254 856
rect 32422 734 32622 856
rect 32790 734 32990 856
rect 33158 734 33358 856
rect 33526 734 33726 856
rect 33894 734 34094 856
rect 34262 734 34462 856
rect 34630 734 34830 856
rect 34998 734 35106 856
rect 35274 734 35474 856
rect 35642 734 35842 856
rect 36010 734 36210 856
rect 36378 734 36578 856
rect 36746 734 36946 856
rect 37114 734 37314 856
rect 37482 734 37682 856
rect 37850 734 38050 856
rect 38218 734 38418 856
rect 38586 734 38786 856
rect 38954 734 39154 856
rect 39322 734 39522 856
rect 39690 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40626 856
rect 40794 734 40902 856
rect 41070 734 41270 856
rect 41438 734 41638 856
rect 41806 734 42006 856
rect 42174 734 42374 856
rect 42542 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43478 856
rect 43646 734 43846 856
rect 44014 734 44214 856
rect 44382 734 44582 856
rect 44750 734 44950 856
rect 45118 734 45318 856
rect 45486 734 45686 856
rect 45854 734 46054 856
rect 46222 734 46422 856
rect 46590 734 46698 856
rect 46866 734 47066 856
rect 47234 734 47434 856
rect 47602 734 47802 856
rect 47970 734 48170 856
rect 48338 734 48538 856
rect 48706 734 48906 856
rect 49074 734 49274 856
rect 49442 734 49642 856
rect 49810 734 50010 856
rect 50178 734 50378 856
rect 50546 734 50746 856
rect 50914 734 51114 856
rect 51282 734 51482 856
rect 51650 734 51850 856
rect 52018 734 52218 856
rect 52386 734 52494 856
rect 52662 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53966 856
rect 54134 734 54334 856
rect 54502 734 54702 856
rect 54870 734 55070 856
rect 55238 734 55438 856
rect 55606 734 55806 856
rect 55974 734 56174 856
rect 56342 734 56542 856
rect 56710 734 56910 856
rect 57078 734 57278 856
rect 57446 734 57646 856
rect 57814 734 58014 856
rect 58182 734 58290 856
rect 58458 734 58658 856
rect 58826 734 59026 856
rect 59194 734 59394 856
rect 59562 734 59762 856
rect 59930 734 60130 856
rect 60298 734 60498 856
rect 60666 734 60866 856
rect 61034 734 61234 856
rect 61402 734 61602 856
rect 61770 734 61970 856
rect 62138 734 62338 856
rect 62506 734 62706 856
rect 62874 734 63074 856
rect 63242 734 63442 856
rect 63610 734 63810 856
rect 63978 734 64086 856
rect 64254 734 64454 856
rect 64622 734 64822 856
rect 64990 734 65190 856
rect 65358 734 65558 856
rect 65726 734 65926 856
rect 66094 734 66294 856
rect 66462 734 66662 856
rect 66830 734 67030 856
rect 67198 734 67398 856
rect 67566 734 67766 856
rect 67934 734 68134 856
rect 68302 734 68502 856
rect 68670 734 68870 856
rect 69038 734 69238 856
rect 69406 734 69606 856
rect 69774 734 69882 856
rect 70050 734 70250 856
rect 70418 734 70618 856
rect 70786 734 70986 856
rect 71154 734 71354 856
rect 71522 734 71722 856
rect 71890 734 72090 856
rect 72258 734 72458 856
rect 72626 734 72826 856
rect 72994 734 73194 856
rect 73362 734 73562 856
rect 73730 734 73930 856
rect 74098 734 74298 856
rect 74466 734 74666 856
rect 74834 734 75034 856
rect 75202 734 75402 856
rect 75570 734 75678 856
rect 75846 734 76046 856
rect 76214 734 76414 856
rect 76582 734 76782 856
rect 76950 734 77150 856
rect 77318 734 77518 856
rect 77686 734 77886 856
rect 78054 734 78254 856
rect 78422 734 78622 856
rect 78790 734 78990 856
rect 79158 734 79358 856
rect 79526 734 79726 856
rect 79894 734 80094 856
rect 80262 734 80462 856
rect 80630 734 80830 856
rect 80998 734 81198 856
rect 81366 734 81474 856
rect 81642 734 81842 856
rect 82010 734 82210 856
rect 82378 734 82578 856
rect 82746 734 82946 856
rect 83114 734 83314 856
rect 83482 734 83682 856
rect 83850 734 84050 856
rect 84218 734 84418 856
rect 84586 734 84786 856
rect 84954 734 85154 856
rect 85322 734 85522 856
rect 85690 734 85890 856
rect 86058 734 86258 856
rect 86426 734 86626 856
rect 86794 734 86994 856
rect 87162 734 87270 856
rect 87438 734 87638 856
rect 87806 734 88006 856
rect 88174 734 88374 856
rect 88542 734 88742 856
rect 88910 734 89110 856
rect 89278 734 89478 856
rect 89646 734 89846 856
rect 90014 734 90214 856
rect 90382 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91318 856
rect 91486 734 91686 856
rect 91854 734 92054 856
rect 92222 734 92422 856
rect 92590 734 92790 856
rect 92958 734 93066 856
rect 93234 734 93434 856
rect 93602 734 93802 856
rect 93970 734 94170 856
rect 94338 734 94538 856
rect 94706 734 94906 856
rect 95074 734 95274 856
rect 95442 734 95642 856
rect 95810 734 96010 856
rect 96178 734 96378 856
rect 96546 734 96746 856
rect 96914 734 97114 856
rect 97282 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98218 856
rect 98386 734 98586 856
rect 98754 734 98862 856
rect 99030 734 99230 856
rect 99398 734 99598 856
rect 99766 734 99966 856
rect 100134 734 100334 856
rect 100502 734 100702 856
rect 100870 734 101070 856
rect 101238 734 101438 856
rect 101606 734 101806 856
rect 101974 734 102174 856
rect 102342 734 102542 856
rect 102710 734 102910 856
rect 103078 734 103278 856
rect 103446 734 103646 856
rect 103814 734 104014 856
rect 104182 734 104382 856
rect 104550 734 104658 856
rect 104826 734 105026 856
rect 105194 734 105394 856
rect 105562 734 105762 856
rect 105930 734 106130 856
rect 106298 734 106498 856
rect 106666 734 106866 856
rect 107034 734 107234 856
rect 107402 734 107602 856
rect 107770 734 107970 856
rect 108138 734 108338 856
rect 108506 734 108706 856
rect 108874 734 109074 856
rect 109242 734 109442 856
rect 109610 734 109810 856
rect 109978 734 110178 856
rect 110346 734 110454 856
rect 110622 734 110822 856
rect 110990 734 111190 856
rect 111358 734 111558 856
rect 111726 734 111926 856
rect 112094 734 112294 856
rect 112462 734 112662 856
rect 112830 734 113030 856
rect 113198 734 113398 856
rect 113566 734 113766 856
rect 113934 734 114134 856
rect 114302 734 114502 856
rect 114670 734 114870 856
rect 115038 734 115238 856
rect 115406 734 115606 856
rect 115774 734 115974 856
rect 116142 734 116250 856
rect 116418 734 116618 856
rect 116786 734 116986 856
rect 117154 734 117354 856
rect 117522 734 117722 856
rect 117890 734 118090 856
rect 118258 734 118458 856
rect 118626 734 118826 856
rect 118994 734 119194 856
rect 119362 734 119562 856
rect 119730 734 119930 856
rect 120098 734 120298 856
rect 120466 734 120666 856
rect 120834 734 121034 856
rect 121202 734 121402 856
rect 121570 734 121770 856
rect 121938 734 122046 856
rect 122214 734 122414 856
rect 122582 734 122782 856
rect 122950 734 123150 856
rect 123318 734 123518 856
rect 123686 734 123886 856
rect 124054 734 124254 856
rect 124422 734 124622 856
rect 124790 734 124990 856
rect 125158 734 125358 856
rect 125526 734 125726 856
rect 125894 734 126094 856
rect 126262 734 126462 856
rect 126630 734 126830 856
rect 126998 734 127198 856
rect 127366 734 127566 856
rect 127734 734 127842 856
rect 128010 734 128210 856
rect 128378 734 128578 856
rect 128746 734 128946 856
rect 129114 734 129314 856
rect 129482 734 129682 856
rect 129850 734 130050 856
rect 130218 734 130418 856
rect 130586 734 130786 856
rect 130954 734 131154 856
rect 131322 734 131522 856
rect 131690 734 131890 856
rect 132058 734 132258 856
rect 132426 734 132626 856
rect 132794 734 132994 856
rect 133162 734 133362 856
rect 133530 734 133638 856
rect 133806 734 134006 856
rect 134174 734 134374 856
rect 134542 734 134742 856
rect 134910 734 135110 856
rect 135278 734 135478 856
rect 135646 734 135846 856
rect 136014 734 136214 856
rect 136382 734 136582 856
rect 136750 734 136950 856
rect 137118 734 137318 856
rect 137486 734 137686 856
rect 137854 734 138054 856
rect 138222 734 138422 856
rect 138590 734 138790 856
rect 138958 734 139158 856
rect 139326 734 139434 856
rect 139602 734 139802 856
rect 139970 734 140170 856
rect 140338 734 140538 856
rect 140706 734 140906 856
rect 141074 734 141274 856
rect 141442 734 141642 856
rect 141810 734 142010 856
rect 142178 734 142378 856
rect 142546 734 142746 856
rect 142914 734 143114 856
rect 143282 734 143482 856
rect 143650 734 143850 856
rect 144018 734 144218 856
rect 144386 734 144586 856
rect 144754 734 144954 856
rect 145122 734 145230 856
rect 145398 734 145598 856
rect 145766 734 145966 856
rect 146134 734 146334 856
rect 146502 734 146702 856
rect 146870 734 147070 856
rect 147238 734 147438 856
rect 147606 734 147806 856
rect 147974 734 148174 856
rect 148342 734 148542 856
rect 148710 734 148910 856
rect 149078 734 149278 856
rect 149446 734 149646 856
rect 149814 734 150014 856
rect 150182 734 150382 856
rect 150550 734 150750 856
rect 150918 734 151026 856
rect 151194 734 151394 856
rect 151562 734 151762 856
rect 151930 734 152130 856
rect 152298 734 152498 856
rect 152666 734 152866 856
rect 153034 734 153234 856
rect 153402 734 153602 856
rect 153770 734 153970 856
rect 154138 734 154338 856
rect 154506 734 154706 856
rect 154874 734 155074 856
rect 155242 734 155442 856
rect 155610 734 155810 856
rect 155978 734 156178 856
rect 156346 734 156546 856
rect 156714 734 156822 856
rect 156990 734 157190 856
rect 157358 734 157558 856
rect 157726 734 157926 856
rect 158094 734 158294 856
rect 158462 734 158662 856
rect 158830 734 159030 856
rect 159198 734 159398 856
rect 159566 734 159766 856
rect 159934 734 160134 856
rect 160302 734 160502 856
rect 160670 734 160870 856
rect 161038 734 161238 856
rect 161406 734 161606 856
rect 161774 734 161974 856
rect 162142 734 162342 856
rect 162510 734 162618 856
rect 162786 734 162986 856
rect 163154 734 163354 856
rect 163522 734 163722 856
rect 163890 734 164090 856
rect 164258 734 164458 856
rect 164626 734 164826 856
rect 164994 734 165194 856
rect 165362 734 165562 856
rect 165730 734 165930 856
rect 166098 734 166298 856
rect 166466 734 166666 856
rect 166834 734 167034 856
rect 167202 734 167402 856
rect 167570 734 167770 856
rect 167938 734 168138 856
rect 168306 734 168414 856
rect 168582 734 168782 856
rect 168950 734 169150 856
rect 169318 734 169518 856
rect 169686 734 169886 856
rect 170054 734 170254 856
rect 170422 734 170622 856
rect 170790 734 170990 856
rect 171158 734 171358 856
rect 171526 734 171726 856
rect 171894 734 172094 856
rect 172262 734 172462 856
rect 172630 734 172830 856
rect 172998 734 173198 856
rect 173366 734 173566 856
rect 173734 734 173934 856
rect 174102 734 174210 856
rect 174378 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175314 856
rect 175482 734 175682 856
rect 175850 734 176050 856
rect 176218 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178186 856
<< metal3 >>
rect 0 113296 800 113416
rect 179200 112344 180000 112464
rect 0 99968 800 100088
rect 179200 97384 180000 97504
rect 0 86640 800 86760
rect 179200 82424 180000 82544
rect 0 73312 800 73432
rect 179200 67464 180000 67584
rect 0 59984 800 60104
rect 179200 52368 180000 52488
rect 0 46656 800 46776
rect 179200 37408 180000 37528
rect 0 33328 800 33448
rect 179200 22448 180000 22568
rect 0 20000 800 20120
rect 179200 7488 180000 7608
rect 0 6672 800 6792
<< obsm3 >>
rect 800 113496 179200 117537
rect 880 113216 179200 113496
rect 800 112544 179200 113216
rect 800 112264 179120 112544
rect 800 100168 179200 112264
rect 880 99888 179200 100168
rect 800 97584 179200 99888
rect 800 97304 179120 97584
rect 800 86840 179200 97304
rect 880 86560 179200 86840
rect 800 82624 179200 86560
rect 800 82344 179120 82624
rect 800 73512 179200 82344
rect 880 73232 179200 73512
rect 800 67664 179200 73232
rect 800 67384 179120 67664
rect 800 60184 179200 67384
rect 880 59904 179200 60184
rect 800 52568 179200 59904
rect 800 52288 179120 52568
rect 800 46856 179200 52288
rect 880 46576 179200 46856
rect 800 37608 179200 46576
rect 800 37328 179120 37608
rect 800 33528 179200 37328
rect 880 33248 179200 33528
rect 800 22648 179200 33248
rect 800 22368 179120 22648
rect 800 20200 179200 22368
rect 880 19920 179200 20200
rect 800 7688 179200 19920
rect 800 7408 179120 7688
rect 800 6872 179200 7408
rect 880 6592 179200 6872
rect 800 2143 179200 6592
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 84699 110875 93229 117333
<< labels >>
rlabel metal3 s 179200 7488 180000 7608 6 active
port 1 nsew signal input
rlabel metal3 s 179200 22448 180000 22568 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 0 86640 800 86760 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal2 s 170494 119200 170550 120000 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 179200 67464 180000 67584 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 0 99968 800 100088 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 171966 119200 172022 120000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal3 s 179200 82424 180000 82544 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal2 s 173438 119200 173494 120000 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 179200 97384 180000 97504 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 179200 37408 180000 37528 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 0 113296 800 113416 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal3 s 179200 112344 180000 112464 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 0 33328 800 33448 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal2 s 167550 119200 167606 120000 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal2 s 169022 119200 169078 120000 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 0 73312 800 73432 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 179200 52368 180000 52488 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 44178 119200 44234 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 48502 119200 48558 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 52918 119200 52974 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 57242 119200 57298 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 61566 119200 61622 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 65982 119200 66038 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 70306 119200 70362 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 74630 119200 74686 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 79046 119200 79102 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 83370 119200 83426 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 4986 119200 5042 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 87694 119200 87750 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 92110 119200 92166 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 96434 119200 96490 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 100758 119200 100814 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 105174 119200 105230 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 109498 119200 109554 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 113914 119200 113970 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 118238 119200 118294 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 122562 119200 122618 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 126978 119200 127034 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9310 119200 9366 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 131302 119200 131358 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 135626 119200 135682 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 140042 119200 140098 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 144366 119200 144422 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 148690 119200 148746 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 153106 119200 153162 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 157430 119200 157486 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 161754 119200 161810 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 13726 119200 13782 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18050 119200 18106 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 22374 119200 22430 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 26790 119200 26846 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31114 119200 31170 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 39854 119200 39910 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2042 119200 2098 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 45650 119200 45706 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 49974 119200 50030 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 54298 119200 54354 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 58714 119200 58770 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 63038 119200 63094 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 67362 119200 67418 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 71778 119200 71834 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 76102 119200 76158 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 80518 119200 80574 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 84842 119200 84898 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6458 119200 6514 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 89166 119200 89222 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 93582 119200 93638 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 97906 119200 97962 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 102230 119200 102286 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 106646 119200 106702 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 110970 119200 111026 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 124034 119200 124090 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 128358 119200 128414 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 10782 119200 10838 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 137098 119200 137154 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 141422 119200 141478 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 145838 119200 145894 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 150162 119200 150218 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 154486 119200 154542 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 158902 119200 158958 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 163226 119200 163282 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15106 119200 15162 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 19522 119200 19578 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 23846 119200 23902 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 32586 119200 32642 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 36910 119200 36966 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 41234 119200 41290 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3514 119200 3570 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 47122 119200 47178 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 51446 119200 51502 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 64510 119200 64566 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 68834 119200 68890 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 73250 119200 73306 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 77574 119200 77630 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 81898 119200 81954 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 86314 119200 86370 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 90638 119200 90694 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 94962 119200 95018 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 99378 119200 99434 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 103702 119200 103758 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 108026 119200 108082 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 112442 119200 112498 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 116766 119200 116822 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 121090 119200 121146 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 125506 119200 125562 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 129830 119200 129886 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12254 119200 12310 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 134154 119200 134210 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 138570 119200 138626 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 142894 119200 142950 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 147310 119200 147366 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 151634 119200 151690 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 155958 119200 156014 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 160374 119200 160430 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 164698 119200 164754 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 16578 119200 16634 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 20902 119200 20958 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25318 119200 25374 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 29642 119200 29698 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 33966 119200 34022 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 38382 119200 38438 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 42706 119200 42762 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 160558 0 160614 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 165986 0 166042 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 167090 0 167146 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 171414 0 171470 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 user_clock2
port 529 nsew signal input
rlabel metal2 s 166170 119200 166226 120000 6 user_irq[0]
port 530 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 user_irq[1]
port 531 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7796784
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_7.magic.gds
string GDS_START 299924
<< end >>

