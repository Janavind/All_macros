magic
tech sky130A
magscale 1 2
timestamp 1653373056
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 14 2128 178848 117552
<< metal2 >>
rect 662 119200 718 120000
rect 1950 119200 2006 120000
rect 3238 119200 3294 120000
rect 4526 119200 4582 120000
rect 5814 119200 5870 120000
rect 7102 119200 7158 120000
rect 8482 119200 8538 120000
rect 9770 119200 9826 120000
rect 11058 119200 11114 120000
rect 12346 119200 12402 120000
rect 13634 119200 13690 120000
rect 14922 119200 14978 120000
rect 16302 119200 16358 120000
rect 17590 119200 17646 120000
rect 18878 119200 18934 120000
rect 20166 119200 20222 120000
rect 21454 119200 21510 120000
rect 22834 119200 22890 120000
rect 24122 119200 24178 120000
rect 25410 119200 25466 120000
rect 26698 119200 26754 120000
rect 27986 119200 28042 120000
rect 29274 119200 29330 120000
rect 30654 119200 30710 120000
rect 31942 119200 31998 120000
rect 33230 119200 33286 120000
rect 34518 119200 34574 120000
rect 35806 119200 35862 120000
rect 37186 119200 37242 120000
rect 38474 119200 38530 120000
rect 39762 119200 39818 120000
rect 41050 119200 41106 120000
rect 42338 119200 42394 120000
rect 43626 119200 43682 120000
rect 45006 119200 45062 120000
rect 46294 119200 46350 120000
rect 47582 119200 47638 120000
rect 48870 119200 48926 120000
rect 50158 119200 50214 120000
rect 51538 119200 51594 120000
rect 52826 119200 52882 120000
rect 54114 119200 54170 120000
rect 55402 119200 55458 120000
rect 56690 119200 56746 120000
rect 57978 119200 58034 120000
rect 59358 119200 59414 120000
rect 60646 119200 60702 120000
rect 61934 119200 61990 120000
rect 63222 119200 63278 120000
rect 64510 119200 64566 120000
rect 65890 119200 65946 120000
rect 67178 119200 67234 120000
rect 68466 119200 68522 120000
rect 69754 119200 69810 120000
rect 71042 119200 71098 120000
rect 72330 119200 72386 120000
rect 73710 119200 73766 120000
rect 74998 119200 75054 120000
rect 76286 119200 76342 120000
rect 77574 119200 77630 120000
rect 78862 119200 78918 120000
rect 80242 119200 80298 120000
rect 81530 119200 81586 120000
rect 82818 119200 82874 120000
rect 84106 119200 84162 120000
rect 85394 119200 85450 120000
rect 86682 119200 86738 120000
rect 88062 119200 88118 120000
rect 89350 119200 89406 120000
rect 90638 119200 90694 120000
rect 91926 119200 91982 120000
rect 93214 119200 93270 120000
rect 94594 119200 94650 120000
rect 95882 119200 95938 120000
rect 97170 119200 97226 120000
rect 98458 119200 98514 120000
rect 99746 119200 99802 120000
rect 101034 119200 101090 120000
rect 102414 119200 102470 120000
rect 103702 119200 103758 120000
rect 104990 119200 105046 120000
rect 106278 119200 106334 120000
rect 107566 119200 107622 120000
rect 108946 119200 109002 120000
rect 110234 119200 110290 120000
rect 111522 119200 111578 120000
rect 112810 119200 112866 120000
rect 114098 119200 114154 120000
rect 115386 119200 115442 120000
rect 116766 119200 116822 120000
rect 118054 119200 118110 120000
rect 119342 119200 119398 120000
rect 120630 119200 120686 120000
rect 121918 119200 121974 120000
rect 123298 119200 123354 120000
rect 124586 119200 124642 120000
rect 125874 119200 125930 120000
rect 127162 119200 127218 120000
rect 128450 119200 128506 120000
rect 129738 119200 129794 120000
rect 131118 119200 131174 120000
rect 132406 119200 132462 120000
rect 133694 119200 133750 120000
rect 134982 119200 135038 120000
rect 136270 119200 136326 120000
rect 137650 119200 137706 120000
rect 138938 119200 138994 120000
rect 140226 119200 140282 120000
rect 141514 119200 141570 120000
rect 142802 119200 142858 120000
rect 144090 119200 144146 120000
rect 145470 119200 145526 120000
rect 146758 119200 146814 120000
rect 148046 119200 148102 120000
rect 149334 119200 149390 120000
rect 150622 119200 150678 120000
rect 152002 119200 152058 120000
rect 153290 119200 153346 120000
rect 154578 119200 154634 120000
rect 155866 119200 155922 120000
rect 157154 119200 157210 120000
rect 158442 119200 158498 120000
rect 159822 119200 159878 120000
rect 161110 119200 161166 120000
rect 162398 119200 162454 120000
rect 163686 119200 163742 120000
rect 164974 119200 165030 120000
rect 166354 119200 166410 120000
rect 167642 119200 167698 120000
rect 168930 119200 168986 120000
rect 170218 119200 170274 120000
rect 171506 119200 171562 120000
rect 172794 119200 172850 120000
rect 174174 119200 174230 120000
rect 175462 119200 175518 120000
rect 176750 119200 176806 120000
rect 178038 119200 178094 120000
rect 179326 119200 179382 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59174 0 59230 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88522 0 88578 800
rect 88890 0 88946 800
rect 89258 0 89314 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91282 0 91338 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92386 0 92442 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 120998 0 121054 800
rect 121366 0 121422 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152462 0 152518 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157430 0 157486 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160190 0 160246 800
rect 160558 0 160614 800
rect 160926 0 160982 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161938 0 161994 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168194 0 168250 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173438 0 173494 800
rect 173806 0 173862 800
rect 174174 0 174230 800
rect 174542 0 174598 800
rect 174910 0 174966 800
rect 175186 0 175242 800
rect 175554 0 175610 800
rect 175922 0 175978 800
rect 176290 0 176346 800
rect 176658 0 176714 800
rect 176934 0 176990 800
rect 177302 0 177358 800
rect 177670 0 177726 800
rect 178038 0 178094 800
rect 178406 0 178462 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 20 119144 606 119354
rect 774 119144 1894 119354
rect 2062 119144 3182 119354
rect 3350 119144 4470 119354
rect 4638 119144 5758 119354
rect 5926 119144 7046 119354
rect 7214 119144 8426 119354
rect 8594 119144 9714 119354
rect 9882 119144 11002 119354
rect 11170 119144 12290 119354
rect 12458 119144 13578 119354
rect 13746 119144 14866 119354
rect 15034 119144 16246 119354
rect 16414 119144 17534 119354
rect 17702 119144 18822 119354
rect 18990 119144 20110 119354
rect 20278 119144 21398 119354
rect 21566 119144 22778 119354
rect 22946 119144 24066 119354
rect 24234 119144 25354 119354
rect 25522 119144 26642 119354
rect 26810 119144 27930 119354
rect 28098 119144 29218 119354
rect 29386 119144 30598 119354
rect 30766 119144 31886 119354
rect 32054 119144 33174 119354
rect 33342 119144 34462 119354
rect 34630 119144 35750 119354
rect 35918 119144 37130 119354
rect 37298 119144 38418 119354
rect 38586 119144 39706 119354
rect 39874 119144 40994 119354
rect 41162 119144 42282 119354
rect 42450 119144 43570 119354
rect 43738 119144 44950 119354
rect 45118 119144 46238 119354
rect 46406 119144 47526 119354
rect 47694 119144 48814 119354
rect 48982 119144 50102 119354
rect 50270 119144 51482 119354
rect 51650 119144 52770 119354
rect 52938 119144 54058 119354
rect 54226 119144 55346 119354
rect 55514 119144 56634 119354
rect 56802 119144 57922 119354
rect 58090 119144 59302 119354
rect 59470 119144 60590 119354
rect 60758 119144 61878 119354
rect 62046 119144 63166 119354
rect 63334 119144 64454 119354
rect 64622 119144 65834 119354
rect 66002 119144 67122 119354
rect 67290 119144 68410 119354
rect 68578 119144 69698 119354
rect 69866 119144 70986 119354
rect 71154 119144 72274 119354
rect 72442 119144 73654 119354
rect 73822 119144 74942 119354
rect 75110 119144 76230 119354
rect 76398 119144 77518 119354
rect 77686 119144 78806 119354
rect 78974 119144 80186 119354
rect 80354 119144 81474 119354
rect 81642 119144 82762 119354
rect 82930 119144 84050 119354
rect 84218 119144 85338 119354
rect 85506 119144 86626 119354
rect 86794 119144 88006 119354
rect 88174 119144 89294 119354
rect 89462 119144 90582 119354
rect 90750 119144 91870 119354
rect 92038 119144 93158 119354
rect 93326 119144 94538 119354
rect 94706 119144 95826 119354
rect 95994 119144 97114 119354
rect 97282 119144 98402 119354
rect 98570 119144 99690 119354
rect 99858 119144 100978 119354
rect 101146 119144 102358 119354
rect 102526 119144 103646 119354
rect 103814 119144 104934 119354
rect 105102 119144 106222 119354
rect 106390 119144 107510 119354
rect 107678 119144 108890 119354
rect 109058 119144 110178 119354
rect 110346 119144 111466 119354
rect 111634 119144 112754 119354
rect 112922 119144 114042 119354
rect 114210 119144 115330 119354
rect 115498 119144 116710 119354
rect 116878 119144 117998 119354
rect 118166 119144 119286 119354
rect 119454 119144 120574 119354
rect 120742 119144 121862 119354
rect 122030 119144 123242 119354
rect 123410 119144 124530 119354
rect 124698 119144 125818 119354
rect 125986 119144 127106 119354
rect 127274 119144 128394 119354
rect 128562 119144 129682 119354
rect 129850 119144 131062 119354
rect 131230 119144 132350 119354
rect 132518 119144 133638 119354
rect 133806 119144 134926 119354
rect 135094 119144 136214 119354
rect 136382 119144 137594 119354
rect 137762 119144 138882 119354
rect 139050 119144 140170 119354
rect 140338 119144 141458 119354
rect 141626 119144 142746 119354
rect 142914 119144 144034 119354
rect 144202 119144 145414 119354
rect 145582 119144 146702 119354
rect 146870 119144 147990 119354
rect 148158 119144 149278 119354
rect 149446 119144 150566 119354
rect 150734 119144 151946 119354
rect 152114 119144 153234 119354
rect 153402 119144 154522 119354
rect 154690 119144 155810 119354
rect 155978 119144 157098 119354
rect 157266 119144 158386 119354
rect 158554 119144 159766 119354
rect 159934 119144 161054 119354
rect 161222 119144 162342 119354
rect 162510 119144 163630 119354
rect 163798 119144 164918 119354
rect 165086 119144 166298 119354
rect 166466 119144 167586 119354
rect 167754 119144 168874 119354
rect 169042 119144 170162 119354
rect 170330 119144 171450 119354
rect 171618 119144 172738 119354
rect 172906 119144 174118 119354
rect 174286 119144 175406 119354
rect 175574 119144 176694 119354
rect 176862 119144 177982 119354
rect 178150 119144 178186 119354
rect 20 856 178186 119144
rect 20 800 54 856
rect 222 800 330 856
rect 498 800 698 856
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2446 856
rect 2614 800 2814 856
rect 2982 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3826 856
rect 3994 800 4194 856
rect 4362 800 4562 856
rect 4730 800 4930 856
rect 5098 800 5298 856
rect 5466 800 5574 856
rect 5742 800 5942 856
rect 6110 800 6310 856
rect 6478 800 6678 856
rect 6846 800 7046 856
rect 7214 800 7322 856
rect 7490 800 7690 856
rect 7858 800 8058 856
rect 8226 800 8426 856
rect 8594 800 8794 856
rect 8962 800 9070 856
rect 9238 800 9438 856
rect 9606 800 9806 856
rect 9974 800 10174 856
rect 10342 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13302 856
rect 13470 800 13670 856
rect 13838 800 14038 856
rect 14206 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15050 856
rect 15218 800 15418 856
rect 15586 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16430 856
rect 16598 800 16798 856
rect 16966 800 17166 856
rect 17334 800 17534 856
rect 17702 800 17810 856
rect 17978 800 18178 856
rect 18346 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19558 856
rect 19726 800 19926 856
rect 20094 800 20294 856
rect 20462 800 20662 856
rect 20830 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23422 856
rect 23590 800 23790 856
rect 23958 800 24158 856
rect 24326 800 24526 856
rect 24694 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25538 856
rect 25706 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26550 856
rect 26718 800 26918 856
rect 27086 800 27286 856
rect 27454 800 27654 856
rect 27822 800 28022 856
rect 28190 800 28298 856
rect 28466 800 28666 856
rect 28834 800 29034 856
rect 29202 800 29402 856
rect 29570 800 29770 856
rect 29938 800 30046 856
rect 30214 800 30414 856
rect 30582 800 30782 856
rect 30950 800 31150 856
rect 31318 800 31518 856
rect 31686 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34646 856
rect 34814 800 35014 856
rect 35182 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37038 856
rect 37206 800 37406 856
rect 37574 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38786 856
rect 38954 800 39154 856
rect 39322 800 39522 856
rect 39690 800 39890 856
rect 40058 800 40258 856
rect 40426 800 40534 856
rect 40702 800 40902 856
rect 41070 800 41270 856
rect 41438 800 41638 856
rect 41806 800 42006 856
rect 42174 800 42282 856
rect 42450 800 42650 856
rect 42818 800 43018 856
rect 43186 800 43386 856
rect 43554 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44398 856
rect 44566 800 44766 856
rect 44934 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45778 856
rect 45946 800 46146 856
rect 46314 800 46514 856
rect 46682 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47526 856
rect 47694 800 47894 856
rect 48062 800 48262 856
rect 48430 800 48630 856
rect 48798 800 48998 856
rect 49166 800 49274 856
rect 49442 800 49642 856
rect 49810 800 50010 856
rect 50178 800 50378 856
rect 50546 800 50746 856
rect 50914 800 51022 856
rect 51190 800 51390 856
rect 51558 800 51758 856
rect 51926 800 52126 856
rect 52294 800 52494 856
rect 52662 800 52770 856
rect 52938 800 53138 856
rect 53306 800 53506 856
rect 53674 800 53874 856
rect 54042 800 54242 856
rect 54410 800 54518 856
rect 54686 800 54886 856
rect 55054 800 55254 856
rect 55422 800 55622 856
rect 55790 800 55990 856
rect 56158 800 56266 856
rect 56434 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57738 856
rect 57906 800 58014 856
rect 58182 800 58382 856
rect 58550 800 58750 856
rect 58918 800 59118 856
rect 59286 800 59486 856
rect 59654 800 59762 856
rect 59930 800 60130 856
rect 60298 800 60498 856
rect 60666 800 60866 856
rect 61034 800 61234 856
rect 61402 800 61510 856
rect 61678 800 61878 856
rect 62046 800 62246 856
rect 62414 800 62614 856
rect 62782 800 62982 856
rect 63150 800 63258 856
rect 63426 800 63626 856
rect 63794 800 63994 856
rect 64162 800 64362 856
rect 64530 800 64730 856
rect 64898 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65742 856
rect 65910 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66754 856
rect 66922 800 67122 856
rect 67290 800 67490 856
rect 67658 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68502 856
rect 68670 800 68870 856
rect 69038 800 69238 856
rect 69406 800 69606 856
rect 69774 800 69974 856
rect 70142 800 70250 856
rect 70418 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71354 856
rect 71522 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73746 856
rect 73914 800 74114 856
rect 74282 800 74482 856
rect 74650 800 74850 856
rect 75018 800 75218 856
rect 75386 800 75494 856
rect 75662 800 75862 856
rect 76030 800 76230 856
rect 76398 800 76598 856
rect 76766 800 76966 856
rect 77134 800 77242 856
rect 77410 800 77610 856
rect 77778 800 77978 856
rect 78146 800 78346 856
rect 78514 800 78714 856
rect 78882 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79726 856
rect 79894 800 80094 856
rect 80262 800 80462 856
rect 80630 800 80738 856
rect 80906 800 81106 856
rect 81274 800 81474 856
rect 81642 800 81842 856
rect 82010 800 82210 856
rect 82378 800 82486 856
rect 82654 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83958 856
rect 84126 800 84234 856
rect 84402 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85338 856
rect 85506 800 85706 856
rect 85874 800 85982 856
rect 86150 800 86350 856
rect 86518 800 86718 856
rect 86886 800 87086 856
rect 87254 800 87454 856
rect 87622 800 87730 856
rect 87898 800 88098 856
rect 88266 800 88466 856
rect 88634 800 88834 856
rect 89002 800 89202 856
rect 89370 800 89478 856
rect 89646 800 89846 856
rect 90014 800 90214 856
rect 90382 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91226 856
rect 91394 800 91594 856
rect 91762 800 91962 856
rect 92130 800 92330 856
rect 92498 800 92698 856
rect 92866 800 92974 856
rect 93142 800 93342 856
rect 93510 800 93710 856
rect 93878 800 94078 856
rect 94246 800 94446 856
rect 94614 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97206 856
rect 97374 800 97574 856
rect 97742 800 97942 856
rect 98110 800 98218 856
rect 98386 800 98586 856
rect 98754 800 98954 856
rect 99122 800 99322 856
rect 99490 800 99690 856
rect 99858 800 99966 856
rect 100134 800 100334 856
rect 100502 800 100702 856
rect 100870 800 101070 856
rect 101238 800 101438 856
rect 101606 800 101714 856
rect 101882 800 102082 856
rect 102250 800 102450 856
rect 102618 800 102818 856
rect 102986 800 103186 856
rect 103354 800 103462 856
rect 103630 800 103830 856
rect 103998 800 104198 856
rect 104366 800 104566 856
rect 104734 800 104934 856
rect 105102 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105946 856
rect 106114 800 106314 856
rect 106482 800 106682 856
rect 106850 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107694 856
rect 107862 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108706 856
rect 108874 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110454 856
rect 110622 800 110822 856
rect 110990 800 111190 856
rect 111358 800 111558 856
rect 111726 800 111926 856
rect 112094 800 112202 856
rect 112370 800 112570 856
rect 112738 800 112938 856
rect 113106 800 113306 856
rect 113474 800 113674 856
rect 113842 800 113950 856
rect 114118 800 114318 856
rect 114486 800 114686 856
rect 114854 800 115054 856
rect 115222 800 115422 856
rect 115590 800 115698 856
rect 115866 800 116066 856
rect 116234 800 116434 856
rect 116602 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117446 856
rect 117614 800 117814 856
rect 117982 800 118182 856
rect 118350 800 118550 856
rect 118718 800 118918 856
rect 119086 800 119194 856
rect 119362 800 119562 856
rect 119730 800 119930 856
rect 120098 800 120298 856
rect 120466 800 120666 856
rect 120834 800 120942 856
rect 121110 800 121310 856
rect 121478 800 121678 856
rect 121846 800 122046 856
rect 122214 800 122414 856
rect 122582 800 122690 856
rect 122858 800 123058 856
rect 123226 800 123426 856
rect 123594 800 123794 856
rect 123962 800 124162 856
rect 124330 800 124438 856
rect 124606 800 124806 856
rect 124974 800 125174 856
rect 125342 800 125542 856
rect 125710 800 125910 856
rect 126078 800 126186 856
rect 126354 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127290 856
rect 127458 800 127658 856
rect 127826 800 127934 856
rect 128102 800 128302 856
rect 128470 800 128670 856
rect 128838 800 129038 856
rect 129206 800 129406 856
rect 129574 800 129682 856
rect 129850 800 130050 856
rect 130218 800 130418 856
rect 130586 800 130786 856
rect 130954 800 131154 856
rect 131322 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132166 856
rect 132334 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133178 856
rect 133346 800 133546 856
rect 133714 800 133914 856
rect 134082 800 134282 856
rect 134450 800 134650 856
rect 134818 800 134926 856
rect 135094 800 135294 856
rect 135462 800 135662 856
rect 135830 800 136030 856
rect 136198 800 136398 856
rect 136566 800 136674 856
rect 136842 800 137042 856
rect 137210 800 137410 856
rect 137578 800 137778 856
rect 137946 800 138146 856
rect 138314 800 138422 856
rect 138590 800 138790 856
rect 138958 800 139158 856
rect 139326 800 139526 856
rect 139694 800 139894 856
rect 140062 800 140170 856
rect 140338 800 140538 856
rect 140706 800 140906 856
rect 141074 800 141274 856
rect 141442 800 141642 856
rect 141810 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142654 856
rect 142822 800 143022 856
rect 143190 800 143390 856
rect 143558 800 143666 856
rect 143834 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145414 856
rect 145582 800 145782 856
rect 145950 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146886 856
rect 147054 800 147162 856
rect 147330 800 147530 856
rect 147698 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 148910 856
rect 149078 800 149278 856
rect 149446 800 149646 856
rect 149814 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150658 856
rect 150826 800 151026 856
rect 151194 800 151394 856
rect 151562 800 151762 856
rect 151930 800 152130 856
rect 152298 800 152406 856
rect 152574 800 152774 856
rect 152942 800 153142 856
rect 153310 800 153510 856
rect 153678 800 153878 856
rect 154046 800 154154 856
rect 154322 800 154522 856
rect 154690 800 154890 856
rect 155058 800 155258 856
rect 155426 800 155626 856
rect 155794 800 155902 856
rect 156070 800 156270 856
rect 156438 800 156638 856
rect 156806 800 157006 856
rect 157174 800 157374 856
rect 157542 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159398 856
rect 159566 800 159766 856
rect 159934 800 160134 856
rect 160302 800 160502 856
rect 160670 800 160870 856
rect 161038 800 161146 856
rect 161314 800 161514 856
rect 161682 800 161882 856
rect 162050 800 162250 856
rect 162418 800 162618 856
rect 162786 800 162894 856
rect 163062 800 163262 856
rect 163430 800 163630 856
rect 163798 800 163998 856
rect 164166 800 164366 856
rect 164534 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166390 856
rect 166558 800 166758 856
rect 166926 800 167126 856
rect 167294 800 167494 856
rect 167662 800 167862 856
rect 168030 800 168138 856
rect 168306 800 168506 856
rect 168674 800 168874 856
rect 169042 800 169242 856
rect 169410 800 169610 856
rect 169778 800 169886 856
rect 170054 800 170254 856
rect 170422 800 170622 856
rect 170790 800 170990 856
rect 171158 800 171358 856
rect 171526 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173106 856
rect 173274 800 173382 856
rect 173550 800 173750 856
rect 173918 800 174118 856
rect 174286 800 174486 856
rect 174654 800 174854 856
rect 175022 800 175130 856
rect 175298 800 175498 856
rect 175666 800 175866 856
rect 176034 800 176234 856
rect 176402 800 176602 856
rect 176770 800 176878 856
rect 177046 800 177246 856
rect 177414 800 177614 856
rect 177782 800 177982 856
rect 178150 800 178186 856
<< metal3 >>
rect 179200 117784 180000 117904
rect 0 116560 800 116680
rect 179200 113840 180000 113960
rect 0 109896 800 110016
rect 179200 109760 180000 109880
rect 179200 105816 180000 105936
rect 0 103232 800 103352
rect 179200 101872 180000 101992
rect 179200 97792 180000 97912
rect 0 96568 800 96688
rect 179200 93848 180000 93968
rect 0 89904 800 90024
rect 179200 89768 180000 89888
rect 179200 85824 180000 85944
rect 0 83240 800 83360
rect 179200 81880 180000 82000
rect 179200 77800 180000 77920
rect 0 76576 800 76696
rect 179200 73856 180000 73976
rect 0 69912 800 70032
rect 179200 69776 180000 69896
rect 179200 65832 180000 65952
rect 0 63248 800 63368
rect 179200 61888 180000 62008
rect 179200 57808 180000 57928
rect 0 56584 800 56704
rect 179200 53864 180000 53984
rect 0 49920 800 50040
rect 179200 49784 180000 49904
rect 179200 45840 180000 45960
rect 0 43256 800 43376
rect 179200 41896 180000 42016
rect 179200 37816 180000 37936
rect 0 36592 800 36712
rect 179200 33872 180000 33992
rect 0 29928 800 30048
rect 179200 29792 180000 29912
rect 179200 25848 180000 25968
rect 0 23264 800 23384
rect 179200 21904 180000 22024
rect 179200 17824 180000 17944
rect 0 16600 800 16720
rect 179200 13880 180000 14000
rect 0 9936 800 10056
rect 179200 9800 180000 9920
rect 179200 5856 180000 5976
rect 0 3272 800 3392
rect 179200 1912 180000 2032
<< obsm3 >>
rect 800 116760 179200 117537
rect 880 116480 179200 116760
rect 800 114040 179200 116480
rect 800 113760 179120 114040
rect 800 110096 179200 113760
rect 880 109960 179200 110096
rect 880 109816 179120 109960
rect 800 109680 179120 109816
rect 800 106016 179200 109680
rect 800 105736 179120 106016
rect 800 103432 179200 105736
rect 880 103152 179200 103432
rect 800 102072 179200 103152
rect 800 101792 179120 102072
rect 800 97992 179200 101792
rect 800 97712 179120 97992
rect 800 96768 179200 97712
rect 880 96488 179200 96768
rect 800 94048 179200 96488
rect 800 93768 179120 94048
rect 800 90104 179200 93768
rect 880 89968 179200 90104
rect 880 89824 179120 89968
rect 800 89688 179120 89824
rect 800 86024 179200 89688
rect 800 85744 179120 86024
rect 800 83440 179200 85744
rect 880 83160 179200 83440
rect 800 82080 179200 83160
rect 800 81800 179120 82080
rect 800 78000 179200 81800
rect 800 77720 179120 78000
rect 800 76776 179200 77720
rect 880 76496 179200 76776
rect 800 74056 179200 76496
rect 800 73776 179120 74056
rect 800 70112 179200 73776
rect 880 69976 179200 70112
rect 880 69832 179120 69976
rect 800 69696 179120 69832
rect 800 66032 179200 69696
rect 800 65752 179120 66032
rect 800 63448 179200 65752
rect 880 63168 179200 63448
rect 800 62088 179200 63168
rect 800 61808 179120 62088
rect 800 58008 179200 61808
rect 800 57728 179120 58008
rect 800 56784 179200 57728
rect 880 56504 179200 56784
rect 800 54064 179200 56504
rect 800 53784 179120 54064
rect 800 50120 179200 53784
rect 880 49984 179200 50120
rect 880 49840 179120 49984
rect 800 49704 179120 49840
rect 800 46040 179200 49704
rect 800 45760 179120 46040
rect 800 43456 179200 45760
rect 880 43176 179200 43456
rect 800 42096 179200 43176
rect 800 41816 179120 42096
rect 800 38016 179200 41816
rect 800 37736 179120 38016
rect 800 36792 179200 37736
rect 880 36512 179200 36792
rect 800 34072 179200 36512
rect 800 33792 179120 34072
rect 800 30128 179200 33792
rect 880 29992 179200 30128
rect 880 29848 179120 29992
rect 800 29712 179120 29848
rect 800 26048 179200 29712
rect 800 25768 179120 26048
rect 800 23464 179200 25768
rect 880 23184 179200 23464
rect 800 22104 179200 23184
rect 800 21824 179120 22104
rect 800 18024 179200 21824
rect 800 17744 179120 18024
rect 800 16800 179200 17744
rect 880 16520 179200 16800
rect 800 14080 179200 16520
rect 800 13800 179120 14080
rect 800 10136 179200 13800
rect 880 10000 179200 10136
rect 880 9856 179120 10000
rect 800 9720 179120 9856
rect 800 6056 179200 9720
rect 800 5776 179120 6056
rect 800 3472 179200 5776
rect 880 3192 179200 3472
rect 800 2112 179200 3192
rect 800 1939 179120 2112
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 74395 4523 80928 117197
rect 81408 4523 96288 117197
rect 96768 4523 104821 117197
<< labels >>
rlabel metal3 s 179200 9800 180000 9920 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 179200 25848 180000 25968 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 179200 61888 180000 62008 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 A1[0]
port 9 nsew signal input
rlabel metal2 s 157154 119200 157210 120000 6 A1[1]
port 10 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 A1[2]
port 11 nsew signal input
rlabel metal3 s 179200 45840 180000 45960 6 A1[3]
port 12 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 A1[4]
port 13 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 A1[5]
port 14 nsew signal input
rlabel metal3 s 179200 73856 180000 73976 6 A1[6]
port 15 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 A1[7]
port 16 nsew signal input
rlabel metal2 s 150622 119200 150678 120000 6 ALU_Out1[0]
port 17 nsew signal output
rlabel metal2 s 158442 119200 158498 120000 6 ALU_Out1[1]
port 18 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 ALU_Out1[2]
port 19 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 ALU_Out1[3]
port 20 nsew signal output
rlabel metal3 s 179200 57808 180000 57928 6 ALU_Out1[4]
port 21 nsew signal output
rlabel metal3 s 179200 65832 180000 65952 6 ALU_Out1[5]
port 22 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 ALU_Out1[6]
port 23 nsew signal output
rlabel metal3 s 179200 89768 180000 89888 6 ALU_Out1[7]
port 24 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 ALU_Out2[0]
port 25 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 ALU_Out2[1]
port 26 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 ALU_Out2[2]
port 27 nsew signal output
rlabel metal3 s 179200 49784 180000 49904 6 ALU_Out2[3]
port 28 nsew signal output
rlabel metal2 s 164974 119200 165030 120000 6 ALU_Out2[4]
port 29 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 ALU_Out2[5]
port 30 nsew signal output
rlabel metal3 s 179200 77800 180000 77920 6 ALU_Out2[6]
port 31 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 ALU_Out2[7]
port 32 nsew signal output
rlabel metal2 s 152002 119200 152058 120000 6 ALU_Sel1[0]
port 33 nsew signal input
rlabel metal2 s 159822 119200 159878 120000 6 ALU_Sel1[1]
port 34 nsew signal input
rlabel metal3 s 179200 13880 180000 14000 6 ALU_Sel2[0]
port 35 nsew signal input
rlabel metal3 s 179200 17824 180000 17944 6 ALU_Sel2[1]
port 36 nsew signal input
rlabel metal2 s 153290 119200 153346 120000 6 B0[0]
port 37 nsew signal input
rlabel metal2 s 161110 119200 161166 120000 6 B0[1]
port 38 nsew signal input
rlabel metal3 s 179200 29792 180000 29912 6 B0[2]
port 39 nsew signal input
rlabel metal3 s 179200 53864 180000 53984 6 B0[3]
port 40 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 B0[4]
port 41 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 B0[5]
port 42 nsew signal input
rlabel metal3 s 179200 81880 180000 82000 6 B0[6]
port 43 nsew signal input
rlabel metal3 s 179200 93848 180000 93968 6 B0[7]
port 44 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 B1[0]
port 45 nsew signal input
rlabel metal3 s 179200 21904 180000 22024 6 B1[1]
port 46 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 B1[2]
port 47 nsew signal input
rlabel metal2 s 163686 119200 163742 120000 6 B1[3]
port 48 nsew signal input
rlabel metal2 s 166354 119200 166410 120000 6 B1[4]
port 49 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 B1[5]
port 50 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 B1[6]
port 51 nsew signal input
rlabel metal3 s 179200 97792 180000 97912 6 B1[7]
port 52 nsew signal input
rlabel metal3 s 179200 1912 180000 2032 6 CarryOut1
port 53 nsew signal output
rlabel metal2 s 171414 0 171470 800 6 CarryOut2
port 54 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 analog_io[0]
port 55 nsew signal bidirectional
rlabel metal3 s 179200 101872 180000 101992 6 analog_io[10]
port 56 nsew signal bidirectional
rlabel metal2 s 174174 119200 174230 120000 6 analog_io[11]
port 57 nsew signal bidirectional
rlabel metal3 s 179200 105816 180000 105936 6 analog_io[12]
port 58 nsew signal bidirectional
rlabel metal2 s 175462 119200 175518 120000 6 analog_io[13]
port 59 nsew signal bidirectional
rlabel metal2 s 178038 0 178094 800 6 analog_io[14]
port 60 nsew signal bidirectional
rlabel metal3 s 0 103232 800 103352 6 analog_io[15]
port 61 nsew signal bidirectional
rlabel metal2 s 176750 119200 176806 120000 6 analog_io[16]
port 62 nsew signal bidirectional
rlabel metal3 s 179200 109760 180000 109880 6 analog_io[17]
port 63 nsew signal bidirectional
rlabel metal2 s 178038 119200 178094 120000 6 analog_io[18]
port 64 nsew signal bidirectional
rlabel metal3 s 0 109896 800 110016 6 analog_io[19]
port 65 nsew signal bidirectional
rlabel metal2 s 162398 119200 162454 120000 6 analog_io[1]
port 66 nsew signal bidirectional
rlabel metal3 s 0 116560 800 116680 6 analog_io[20]
port 67 nsew signal bidirectional
rlabel metal2 s 178406 0 178462 800 6 analog_io[21]
port 68 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[22]
port 69 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[23]
port 70 nsew signal bidirectional
rlabel metal3 s 179200 113840 180000 113960 6 analog_io[24]
port 71 nsew signal bidirectional
rlabel metal2 s 179326 119200 179382 120000 6 analog_io[25]
port 72 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[26]
port 73 nsew signal bidirectional
rlabel metal3 s 179200 117784 180000 117904 6 analog_io[27]
port 74 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 75 nsew signal bidirectional
rlabel metal3 s 179200 33872 180000 33992 6 analog_io[2]
port 76 nsew signal bidirectional
rlabel metal3 s 0 56584 800 56704 6 analog_io[3]
port 77 nsew signal bidirectional
rlabel metal2 s 167642 119200 167698 120000 6 analog_io[4]
port 78 nsew signal bidirectional
rlabel metal2 s 168930 119200 168986 120000 6 analog_io[5]
port 79 nsew signal bidirectional
rlabel metal2 s 176934 0 176990 800 6 analog_io[6]
port 80 nsew signal bidirectional
rlabel metal2 s 170218 119200 170274 120000 6 analog_io[7]
port 81 nsew signal bidirectional
rlabel metal2 s 171506 119200 171562 120000 6 analog_io[8]
port 82 nsew signal bidirectional
rlabel metal2 s 172794 119200 172850 120000 6 analog_io[9]
port 83 nsew signal bidirectional
rlabel metal2 s 149334 119200 149390 120000 6 clk
port 84 nsew signal input
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 85 nsew signal input
rlabel metal2 s 39762 119200 39818 120000 6 io_in[10]
port 86 nsew signal input
rlabel metal2 s 43626 119200 43682 120000 6 io_in[11]
port 87 nsew signal input
rlabel metal2 s 47582 119200 47638 120000 6 io_in[12]
port 88 nsew signal input
rlabel metal2 s 51538 119200 51594 120000 6 io_in[13]
port 89 nsew signal input
rlabel metal2 s 55402 119200 55458 120000 6 io_in[14]
port 90 nsew signal input
rlabel metal2 s 59358 119200 59414 120000 6 io_in[15]
port 91 nsew signal input
rlabel metal2 s 63222 119200 63278 120000 6 io_in[16]
port 92 nsew signal input
rlabel metal2 s 67178 119200 67234 120000 6 io_in[17]
port 93 nsew signal input
rlabel metal2 s 71042 119200 71098 120000 6 io_in[18]
port 94 nsew signal input
rlabel metal2 s 74998 119200 75054 120000 6 io_in[19]
port 95 nsew signal input
rlabel metal2 s 4526 119200 4582 120000 6 io_in[1]
port 96 nsew signal input
rlabel metal2 s 78862 119200 78918 120000 6 io_in[20]
port 97 nsew signal input
rlabel metal2 s 82818 119200 82874 120000 6 io_in[21]
port 98 nsew signal input
rlabel metal2 s 86682 119200 86738 120000 6 io_in[22]
port 99 nsew signal input
rlabel metal2 s 90638 119200 90694 120000 6 io_in[23]
port 100 nsew signal input
rlabel metal2 s 94594 119200 94650 120000 6 io_in[24]
port 101 nsew signal input
rlabel metal2 s 98458 119200 98514 120000 6 io_in[25]
port 102 nsew signal input
rlabel metal2 s 102414 119200 102470 120000 6 io_in[26]
port 103 nsew signal input
rlabel metal2 s 106278 119200 106334 120000 6 io_in[27]
port 104 nsew signal input
rlabel metal2 s 110234 119200 110290 120000 6 io_in[28]
port 105 nsew signal input
rlabel metal2 s 114098 119200 114154 120000 6 io_in[29]
port 106 nsew signal input
rlabel metal2 s 8482 119200 8538 120000 6 io_in[2]
port 107 nsew signal input
rlabel metal2 s 118054 119200 118110 120000 6 io_in[30]
port 108 nsew signal input
rlabel metal2 s 121918 119200 121974 120000 6 io_in[31]
port 109 nsew signal input
rlabel metal2 s 125874 119200 125930 120000 6 io_in[32]
port 110 nsew signal input
rlabel metal2 s 129738 119200 129794 120000 6 io_in[33]
port 111 nsew signal input
rlabel metal2 s 133694 119200 133750 120000 6 io_in[34]
port 112 nsew signal input
rlabel metal2 s 137650 119200 137706 120000 6 io_in[35]
port 113 nsew signal input
rlabel metal2 s 141514 119200 141570 120000 6 io_in[36]
port 114 nsew signal input
rlabel metal2 s 145470 119200 145526 120000 6 io_in[37]
port 115 nsew signal input
rlabel metal2 s 12346 119200 12402 120000 6 io_in[3]
port 116 nsew signal input
rlabel metal2 s 16302 119200 16358 120000 6 io_in[4]
port 117 nsew signal input
rlabel metal2 s 20166 119200 20222 120000 6 io_in[5]
port 118 nsew signal input
rlabel metal2 s 24122 119200 24178 120000 6 io_in[6]
port 119 nsew signal input
rlabel metal2 s 27986 119200 28042 120000 6 io_in[7]
port 120 nsew signal input
rlabel metal2 s 31942 119200 31998 120000 6 io_in[8]
port 121 nsew signal input
rlabel metal2 s 35806 119200 35862 120000 6 io_in[9]
port 122 nsew signal input
rlabel metal2 s 1950 119200 2006 120000 6 io_oeb[0]
port 123 nsew signal output
rlabel metal2 s 41050 119200 41106 120000 6 io_oeb[10]
port 124 nsew signal output
rlabel metal2 s 45006 119200 45062 120000 6 io_oeb[11]
port 125 nsew signal output
rlabel metal2 s 48870 119200 48926 120000 6 io_oeb[12]
port 126 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_oeb[13]
port 127 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 io_oeb[14]
port 128 nsew signal output
rlabel metal2 s 60646 119200 60702 120000 6 io_oeb[15]
port 129 nsew signal output
rlabel metal2 s 64510 119200 64566 120000 6 io_oeb[16]
port 130 nsew signal output
rlabel metal2 s 68466 119200 68522 120000 6 io_oeb[17]
port 131 nsew signal output
rlabel metal2 s 72330 119200 72386 120000 6 io_oeb[18]
port 132 nsew signal output
rlabel metal2 s 76286 119200 76342 120000 6 io_oeb[19]
port 133 nsew signal output
rlabel metal2 s 5814 119200 5870 120000 6 io_oeb[1]
port 134 nsew signal output
rlabel metal2 s 80242 119200 80298 120000 6 io_oeb[20]
port 135 nsew signal output
rlabel metal2 s 84106 119200 84162 120000 6 io_oeb[21]
port 136 nsew signal output
rlabel metal2 s 88062 119200 88118 120000 6 io_oeb[22]
port 137 nsew signal output
rlabel metal2 s 91926 119200 91982 120000 6 io_oeb[23]
port 138 nsew signal output
rlabel metal2 s 95882 119200 95938 120000 6 io_oeb[24]
port 139 nsew signal output
rlabel metal2 s 99746 119200 99802 120000 6 io_oeb[25]
port 140 nsew signal output
rlabel metal2 s 103702 119200 103758 120000 6 io_oeb[26]
port 141 nsew signal output
rlabel metal2 s 107566 119200 107622 120000 6 io_oeb[27]
port 142 nsew signal output
rlabel metal2 s 111522 119200 111578 120000 6 io_oeb[28]
port 143 nsew signal output
rlabel metal2 s 115386 119200 115442 120000 6 io_oeb[29]
port 144 nsew signal output
rlabel metal2 s 9770 119200 9826 120000 6 io_oeb[2]
port 145 nsew signal output
rlabel metal2 s 119342 119200 119398 120000 6 io_oeb[30]
port 146 nsew signal output
rlabel metal2 s 123298 119200 123354 120000 6 io_oeb[31]
port 147 nsew signal output
rlabel metal2 s 127162 119200 127218 120000 6 io_oeb[32]
port 148 nsew signal output
rlabel metal2 s 131118 119200 131174 120000 6 io_oeb[33]
port 149 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[34]
port 150 nsew signal output
rlabel metal2 s 138938 119200 138994 120000 6 io_oeb[35]
port 151 nsew signal output
rlabel metal2 s 142802 119200 142858 120000 6 io_oeb[36]
port 152 nsew signal output
rlabel metal2 s 146758 119200 146814 120000 6 io_oeb[37]
port 153 nsew signal output
rlabel metal2 s 13634 119200 13690 120000 6 io_oeb[3]
port 154 nsew signal output
rlabel metal2 s 17590 119200 17646 120000 6 io_oeb[4]
port 155 nsew signal output
rlabel metal2 s 21454 119200 21510 120000 6 io_oeb[5]
port 156 nsew signal output
rlabel metal2 s 25410 119200 25466 120000 6 io_oeb[6]
port 157 nsew signal output
rlabel metal2 s 29274 119200 29330 120000 6 io_oeb[7]
port 158 nsew signal output
rlabel metal2 s 33230 119200 33286 120000 6 io_oeb[8]
port 159 nsew signal output
rlabel metal2 s 37186 119200 37242 120000 6 io_oeb[9]
port 160 nsew signal output
rlabel metal2 s 3238 119200 3294 120000 6 io_out[0]
port 161 nsew signal output
rlabel metal2 s 42338 119200 42394 120000 6 io_out[10]
port 162 nsew signal output
rlabel metal2 s 46294 119200 46350 120000 6 io_out[11]
port 163 nsew signal output
rlabel metal2 s 50158 119200 50214 120000 6 io_out[12]
port 164 nsew signal output
rlabel metal2 s 54114 119200 54170 120000 6 io_out[13]
port 165 nsew signal output
rlabel metal2 s 57978 119200 58034 120000 6 io_out[14]
port 166 nsew signal output
rlabel metal2 s 61934 119200 61990 120000 6 io_out[15]
port 167 nsew signal output
rlabel metal2 s 65890 119200 65946 120000 6 io_out[16]
port 168 nsew signal output
rlabel metal2 s 69754 119200 69810 120000 6 io_out[17]
port 169 nsew signal output
rlabel metal2 s 73710 119200 73766 120000 6 io_out[18]
port 170 nsew signal output
rlabel metal2 s 77574 119200 77630 120000 6 io_out[19]
port 171 nsew signal output
rlabel metal2 s 7102 119200 7158 120000 6 io_out[1]
port 172 nsew signal output
rlabel metal2 s 81530 119200 81586 120000 6 io_out[20]
port 173 nsew signal output
rlabel metal2 s 85394 119200 85450 120000 6 io_out[21]
port 174 nsew signal output
rlabel metal2 s 89350 119200 89406 120000 6 io_out[22]
port 175 nsew signal output
rlabel metal2 s 93214 119200 93270 120000 6 io_out[23]
port 176 nsew signal output
rlabel metal2 s 97170 119200 97226 120000 6 io_out[24]
port 177 nsew signal output
rlabel metal2 s 101034 119200 101090 120000 6 io_out[25]
port 178 nsew signal output
rlabel metal2 s 104990 119200 105046 120000 6 io_out[26]
port 179 nsew signal output
rlabel metal2 s 108946 119200 109002 120000 6 io_out[27]
port 180 nsew signal output
rlabel metal2 s 112810 119200 112866 120000 6 io_out[28]
port 181 nsew signal output
rlabel metal2 s 116766 119200 116822 120000 6 io_out[29]
port 182 nsew signal output
rlabel metal2 s 11058 119200 11114 120000 6 io_out[2]
port 183 nsew signal output
rlabel metal2 s 120630 119200 120686 120000 6 io_out[30]
port 184 nsew signal output
rlabel metal2 s 124586 119200 124642 120000 6 io_out[31]
port 185 nsew signal output
rlabel metal2 s 128450 119200 128506 120000 6 io_out[32]
port 186 nsew signal output
rlabel metal2 s 132406 119200 132462 120000 6 io_out[33]
port 187 nsew signal output
rlabel metal2 s 136270 119200 136326 120000 6 io_out[34]
port 188 nsew signal output
rlabel metal2 s 140226 119200 140282 120000 6 io_out[35]
port 189 nsew signal output
rlabel metal2 s 144090 119200 144146 120000 6 io_out[36]
port 190 nsew signal output
rlabel metal2 s 148046 119200 148102 120000 6 io_out[37]
port 191 nsew signal output
rlabel metal2 s 14922 119200 14978 120000 6 io_out[3]
port 192 nsew signal output
rlabel metal2 s 18878 119200 18934 120000 6 io_out[4]
port 193 nsew signal output
rlabel metal2 s 22834 119200 22890 120000 6 io_out[5]
port 194 nsew signal output
rlabel metal2 s 26698 119200 26754 120000 6 io_out[6]
port 195 nsew signal output
rlabel metal2 s 30654 119200 30710 120000 6 io_out[7]
port 196 nsew signal output
rlabel metal2 s 34518 119200 34574 120000 6 io_out[8]
port 197 nsew signal output
rlabel metal2 s 38474 119200 38530 120000 6 io_out[9]
port 198 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_in[0]
port 199 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[100]
port 200 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[101]
port 201 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[102]
port 202 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[103]
port 203 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[104]
port 204 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[105]
port 205 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[106]
port 206 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[107]
port 207 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[108]
port 208 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[109]
port 209 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[10]
port 210 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[110]
port 211 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[111]
port 212 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[112]
port 213 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[113]
port 214 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[114]
port 215 nsew signal input
rlabel metal2 s 157706 0 157762 800 6 la_data_in[115]
port 216 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 la_data_in[116]
port 217 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[117]
port 218 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[118]
port 219 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[119]
port 220 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[11]
port 221 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_data_in[120]
port 222 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_data_in[121]
port 223 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[122]
port 224 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[123]
port 225 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[124]
port 226 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_data_in[125]
port 227 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_data_in[126]
port 228 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[127]
port 229 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[12]
port 230 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[13]
port 231 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[14]
port 232 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[15]
port 233 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[16]
port 234 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[17]
port 235 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[18]
port 236 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[19]
port 237 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_data_in[1]
port 238 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[20]
port 239 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_data_in[21]
port 240 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[22]
port 241 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[23]
port 242 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[24]
port 243 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[25]
port 244 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_data_in[26]
port 245 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[27]
port 246 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[28]
port 247 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[29]
port 248 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[2]
port 249 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[30]
port 250 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[31]
port 251 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[32]
port 252 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[33]
port 253 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[34]
port 254 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[35]
port 255 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[36]
port 256 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[37]
port 257 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[38]
port 258 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[39]
port 259 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[3]
port 260 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[40]
port 261 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[41]
port 262 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[42]
port 263 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[43]
port 264 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[44]
port 265 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[45]
port 266 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[46]
port 267 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[47]
port 268 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[48]
port 269 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[49]
port 270 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[4]
port 271 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_data_in[50]
port 272 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[51]
port 273 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[52]
port 274 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[53]
port 275 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 la_data_in[54]
port 276 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[55]
port 277 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[56]
port 278 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[57]
port 279 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[58]
port 280 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[59]
port 281 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[5]
port 282 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[60]
port 283 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[61]
port 284 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[62]
port 285 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[63]
port 286 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[64]
port 287 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[65]
port 288 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_data_in[66]
port 289 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[67]
port 290 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[68]
port 291 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[69]
port 292 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[6]
port 293 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_data_in[70]
port 294 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_data_in[71]
port 295 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[72]
port 296 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[73]
port 297 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[74]
port 298 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[75]
port 299 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[76]
port 300 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_data_in[77]
port 301 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[78]
port 302 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[79]
port 303 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[7]
port 304 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_data_in[80]
port 305 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[81]
port 306 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[82]
port 307 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[83]
port 308 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[84]
port 309 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[85]
port 310 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[86]
port 311 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[87]
port 312 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[88]
port 313 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[89]
port 314 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[8]
port 315 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[90]
port 316 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[91]
port 317 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[92]
port 318 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[93]
port 319 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[94]
port 320 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[95]
port 321 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[96]
port 322 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[97]
port 323 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[98]
port 324 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_data_in[99]
port 325 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[9]
port 326 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_out[0]
port 327 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[100]
port 328 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[101]
port 329 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[102]
port 330 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[103]
port 331 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[104]
port 332 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[105]
port 333 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[106]
port 334 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[107]
port 335 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[108]
port 336 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[109]
port 337 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[10]
port 338 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[110]
port 339 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[111]
port 340 nsew signal output
rlabel metal2 s 154946 0 155002 800 6 la_data_out[112]
port 341 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[113]
port 342 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[114]
port 343 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[115]
port 344 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[116]
port 345 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[117]
port 346 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[118]
port 347 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[119]
port 348 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[11]
port 349 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 la_data_out[120]
port 350 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[121]
port 351 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[122]
port 352 nsew signal output
rlabel metal2 s 166446 0 166502 800 6 la_data_out[123]
port 353 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 la_data_out[124]
port 354 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 la_data_out[125]
port 355 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 la_data_out[126]
port 356 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[127]
port 357 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[12]
port 358 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[13]
port 359 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[14]
port 360 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[15]
port 361 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[16]
port 362 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[17]
port 363 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[18]
port 364 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[19]
port 365 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[1]
port 366 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[20]
port 367 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[21]
port 368 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[22]
port 369 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[23]
port 370 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[24]
port 371 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[25]
port 372 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 la_data_out[26]
port 373 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[27]
port 374 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[28]
port 375 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[29]
port 376 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[2]
port 377 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[30]
port 378 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[31]
port 379 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[32]
port 380 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[33]
port 381 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[34]
port 382 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[35]
port 383 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[36]
port 384 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[37]
port 385 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[38]
port 386 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[39]
port 387 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[3]
port 388 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[40]
port 389 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[41]
port 390 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[42]
port 391 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[43]
port 392 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[44]
port 393 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[45]
port 394 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[46]
port 395 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[47]
port 396 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 la_data_out[48]
port 397 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 la_data_out[49]
port 398 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[4]
port 399 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[50]
port 400 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[51]
port 401 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[52]
port 402 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[53]
port 403 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[54]
port 404 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[55]
port 405 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[56]
port 406 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[57]
port 407 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[58]
port 408 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[59]
port 409 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[5]
port 410 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[60]
port 411 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[61]
port 412 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[62]
port 413 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[63]
port 414 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[64]
port 415 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[65]
port 416 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[66]
port 417 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[67]
port 418 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[68]
port 419 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[69]
port 420 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[6]
port 421 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[70]
port 422 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[71]
port 423 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[72]
port 424 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[73]
port 425 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[74]
port 426 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[75]
port 427 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[76]
port 428 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[77]
port 429 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[78]
port 430 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 la_data_out[79]
port 431 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[7]
port 432 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[80]
port 433 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 la_data_out[81]
port 434 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 la_data_out[82]
port 435 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 la_data_out[83]
port 436 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[84]
port 437 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[85]
port 438 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[86]
port 439 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[87]
port 440 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[88]
port 441 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[89]
port 442 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[8]
port 443 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[90]
port 444 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[91]
port 445 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[92]
port 446 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[93]
port 447 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[94]
port 448 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[95]
port 449 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[96]
port 450 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[97]
port 451 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[98]
port 452 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[99]
port 453 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[9]
port 454 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_oenb[0]
port 455 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[100]
port 456 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[101]
port 457 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[102]
port 458 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[103]
port 459 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oenb[104]
port 460 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[105]
port 461 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[106]
port 462 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_oenb[107]
port 463 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[108]
port 464 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_oenb[109]
port 465 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[10]
port 466 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[110]
port 467 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[111]
port 468 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[112]
port 469 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_oenb[113]
port 470 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oenb[114]
port 471 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[115]
port 472 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_oenb[116]
port 473 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[117]
port 474 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[118]
port 475 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[119]
port 476 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[11]
port 477 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_oenb[120]
port 478 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_oenb[121]
port 479 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[122]
port 480 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_oenb[123]
port 481 nsew signal input
rlabel metal2 s 167918 0 167974 800 6 la_oenb[124]
port 482 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[125]
port 483 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oenb[126]
port 484 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oenb[127]
port 485 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[12]
port 486 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[13]
port 487 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[14]
port 488 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[15]
port 489 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[16]
port 490 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[17]
port 491 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[18]
port 492 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[19]
port 493 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_oenb[1]
port 494 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[20]
port 495 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[21]
port 496 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_oenb[22]
port 497 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[23]
port 498 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[24]
port 499 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[25]
port 500 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_oenb[26]
port 501 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[27]
port 502 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[28]
port 503 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[29]
port 504 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[2]
port 505 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[30]
port 506 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[31]
port 507 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[32]
port 508 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[33]
port 509 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[34]
port 510 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[35]
port 511 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[36]
port 512 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[37]
port 513 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[38]
port 514 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[39]
port 515 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[3]
port 516 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[40]
port 517 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[41]
port 518 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[42]
port 519 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[43]
port 520 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[44]
port 521 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[45]
port 522 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[46]
port 523 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[47]
port 524 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[48]
port 525 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[49]
port 526 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[4]
port 527 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[50]
port 528 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[51]
port 529 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[52]
port 530 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[53]
port 531 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[54]
port 532 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[55]
port 533 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[56]
port 534 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[57]
port 535 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[58]
port 536 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[59]
port 537 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[5]
port 538 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[60]
port 539 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[61]
port 540 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[62]
port 541 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[63]
port 542 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[64]
port 543 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_oenb[65]
port 544 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[66]
port 545 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[67]
port 546 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[68]
port 547 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[69]
port 548 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[6]
port 549 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_oenb[70]
port 550 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[71]
port 551 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[72]
port 552 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_oenb[73]
port 553 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[74]
port 554 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[75]
port 555 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[76]
port 556 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[77]
port 557 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[78]
port 558 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[79]
port 559 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[7]
port 560 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[80]
port 561 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[81]
port 562 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[82]
port 563 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[83]
port 564 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_oenb[84]
port 565 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[85]
port 566 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[86]
port 567 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[87]
port 568 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oenb[88]
port 569 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[89]
port 570 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_oenb[8]
port 571 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_oenb[90]
port 572 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_oenb[91]
port 573 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[92]
port 574 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[93]
port 575 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[94]
port 576 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[95]
port 577 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[96]
port 578 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[97]
port 579 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[98]
port 580 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[99]
port 581 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[9]
port 582 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 user_clock2
port 583 nsew signal input
rlabel metal2 s 154578 119200 154634 120000 6 user_irq[0]
port 584 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 user_irq[1]
port 585 nsew signal output
rlabel metal3 s 179200 37816 180000 37936 6 user_irq[2]
port 586 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 587 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 588 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 588 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 588 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 588 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 588 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 588 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 589 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 590 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 591 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[0]
port 592 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[10]
port 593 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[11]
port 594 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[12]
port 595 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[13]
port 596 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[14]
port 597 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[15]
port 598 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[16]
port 599 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[17]
port 600 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_adr_i[18]
port 601 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[19]
port 602 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[1]
port 603 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[20]
port 604 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[21]
port 605 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[22]
port 606 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[23]
port 607 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[24]
port 608 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[25]
port 609 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[26]
port 610 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[27]
port 611 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[28]
port 612 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[29]
port 613 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_adr_i[2]
port 614 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_adr_i[30]
port 615 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[31]
port 616 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[3]
port 617 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_adr_i[4]
port 618 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_adr_i[5]
port 619 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[6]
port 620 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[7]
port 621 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[8]
port 622 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[9]
port 623 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 624 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_i[0]
port 625 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[10]
port 626 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_i[11]
port 627 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[12]
port 628 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[13]
port 629 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[14]
port 630 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[15]
port 631 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_i[16]
port 632 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[17]
port 633 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[18]
port 634 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[19]
port 635 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[1]
port 636 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[20]
port 637 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[21]
port 638 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[22]
port 639 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[23]
port 640 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[24]
port 641 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[25]
port 642 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[26]
port 643 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[27]
port 644 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[28]
port 645 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[29]
port 646 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[2]
port 647 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[30]
port 648 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[31]
port 649 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[3]
port 650 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[4]
port 651 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[5]
port 652 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[6]
port 653 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_i[7]
port 654 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[8]
port 655 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[9]
port 656 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_o[0]
port 657 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_o[10]
port 658 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[11]
port 659 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[12]
port 660 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[13]
port 661 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[14]
port 662 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[15]
port 663 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[16]
port 664 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[17]
port 665 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[18]
port 666 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[19]
port 667 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[1]
port 668 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[20]
port 669 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[21]
port 670 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[22]
port 671 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[23]
port 672 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[24]
port 673 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[25]
port 674 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_o[26]
port 675 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[27]
port 676 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[28]
port 677 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[29]
port 678 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[2]
port 679 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[30]
port 680 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[31]
port 681 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_o[3]
port 682 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[4]
port 683 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[5]
port 684 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[6]
port 685 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_o[7]
port 686 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[8]
port 687 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[9]
port 688 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[0]
port 689 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_sel_i[1]
port 690 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_sel_i[2]
port 691 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_sel_i[3]
port 692 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 693 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 694 nsew signal input
rlabel metal2 s 155866 119200 155922 120000 6 x[0]
port 695 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 x[1]
port 696 nsew signal output
rlabel metal3 s 179200 41896 180000 42016 6 x[2]
port 697 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 x[3]
port 698 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 x[4]
port 699 nsew signal output
rlabel metal3 s 179200 69776 180000 69896 6 x[5]
port 700 nsew signal output
rlabel metal3 s 179200 85824 180000 85944 6 x[6]
port 701 nsew signal output
rlabel metal2 s 177670 0 177726 800 6 x[7]
port 702 nsew signal output
rlabel metal3 s 179200 5856 180000 5976 6 y
port 703 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6950022
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/sample.magic.gds
string GDS_START 349090
<< end >>

