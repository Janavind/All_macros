magic
tech sky130A
magscale 1 2
timestamp 1654236653
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118108
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9678 119200 9734 120000
rect 11150 119200 11206 120000
rect 12622 119200 12678 120000
rect 14094 119200 14150 120000
rect 15566 119200 15622 120000
rect 17038 119200 17094 120000
rect 18602 119200 18658 120000
rect 20074 119200 20130 120000
rect 21546 119200 21602 120000
rect 23018 119200 23074 120000
rect 24490 119200 24546 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30470 119200 30526 120000
rect 31942 119200 31998 120000
rect 33414 119200 33470 120000
rect 34886 119200 34942 120000
rect 36450 119200 36506 120000
rect 37922 119200 37978 120000
rect 39394 119200 39450 120000
rect 40866 119200 40922 120000
rect 42338 119200 42394 120000
rect 43902 119200 43958 120000
rect 45374 119200 45430 120000
rect 46846 119200 46902 120000
rect 48318 119200 48374 120000
rect 49790 119200 49846 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54298 119200 54354 120000
rect 55770 119200 55826 120000
rect 57242 119200 57298 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63222 119200 63278 120000
rect 64694 119200 64750 120000
rect 66166 119200 66222 120000
rect 67638 119200 67694 120000
rect 69110 119200 69166 120000
rect 70674 119200 70730 120000
rect 72146 119200 72202 120000
rect 73618 119200 73674 120000
rect 75090 119200 75146 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79598 119200 79654 120000
rect 81070 119200 81126 120000
rect 82542 119200 82598 120000
rect 84014 119200 84070 120000
rect 85486 119200 85542 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89994 119200 90050 120000
rect 91466 119200 91522 120000
rect 92938 119200 92994 120000
rect 94410 119200 94466 120000
rect 95974 119200 96030 120000
rect 97446 119200 97502 120000
rect 98918 119200 98974 120000
rect 100390 119200 100446 120000
rect 101862 119200 101918 120000
rect 103334 119200 103390 120000
rect 104898 119200 104954 120000
rect 106370 119200 106426 120000
rect 107842 119200 107898 120000
rect 109314 119200 109370 120000
rect 110786 119200 110842 120000
rect 112350 119200 112406 120000
rect 113822 119200 113878 120000
rect 115294 119200 115350 120000
rect 116766 119200 116822 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122746 119200 122802 120000
rect 124218 119200 124274 120000
rect 125690 119200 125746 120000
rect 127162 119200 127218 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131670 119200 131726 120000
rect 133142 119200 133198 120000
rect 134614 119200 134670 120000
rect 136086 119200 136142 120000
rect 137558 119200 137614 120000
rect 139122 119200 139178 120000
rect 140594 119200 140650 120000
rect 142066 119200 142122 120000
rect 143538 119200 143594 120000
rect 145010 119200 145066 120000
rect 146574 119200 146630 120000
rect 148046 119200 148102 120000
rect 149518 119200 149574 120000
rect 150990 119200 151046 120000
rect 152462 119200 152518 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 156970 119200 157026 120000
rect 158442 119200 158498 120000
rect 159914 119200 159970 120000
rect 161386 119200 161442 120000
rect 162858 119200 162914 120000
rect 164422 119200 164478 120000
rect 165894 119200 165950 120000
rect 167366 119200 167422 120000
rect 168838 119200 168894 120000
rect 170310 119200 170366 120000
rect 171782 119200 171838 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29642 0 29698 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92386 0 92442 800
rect 92754 0 92810 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95330 0 95386 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125598 0 125654 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126702 0 126758 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129922 0 129978 800
rect 130290 0 130346 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132866 0 132922 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153750 0 153806 800
rect 154118 0 154174 800
rect 154486 0 154542 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155590 0 155646 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157338 0 157394 800
rect 157706 0 157762 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161662 0 161718 800
rect 162030 0 162086 800
rect 162398 0 162454 800
rect 162766 0 162822 800
rect 163134 0 163190 800
rect 163502 0 163558 800
rect 163870 0 163926 800
rect 164238 0 164294 800
rect 164606 0 164662 800
rect 164974 0 165030 800
rect 165342 0 165398 800
rect 165710 0 165766 800
rect 166078 0 166134 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 167090 0 167146 800
rect 167458 0 167514 800
rect 167826 0 167882 800
rect 168194 0 168250 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 170034 0 170090 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6586 119354
rect 6754 119144 8058 119354
rect 8226 119144 9622 119354
rect 9790 119144 11094 119354
rect 11262 119144 12566 119354
rect 12734 119144 14038 119354
rect 14206 119144 15510 119354
rect 15678 119144 16982 119354
rect 17150 119144 18546 119354
rect 18714 119144 20018 119354
rect 20186 119144 21490 119354
rect 21658 119144 22962 119354
rect 23130 119144 24434 119354
rect 24602 119144 25906 119354
rect 26074 119144 27470 119354
rect 27638 119144 28942 119354
rect 29110 119144 30414 119354
rect 30582 119144 31886 119354
rect 32054 119144 33358 119354
rect 33526 119144 34830 119354
rect 34998 119144 36394 119354
rect 36562 119144 37866 119354
rect 38034 119144 39338 119354
rect 39506 119144 40810 119354
rect 40978 119144 42282 119354
rect 42450 119144 43846 119354
rect 44014 119144 45318 119354
rect 45486 119144 46790 119354
rect 46958 119144 48262 119354
rect 48430 119144 49734 119354
rect 49902 119144 51206 119354
rect 51374 119144 52770 119354
rect 52938 119144 54242 119354
rect 54410 119144 55714 119354
rect 55882 119144 57186 119354
rect 57354 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61694 119354
rect 61862 119144 63166 119354
rect 63334 119144 64638 119354
rect 64806 119144 66110 119354
rect 66278 119144 67582 119354
rect 67750 119144 69054 119354
rect 69222 119144 70618 119354
rect 70786 119144 72090 119354
rect 72258 119144 73562 119354
rect 73730 119144 75034 119354
rect 75202 119144 76506 119354
rect 76674 119144 78070 119354
rect 78238 119144 79542 119354
rect 79710 119144 81014 119354
rect 81182 119144 82486 119354
rect 82654 119144 83958 119354
rect 84126 119144 85430 119354
rect 85598 119144 86994 119354
rect 87162 119144 88466 119354
rect 88634 119144 89938 119354
rect 90106 119144 91410 119354
rect 91578 119144 92882 119354
rect 93050 119144 94354 119354
rect 94522 119144 95918 119354
rect 96086 119144 97390 119354
rect 97558 119144 98862 119354
rect 99030 119144 100334 119354
rect 100502 119144 101806 119354
rect 101974 119144 103278 119354
rect 103446 119144 104842 119354
rect 105010 119144 106314 119354
rect 106482 119144 107786 119354
rect 107954 119144 109258 119354
rect 109426 119144 110730 119354
rect 110898 119144 112294 119354
rect 112462 119144 113766 119354
rect 113934 119144 115238 119354
rect 115406 119144 116710 119354
rect 116878 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121218 119354
rect 121386 119144 122690 119354
rect 122858 119144 124162 119354
rect 124330 119144 125634 119354
rect 125802 119144 127106 119354
rect 127274 119144 128578 119354
rect 128746 119144 130142 119354
rect 130310 119144 131614 119354
rect 131782 119144 133086 119354
rect 133254 119144 134558 119354
rect 134726 119144 136030 119354
rect 136198 119144 137502 119354
rect 137670 119144 139066 119354
rect 139234 119144 140538 119354
rect 140706 119144 142010 119354
rect 142178 119144 143482 119354
rect 143650 119144 144954 119354
rect 145122 119144 146518 119354
rect 146686 119144 147990 119354
rect 148158 119144 149462 119354
rect 149630 119144 150934 119354
rect 151102 119144 152406 119354
rect 152574 119144 153878 119354
rect 154046 119144 155442 119354
rect 155610 119144 156914 119354
rect 157082 119144 158386 119354
rect 158554 119144 159858 119354
rect 160026 119144 161330 119354
rect 161498 119144 162802 119354
rect 162970 119144 164366 119354
rect 164534 119144 165838 119354
rect 166006 119144 167310 119354
rect 167478 119144 168782 119354
rect 168950 119144 170254 119354
rect 170422 119144 171726 119354
rect 171894 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177632 119354
rect 756 856 177632 119144
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4378 856
rect 4546 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6862 856
rect 7030 800 7230 856
rect 7398 800 7598 856
rect 7766 800 7966 856
rect 8134 800 8334 856
rect 8502 800 8702 856
rect 8870 800 9070 856
rect 9238 800 9346 856
rect 9514 800 9714 856
rect 9882 800 10082 856
rect 10250 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 13026 856
rect 13194 800 13394 856
rect 13562 800 13762 856
rect 13930 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16614 856
rect 16782 800 16982 856
rect 17150 800 17350 856
rect 17518 800 17718 856
rect 17886 800 18086 856
rect 18254 800 18454 856
rect 18622 800 18730 856
rect 18898 800 19098 856
rect 19266 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23054 856
rect 23222 800 23422 856
rect 23590 800 23790 856
rect 23958 800 24158 856
rect 24326 800 24526 856
rect 24694 800 24894 856
rect 25062 800 25262 856
rect 25430 800 25630 856
rect 25798 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26734 856
rect 26902 800 27102 856
rect 27270 800 27470 856
rect 27638 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29586 856
rect 29754 800 29954 856
rect 30122 800 30322 856
rect 30490 800 30690 856
rect 30858 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33174 856
rect 33342 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34646 856
rect 34814 800 35014 856
rect 35182 800 35382 856
rect 35550 800 35750 856
rect 35918 800 36118 856
rect 36286 800 36486 856
rect 36654 800 36854 856
rect 37022 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38234 856
rect 38402 800 38602 856
rect 38770 800 38970 856
rect 39138 800 39338 856
rect 39506 800 39706 856
rect 39874 800 40074 856
rect 40242 800 40442 856
rect 40610 800 40810 856
rect 40978 800 41178 856
rect 41346 800 41546 856
rect 41714 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42558 856
rect 42726 800 42926 856
rect 43094 800 43294 856
rect 43462 800 43662 856
rect 43830 800 44030 856
rect 44198 800 44398 856
rect 44566 800 44766 856
rect 44934 800 45134 856
rect 45302 800 45502 856
rect 45670 800 45870 856
rect 46038 800 46146 856
rect 46314 800 46514 856
rect 46682 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47618 856
rect 47786 800 47986 856
rect 48154 800 48354 856
rect 48522 800 48722 856
rect 48890 800 49090 856
rect 49258 800 49458 856
rect 49626 800 49826 856
rect 49994 800 50194 856
rect 50362 800 50562 856
rect 50730 800 50838 856
rect 51006 800 51206 856
rect 51374 800 51574 856
rect 51742 800 51942 856
rect 52110 800 52310 856
rect 52478 800 52678 856
rect 52846 800 53046 856
rect 53214 800 53414 856
rect 53582 800 53782 856
rect 53950 800 54150 856
rect 54318 800 54518 856
rect 54686 800 54886 856
rect 55054 800 55254 856
rect 55422 800 55530 856
rect 55698 800 55898 856
rect 56066 800 56266 856
rect 56434 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57370 856
rect 57538 800 57738 856
rect 57906 800 58106 856
rect 58274 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59210 856
rect 59378 800 59578 856
rect 59746 800 59946 856
rect 60114 800 60222 856
rect 60390 800 60590 856
rect 60758 800 60958 856
rect 61126 800 61326 856
rect 61494 800 61694 856
rect 61862 800 62062 856
rect 62230 800 62430 856
rect 62598 800 62798 856
rect 62966 800 63166 856
rect 63334 800 63534 856
rect 63702 800 63902 856
rect 64070 800 64270 856
rect 64438 800 64638 856
rect 64806 800 64914 856
rect 65082 800 65282 856
rect 65450 800 65650 856
rect 65818 800 66018 856
rect 66186 800 66386 856
rect 66554 800 66754 856
rect 66922 800 67122 856
rect 67290 800 67490 856
rect 67658 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68594 856
rect 68762 800 68962 856
rect 69130 800 69238 856
rect 69406 800 69606 856
rect 69774 800 69974 856
rect 70142 800 70342 856
rect 70510 800 70710 856
rect 70878 800 71078 856
rect 71246 800 71446 856
rect 71614 800 71814 856
rect 71982 800 72182 856
rect 72350 800 72550 856
rect 72718 800 72918 856
rect 73086 800 73286 856
rect 73454 800 73654 856
rect 73822 800 73930 856
rect 74098 800 74298 856
rect 74466 800 74666 856
rect 74834 800 75034 856
rect 75202 800 75402 856
rect 75570 800 75770 856
rect 75938 800 76138 856
rect 76306 800 76506 856
rect 76674 800 76874 856
rect 77042 800 77242 856
rect 77410 800 77610 856
rect 77778 800 77978 856
rect 78146 800 78346 856
rect 78514 800 78622 856
rect 78790 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79726 856
rect 79894 800 80094 856
rect 80262 800 80462 856
rect 80630 800 80830 856
rect 80998 800 81198 856
rect 81366 800 81566 856
rect 81734 800 81934 856
rect 82102 800 82302 856
rect 82470 800 82670 856
rect 82838 800 83038 856
rect 83206 800 83314 856
rect 83482 800 83682 856
rect 83850 800 84050 856
rect 84218 800 84418 856
rect 84586 800 84786 856
rect 84954 800 85154 856
rect 85322 800 85522 856
rect 85690 800 85890 856
rect 86058 800 86258 856
rect 86426 800 86626 856
rect 86794 800 86994 856
rect 87162 800 87362 856
rect 87530 800 87730 856
rect 87898 800 88006 856
rect 88174 800 88374 856
rect 88542 800 88742 856
rect 88910 800 89110 856
rect 89278 800 89478 856
rect 89646 800 89846 856
rect 90014 800 90214 856
rect 90382 800 90582 856
rect 90750 800 90950 856
rect 91118 800 91318 856
rect 91486 800 91686 856
rect 91854 800 92054 856
rect 92222 800 92330 856
rect 92498 800 92698 856
rect 92866 800 93066 856
rect 93234 800 93434 856
rect 93602 800 93802 856
rect 93970 800 94170 856
rect 94338 800 94538 856
rect 94706 800 94906 856
rect 95074 800 95274 856
rect 95442 800 95642 856
rect 95810 800 96010 856
rect 96178 800 96378 856
rect 96546 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97390 856
rect 97558 800 97758 856
rect 97926 800 98126 856
rect 98294 800 98494 856
rect 98662 800 98862 856
rect 99030 800 99230 856
rect 99398 800 99598 856
rect 99766 800 99966 856
rect 100134 800 100334 856
rect 100502 800 100702 856
rect 100870 800 101070 856
rect 101238 800 101438 856
rect 101606 800 101714 856
rect 101882 800 102082 856
rect 102250 800 102450 856
rect 102618 800 102818 856
rect 102986 800 103186 856
rect 103354 800 103554 856
rect 103722 800 103922 856
rect 104090 800 104290 856
rect 104458 800 104658 856
rect 104826 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105762 856
rect 105930 800 106130 856
rect 106298 800 106406 856
rect 106574 800 106774 856
rect 106942 800 107142 856
rect 107310 800 107510 856
rect 107678 800 107878 856
rect 108046 800 108246 856
rect 108414 800 108614 856
rect 108782 800 108982 856
rect 109150 800 109350 856
rect 109518 800 109718 856
rect 109886 800 110086 856
rect 110254 800 110454 856
rect 110622 800 110822 856
rect 110990 800 111098 856
rect 111266 800 111466 856
rect 111634 800 111834 856
rect 112002 800 112202 856
rect 112370 800 112570 856
rect 112738 800 112938 856
rect 113106 800 113306 856
rect 113474 800 113674 856
rect 113842 800 114042 856
rect 114210 800 114410 856
rect 114578 800 114778 856
rect 114946 800 115146 856
rect 115314 800 115422 856
rect 115590 800 115790 856
rect 115958 800 116158 856
rect 116326 800 116526 856
rect 116694 800 116894 856
rect 117062 800 117262 856
rect 117430 800 117630 856
rect 117798 800 117998 856
rect 118166 800 118366 856
rect 118534 800 118734 856
rect 118902 800 119102 856
rect 119270 800 119470 856
rect 119638 800 119838 856
rect 120006 800 120114 856
rect 120282 800 120482 856
rect 120650 800 120850 856
rect 121018 800 121218 856
rect 121386 800 121586 856
rect 121754 800 121954 856
rect 122122 800 122322 856
rect 122490 800 122690 856
rect 122858 800 123058 856
rect 123226 800 123426 856
rect 123594 800 123794 856
rect 123962 800 124162 856
rect 124330 800 124530 856
rect 124698 800 124806 856
rect 124974 800 125174 856
rect 125342 800 125542 856
rect 125710 800 125910 856
rect 126078 800 126278 856
rect 126446 800 126646 856
rect 126814 800 127014 856
rect 127182 800 127382 856
rect 127550 800 127750 856
rect 127918 800 128118 856
rect 128286 800 128486 856
rect 128654 800 128854 856
rect 129022 800 129222 856
rect 129390 800 129498 856
rect 129666 800 129866 856
rect 130034 800 130234 856
rect 130402 800 130602 856
rect 130770 800 130970 856
rect 131138 800 131338 856
rect 131506 800 131706 856
rect 131874 800 132074 856
rect 132242 800 132442 856
rect 132610 800 132810 856
rect 132978 800 133178 856
rect 133346 800 133546 856
rect 133714 800 133914 856
rect 134082 800 134190 856
rect 134358 800 134558 856
rect 134726 800 134926 856
rect 135094 800 135294 856
rect 135462 800 135662 856
rect 135830 800 136030 856
rect 136198 800 136398 856
rect 136566 800 136766 856
rect 136934 800 137134 856
rect 137302 800 137502 856
rect 137670 800 137870 856
rect 138038 800 138238 856
rect 138406 800 138514 856
rect 138682 800 138882 856
rect 139050 800 139250 856
rect 139418 800 139618 856
rect 139786 800 139986 856
rect 140154 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141090 856
rect 141258 800 141458 856
rect 141626 800 141826 856
rect 141994 800 142194 856
rect 142362 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143206 856
rect 143374 800 143574 856
rect 143742 800 143942 856
rect 144110 800 144310 856
rect 144478 800 144678 856
rect 144846 800 145046 856
rect 145214 800 145414 856
rect 145582 800 145782 856
rect 145950 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146886 856
rect 147054 800 147254 856
rect 147422 800 147622 856
rect 147790 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 149002 856
rect 149170 800 149370 856
rect 149538 800 149738 856
rect 149906 800 150106 856
rect 150274 800 150474 856
rect 150642 800 150842 856
rect 151010 800 151210 856
rect 151378 800 151578 856
rect 151746 800 151946 856
rect 152114 800 152314 856
rect 152482 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153326 856
rect 153494 800 153694 856
rect 153862 800 154062 856
rect 154230 800 154430 856
rect 154598 800 154798 856
rect 154966 800 155166 856
rect 155334 800 155534 856
rect 155702 800 155902 856
rect 156070 800 156270 856
rect 156438 800 156638 856
rect 156806 800 157006 856
rect 157174 800 157282 856
rect 157450 800 157650 856
rect 157818 800 158018 856
rect 158186 800 158386 856
rect 158554 800 158754 856
rect 158922 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160594 856
rect 160762 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161606 856
rect 161774 800 161974 856
rect 162142 800 162342 856
rect 162510 800 162710 856
rect 162878 800 163078 856
rect 163246 800 163446 856
rect 163614 800 163814 856
rect 163982 800 164182 856
rect 164350 800 164550 856
rect 164718 800 164918 856
rect 165086 800 165286 856
rect 165454 800 165654 856
rect 165822 800 166022 856
rect 166190 800 166298 856
rect 166466 800 166666 856
rect 166834 800 167034 856
rect 167202 800 167402 856
rect 167570 800 167770 856
rect 167938 800 168138 856
rect 168306 800 168506 856
rect 168674 800 168874 856
rect 169042 800 169242 856
rect 169410 800 169610 856
rect 169778 800 169978 856
rect 170146 800 170346 856
rect 170514 800 170714 856
rect 170882 800 170990 856
rect 171158 800 171358 856
rect 171526 800 171726 856
rect 171894 800 172094 856
rect 172262 800 172462 856
rect 172630 800 172830 856
rect 172998 800 173198 856
rect 173366 800 173566 856
rect 173734 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
rect 175574 800 175682 856
rect 175850 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
<< metal3 >>
rect 0 113840 800 113960
rect 179200 112344 180000 112464
rect 0 101872 800 101992
rect 179200 97384 180000 97504
rect 0 89904 800 90024
rect 179200 82424 180000 82544
rect 0 77936 800 78056
rect 179200 67464 180000 67584
rect 0 65968 800 66088
rect 0 53864 800 53984
rect 179200 52368 180000 52488
rect 0 41896 800 42016
rect 179200 37408 180000 37528
rect 0 29928 800 30048
rect 179200 22448 180000 22568
rect 0 17960 800 18080
rect 179200 7488 180000 7608
rect 0 5992 800 6112
<< obsm3 >>
rect 800 114040 173488 117605
rect 880 113760 173488 114040
rect 800 102072 173488 113760
rect 880 101792 173488 102072
rect 800 90104 173488 101792
rect 880 89824 173488 90104
rect 800 78136 173488 89824
rect 880 77856 173488 78136
rect 800 66168 173488 77856
rect 880 65888 173488 66168
rect 800 54064 173488 65888
rect 880 53784 173488 54064
rect 800 42096 173488 53784
rect 880 41816 173488 42096
rect 800 30128 173488 41816
rect 880 29848 173488 30128
rect 800 18160 173488 29848
rect 880 17880 173488 18160
rect 800 6192 173488 17880
rect 880 5912 173488 6192
rect 800 2143 173488 5912
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 84147 3299 94333 117469
<< labels >>
rlabel metal3 s 0 5992 800 6112 6 active
port 1 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 0 65968 800 66088 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal3 s 179200 67464 180000 67584 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 179200 82424 180000 82544 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 179200 97384 180000 97504 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal3 s 0 77936 800 78056 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 179200 112344 180000 112464 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal3 s 0 89904 800 90024 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal2 s 176842 0 176898 800 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal3 s 0 101872 800 101992 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 0 113840 800 113960 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 0 41896 800 42016 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 0 53864 800 53984 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 179200 7488 180000 7608 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 179200 22448 180000 22568 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 179200 37408 180000 37528 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 179200 52368 180000 52488 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 45374 119200 45430 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 49790 119200 49846 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 54298 119200 54354 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 58714 119200 58770 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 63222 119200 63278 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 67638 119200 67694 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 81070 119200 81126 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 85486 119200 85542 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 89994 119200 90050 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 94410 119200 94466 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 98918 119200 98974 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 103334 119200 103390 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 107842 119200 107898 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 116766 119200 116822 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 121274 119200 121330 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 125690 119200 125746 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 130198 119200 130254 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 148046 119200 148102 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 152462 119200 152518 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 156970 119200 157026 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 161386 119200 161442 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 165894 119200 165950 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 14094 119200 14150 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18602 119200 18658 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 23018 119200 23074 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 27526 119200 27582 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31942 119200 31998 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 36450 119200 36506 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 40866 119200 40922 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 46846 119200 46902 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 69110 119200 69166 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 73618 119200 73674 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 95974 119200 96030 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 100390 119200 100446 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 104898 119200 104954 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 109314 119200 109370 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 113822 119200 113878 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 122746 119200 122802 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 127162 119200 127218 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 131670 119200 131726 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 11150 119200 11206 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 140594 119200 140650 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 145010 119200 145066 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 149518 119200 149574 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 158442 119200 158498 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 162858 119200 162914 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15566 119200 15622 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 33414 119200 33470 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 37922 119200 37978 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 42338 119200 42394 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 48318 119200 48374 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 57242 119200 57298 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 61750 119200 61806 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 66166 119200 66222 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 84014 119200 84070 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 92938 119200 92994 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 101862 119200 101918 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 128634 119200 128690 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 133142 119200 133198 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12622 119200 12678 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 137558 119200 137614 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 142066 119200 142122 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 146574 119200 146630 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 150990 119200 151046 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 159914 119200 159970 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 164422 119200 164478 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 168838 119200 168894 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 17038 119200 17094 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21546 119200 21602 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 43902 119200 43958 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 151266 0 151322 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 171782 0 171838 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 175094 0 175150 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 164606 0 164662 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal2 s 170310 119200 170366 120000 6 user_clock2
port 529 nsew signal input
rlabel metal2 s 171782 119200 171838 120000 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 user_irq[1]
port 531 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6486174
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_13.magic.gds
string GDS_START 307724
<< end >>

