magic
tech sky130A
magscale 1 2
timestamp 1654284974
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 117904
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6734 119200 6790 120000
rect 8206 119200 8262 120000
rect 9678 119200 9734 120000
rect 11242 119200 11298 120000
rect 12714 119200 12770 120000
rect 14186 119200 14242 120000
rect 15750 119200 15806 120000
rect 17222 119200 17278 120000
rect 18694 119200 18750 120000
rect 20258 119200 20314 120000
rect 21730 119200 21786 120000
rect 23202 119200 23258 120000
rect 24674 119200 24730 120000
rect 26238 119200 26294 120000
rect 27710 119200 27766 120000
rect 29182 119200 29238 120000
rect 30746 119200 30802 120000
rect 32218 119200 32274 120000
rect 33690 119200 33746 120000
rect 35254 119200 35310 120000
rect 36726 119200 36782 120000
rect 38198 119200 38254 120000
rect 39762 119200 39818 120000
rect 41234 119200 41290 120000
rect 42706 119200 42762 120000
rect 44178 119200 44234 120000
rect 45742 119200 45798 120000
rect 47214 119200 47270 120000
rect 48686 119200 48742 120000
rect 50250 119200 50306 120000
rect 51722 119200 51778 120000
rect 53194 119200 53250 120000
rect 54758 119200 54814 120000
rect 56230 119200 56286 120000
rect 57702 119200 57758 120000
rect 59266 119200 59322 120000
rect 60738 119200 60794 120000
rect 62210 119200 62266 120000
rect 63682 119200 63738 120000
rect 65246 119200 65302 120000
rect 66718 119200 66774 120000
rect 68190 119200 68246 120000
rect 69754 119200 69810 120000
rect 71226 119200 71282 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75734 119200 75790 120000
rect 77206 119200 77262 120000
rect 78770 119200 78826 120000
rect 80242 119200 80298 120000
rect 81714 119200 81770 120000
rect 83186 119200 83242 120000
rect 84750 119200 84806 120000
rect 86222 119200 86278 120000
rect 87694 119200 87750 120000
rect 89258 119200 89314 120000
rect 90730 119200 90786 120000
rect 92202 119200 92258 120000
rect 93766 119200 93822 120000
rect 95238 119200 95294 120000
rect 96710 119200 96766 120000
rect 98274 119200 98330 120000
rect 99746 119200 99802 120000
rect 101218 119200 101274 120000
rect 102690 119200 102746 120000
rect 104254 119200 104310 120000
rect 105726 119200 105782 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110234 119200 110290 120000
rect 111706 119200 111762 120000
rect 113270 119200 113326 120000
rect 114742 119200 114798 120000
rect 116214 119200 116270 120000
rect 117778 119200 117834 120000
rect 119250 119200 119306 120000
rect 120722 119200 120778 120000
rect 122194 119200 122250 120000
rect 123758 119200 123814 120000
rect 125230 119200 125286 120000
rect 126702 119200 126758 120000
rect 128266 119200 128322 120000
rect 129738 119200 129794 120000
rect 131210 119200 131266 120000
rect 132774 119200 132830 120000
rect 134246 119200 134302 120000
rect 135718 119200 135774 120000
rect 137282 119200 137338 120000
rect 138754 119200 138810 120000
rect 140226 119200 140282 120000
rect 141698 119200 141754 120000
rect 143262 119200 143318 120000
rect 144734 119200 144790 120000
rect 146206 119200 146262 120000
rect 147770 119200 147826 120000
rect 149242 119200 149298 120000
rect 150714 119200 150770 120000
rect 152278 119200 152334 120000
rect 153750 119200 153806 120000
rect 155222 119200 155278 120000
rect 156786 119200 156842 120000
rect 158258 119200 158314 120000
rect 159730 119200 159786 120000
rect 161202 119200 161258 120000
rect 162766 119200 162822 120000
rect 164238 119200 164294 120000
rect 165710 119200 165766 120000
rect 167274 119200 167330 120000
rect 168746 119200 168802 120000
rect 170218 119200 170274 120000
rect 171782 119200 171838 120000
rect 173254 119200 173310 120000
rect 174726 119200 174782 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42982 0 43038 800
rect 43350 0 43406 800
rect 43718 0 43774 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46662 0 46718 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49514 0 49570 800
rect 49882 0 49938 800
rect 50250 0 50306 800
rect 50618 0 50674 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 52090 0 52146 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53194 0 53250 800
rect 53562 0 53618 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65154 0 65210 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70582 0 70638 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76102 0 76158 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83002 0 83058 800
rect 83370 0 83426 800
rect 83738 0 83794 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95330 0 95386 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100482 0 100538 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109222 0 109278 800
rect 109590 0 109646 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113914 0 113970 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118238 0 118294 800
rect 118606 0 118662 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124494 0 124550 800
rect 124862 0 124918 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 128082 0 128138 800
rect 128450 0 128506 800
rect 128818 0 128874 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129922 0 129978 800
rect 130290 0 130346 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131394 0 131450 800
rect 131762 0 131818 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132866 0 132922 800
rect 133142 0 133198 800
rect 133510 0 133566 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152462 0 152518 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155406 0 155462 800
rect 155774 0 155830 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157522 0 157578 800
rect 157890 0 157946 800
rect 158258 0 158314 800
rect 158626 0 158682 800
rect 158994 0 159050 800
rect 159362 0 159418 800
rect 159730 0 159786 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161938 0 161994 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163778 0 163834 800
rect 164146 0 164202 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166262 0 166318 800
rect 166630 0 166686 800
rect 166998 0 167054 800
rect 167366 0 167422 800
rect 167734 0 167790 800
rect 168102 0 168158 800
rect 168470 0 168526 800
rect 168838 0 168894 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6678 119354
rect 6846 119144 8150 119354
rect 8318 119144 9622 119354
rect 9790 119144 11186 119354
rect 11354 119144 12658 119354
rect 12826 119144 14130 119354
rect 14298 119144 15694 119354
rect 15862 119144 17166 119354
rect 17334 119144 18638 119354
rect 18806 119144 20202 119354
rect 20370 119144 21674 119354
rect 21842 119144 23146 119354
rect 23314 119144 24618 119354
rect 24786 119144 26182 119354
rect 26350 119144 27654 119354
rect 27822 119144 29126 119354
rect 29294 119144 30690 119354
rect 30858 119144 32162 119354
rect 32330 119144 33634 119354
rect 33802 119144 35198 119354
rect 35366 119144 36670 119354
rect 36838 119144 38142 119354
rect 38310 119144 39706 119354
rect 39874 119144 41178 119354
rect 41346 119144 42650 119354
rect 42818 119144 44122 119354
rect 44290 119144 45686 119354
rect 45854 119144 47158 119354
rect 47326 119144 48630 119354
rect 48798 119144 50194 119354
rect 50362 119144 51666 119354
rect 51834 119144 53138 119354
rect 53306 119144 54702 119354
rect 54870 119144 56174 119354
rect 56342 119144 57646 119354
rect 57814 119144 59210 119354
rect 59378 119144 60682 119354
rect 60850 119144 62154 119354
rect 62322 119144 63626 119354
rect 63794 119144 65190 119354
rect 65358 119144 66662 119354
rect 66830 119144 68134 119354
rect 68302 119144 69698 119354
rect 69866 119144 71170 119354
rect 71338 119144 72642 119354
rect 72810 119144 74206 119354
rect 74374 119144 75678 119354
rect 75846 119144 77150 119354
rect 77318 119144 78714 119354
rect 78882 119144 80186 119354
rect 80354 119144 81658 119354
rect 81826 119144 83130 119354
rect 83298 119144 84694 119354
rect 84862 119144 86166 119354
rect 86334 119144 87638 119354
rect 87806 119144 89202 119354
rect 89370 119144 90674 119354
rect 90842 119144 92146 119354
rect 92314 119144 93710 119354
rect 93878 119144 95182 119354
rect 95350 119144 96654 119354
rect 96822 119144 98218 119354
rect 98386 119144 99690 119354
rect 99858 119144 101162 119354
rect 101330 119144 102634 119354
rect 102802 119144 104198 119354
rect 104366 119144 105670 119354
rect 105838 119144 107142 119354
rect 107310 119144 108706 119354
rect 108874 119144 110178 119354
rect 110346 119144 111650 119354
rect 111818 119144 113214 119354
rect 113382 119144 114686 119354
rect 114854 119144 116158 119354
rect 116326 119144 117722 119354
rect 117890 119144 119194 119354
rect 119362 119144 120666 119354
rect 120834 119144 122138 119354
rect 122306 119144 123702 119354
rect 123870 119144 125174 119354
rect 125342 119144 126646 119354
rect 126814 119144 128210 119354
rect 128378 119144 129682 119354
rect 129850 119144 131154 119354
rect 131322 119144 132718 119354
rect 132886 119144 134190 119354
rect 134358 119144 135662 119354
rect 135830 119144 137226 119354
rect 137394 119144 138698 119354
rect 138866 119144 140170 119354
rect 140338 119144 141642 119354
rect 141810 119144 143206 119354
rect 143374 119144 144678 119354
rect 144846 119144 146150 119354
rect 146318 119144 147714 119354
rect 147882 119144 149186 119354
rect 149354 119144 150658 119354
rect 150826 119144 152222 119354
rect 152390 119144 153694 119354
rect 153862 119144 155166 119354
rect 155334 119144 156730 119354
rect 156898 119144 158202 119354
rect 158370 119144 159674 119354
rect 159842 119144 161146 119354
rect 161314 119144 162710 119354
rect 162878 119144 164182 119354
rect 164350 119144 165654 119354
rect 165822 119144 167218 119354
rect 167386 119144 168690 119354
rect 168858 119144 170162 119354
rect 170330 119144 171726 119354
rect 171894 119144 173198 119354
rect 173366 119144 174670 119354
rect 174838 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7322 856
rect 7490 734 7690 856
rect 7858 734 7966 856
rect 8134 734 8334 856
rect 8502 734 8702 856
rect 8870 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9806 856
rect 9974 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12750 856
rect 12918 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14222 856
rect 14390 734 14590 856
rect 14758 734 14958 856
rect 15126 734 15326 856
rect 15494 734 15694 856
rect 15862 734 15970 856
rect 16138 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17810 856
rect 17978 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18914 856
rect 19082 734 19282 856
rect 19450 734 19650 856
rect 19818 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20754 856
rect 20922 734 21122 856
rect 21290 734 21490 856
rect 21658 734 21858 856
rect 22026 734 22226 856
rect 22394 734 22594 856
rect 22762 734 22962 856
rect 23130 734 23330 856
rect 23498 734 23606 856
rect 23774 734 23974 856
rect 24142 734 24342 856
rect 24510 734 24710 856
rect 24878 734 25078 856
rect 25246 734 25446 856
rect 25614 734 25814 856
rect 25982 734 26182 856
rect 26350 734 26550 856
rect 26718 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27654 856
rect 27822 734 28022 856
rect 28190 734 28390 856
rect 28558 734 28758 856
rect 28926 734 29126 856
rect 29294 734 29494 856
rect 29662 734 29862 856
rect 30030 734 30230 856
rect 30398 734 30598 856
rect 30766 734 30966 856
rect 31134 734 31334 856
rect 31502 734 31610 856
rect 31778 734 31978 856
rect 32146 734 32346 856
rect 32514 734 32714 856
rect 32882 734 33082 856
rect 33250 734 33450 856
rect 33618 734 33818 856
rect 33986 734 34186 856
rect 34354 734 34554 856
rect 34722 734 34922 856
rect 35090 734 35290 856
rect 35458 734 35658 856
rect 35826 734 36026 856
rect 36194 734 36394 856
rect 36562 734 36762 856
rect 36930 734 37130 856
rect 37298 734 37498 856
rect 37666 734 37866 856
rect 38034 734 38234 856
rect 38402 734 38602 856
rect 38770 734 38970 856
rect 39138 734 39246 856
rect 39414 734 39614 856
rect 39782 734 39982 856
rect 40150 734 40350 856
rect 40518 734 40718 856
rect 40886 734 41086 856
rect 41254 734 41454 856
rect 41622 734 41822 856
rect 41990 734 42190 856
rect 42358 734 42558 856
rect 42726 734 42926 856
rect 43094 734 43294 856
rect 43462 734 43662 856
rect 43830 734 44030 856
rect 44198 734 44398 856
rect 44566 734 44766 856
rect 44934 734 45134 856
rect 45302 734 45502 856
rect 45670 734 45870 856
rect 46038 734 46238 856
rect 46406 734 46606 856
rect 46774 734 46974 856
rect 47142 734 47250 856
rect 47418 734 47618 856
rect 47786 734 47986 856
rect 48154 734 48354 856
rect 48522 734 48722 856
rect 48890 734 49090 856
rect 49258 734 49458 856
rect 49626 734 49826 856
rect 49994 734 50194 856
rect 50362 734 50562 856
rect 50730 734 50930 856
rect 51098 734 51298 856
rect 51466 734 51666 856
rect 51834 734 52034 856
rect 52202 734 52402 856
rect 52570 734 52770 856
rect 52938 734 53138 856
rect 53306 734 53506 856
rect 53674 734 53874 856
rect 54042 734 54242 856
rect 54410 734 54610 856
rect 54778 734 54886 856
rect 55054 734 55254 856
rect 55422 734 55622 856
rect 55790 734 55990 856
rect 56158 734 56358 856
rect 56526 734 56726 856
rect 56894 734 57094 856
rect 57262 734 57462 856
rect 57630 734 57830 856
rect 57998 734 58198 856
rect 58366 734 58566 856
rect 58734 734 58934 856
rect 59102 734 59302 856
rect 59470 734 59670 856
rect 59838 734 60038 856
rect 60206 734 60406 856
rect 60574 734 60774 856
rect 60942 734 61142 856
rect 61310 734 61510 856
rect 61678 734 61878 856
rect 62046 734 62246 856
rect 62414 734 62614 856
rect 62782 734 62890 856
rect 63058 734 63258 856
rect 63426 734 63626 856
rect 63794 734 63994 856
rect 64162 734 64362 856
rect 64530 734 64730 856
rect 64898 734 65098 856
rect 65266 734 65466 856
rect 65634 734 65834 856
rect 66002 734 66202 856
rect 66370 734 66570 856
rect 66738 734 66938 856
rect 67106 734 67306 856
rect 67474 734 67674 856
rect 67842 734 68042 856
rect 68210 734 68410 856
rect 68578 734 68778 856
rect 68946 734 69146 856
rect 69314 734 69514 856
rect 69682 734 69882 856
rect 70050 734 70250 856
rect 70418 734 70526 856
rect 70694 734 70894 856
rect 71062 734 71262 856
rect 71430 734 71630 856
rect 71798 734 71998 856
rect 72166 734 72366 856
rect 72534 734 72734 856
rect 72902 734 73102 856
rect 73270 734 73470 856
rect 73638 734 73838 856
rect 74006 734 74206 856
rect 74374 734 74574 856
rect 74742 734 74942 856
rect 75110 734 75310 856
rect 75478 734 75678 856
rect 75846 734 76046 856
rect 76214 734 76414 856
rect 76582 734 76782 856
rect 76950 734 77150 856
rect 77318 734 77518 856
rect 77686 734 77886 856
rect 78054 734 78254 856
rect 78422 734 78530 856
rect 78698 734 78898 856
rect 79066 734 79266 856
rect 79434 734 79634 856
rect 79802 734 80002 856
rect 80170 734 80370 856
rect 80538 734 80738 856
rect 80906 734 81106 856
rect 81274 734 81474 856
rect 81642 734 81842 856
rect 82010 734 82210 856
rect 82378 734 82578 856
rect 82746 734 82946 856
rect 83114 734 83314 856
rect 83482 734 83682 856
rect 83850 734 84050 856
rect 84218 734 84418 856
rect 84586 734 84786 856
rect 84954 734 85154 856
rect 85322 734 85522 856
rect 85690 734 85890 856
rect 86058 734 86166 856
rect 86334 734 86534 856
rect 86702 734 86902 856
rect 87070 734 87270 856
rect 87438 734 87638 856
rect 87806 734 88006 856
rect 88174 734 88374 856
rect 88542 734 88742 856
rect 88910 734 89110 856
rect 89278 734 89478 856
rect 89646 734 89846 856
rect 90014 734 90214 856
rect 90382 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91318 856
rect 91486 734 91686 856
rect 91854 734 92054 856
rect 92222 734 92422 856
rect 92590 734 92790 856
rect 92958 734 93158 856
rect 93326 734 93526 856
rect 93694 734 93894 856
rect 94062 734 94170 856
rect 94338 734 94538 856
rect 94706 734 94906 856
rect 95074 734 95274 856
rect 95442 734 95642 856
rect 95810 734 96010 856
rect 96178 734 96378 856
rect 96546 734 96746 856
rect 96914 734 97114 856
rect 97282 734 97482 856
rect 97650 734 97850 856
rect 98018 734 98218 856
rect 98386 734 98586 856
rect 98754 734 98954 856
rect 99122 734 99322 856
rect 99490 734 99690 856
rect 99858 734 100058 856
rect 100226 734 100426 856
rect 100594 734 100794 856
rect 100962 734 101162 856
rect 101330 734 101530 856
rect 101698 734 101806 856
rect 101974 734 102174 856
rect 102342 734 102542 856
rect 102710 734 102910 856
rect 103078 734 103278 856
rect 103446 734 103646 856
rect 103814 734 104014 856
rect 104182 734 104382 856
rect 104550 734 104750 856
rect 104918 734 105118 856
rect 105286 734 105486 856
rect 105654 734 105854 856
rect 106022 734 106222 856
rect 106390 734 106590 856
rect 106758 734 106958 856
rect 107126 734 107326 856
rect 107494 734 107694 856
rect 107862 734 108062 856
rect 108230 734 108430 856
rect 108598 734 108798 856
rect 108966 734 109166 856
rect 109334 734 109534 856
rect 109702 734 109810 856
rect 109978 734 110178 856
rect 110346 734 110546 856
rect 110714 734 110914 856
rect 111082 734 111282 856
rect 111450 734 111650 856
rect 111818 734 112018 856
rect 112186 734 112386 856
rect 112554 734 112754 856
rect 112922 734 113122 856
rect 113290 734 113490 856
rect 113658 734 113858 856
rect 114026 734 114226 856
rect 114394 734 114594 856
rect 114762 734 114962 856
rect 115130 734 115330 856
rect 115498 734 115698 856
rect 115866 734 116066 856
rect 116234 734 116434 856
rect 116602 734 116802 856
rect 116970 734 117170 856
rect 117338 734 117446 856
rect 117614 734 117814 856
rect 117982 734 118182 856
rect 118350 734 118550 856
rect 118718 734 118918 856
rect 119086 734 119286 856
rect 119454 734 119654 856
rect 119822 734 120022 856
rect 120190 734 120390 856
rect 120558 734 120758 856
rect 120926 734 121126 856
rect 121294 734 121494 856
rect 121662 734 121862 856
rect 122030 734 122230 856
rect 122398 734 122598 856
rect 122766 734 122966 856
rect 123134 734 123334 856
rect 123502 734 123702 856
rect 123870 734 124070 856
rect 124238 734 124438 856
rect 124606 734 124806 856
rect 124974 734 125174 856
rect 125342 734 125450 856
rect 125618 734 125818 856
rect 125986 734 126186 856
rect 126354 734 126554 856
rect 126722 734 126922 856
rect 127090 734 127290 856
rect 127458 734 127658 856
rect 127826 734 128026 856
rect 128194 734 128394 856
rect 128562 734 128762 856
rect 128930 734 129130 856
rect 129298 734 129498 856
rect 129666 734 129866 856
rect 130034 734 130234 856
rect 130402 734 130602 856
rect 130770 734 130970 856
rect 131138 734 131338 856
rect 131506 734 131706 856
rect 131874 734 132074 856
rect 132242 734 132442 856
rect 132610 734 132810 856
rect 132978 734 133086 856
rect 133254 734 133454 856
rect 133622 734 133822 856
rect 133990 734 134190 856
rect 134358 734 134558 856
rect 134726 734 134926 856
rect 135094 734 135294 856
rect 135462 734 135662 856
rect 135830 734 136030 856
rect 136198 734 136398 856
rect 136566 734 136766 856
rect 136934 734 137134 856
rect 137302 734 137502 856
rect 137670 734 137870 856
rect 138038 734 138238 856
rect 138406 734 138606 856
rect 138774 734 138974 856
rect 139142 734 139342 856
rect 139510 734 139710 856
rect 139878 734 140078 856
rect 140246 734 140446 856
rect 140614 734 140814 856
rect 140982 734 141090 856
rect 141258 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142194 856
rect 142362 734 142562 856
rect 142730 734 142930 856
rect 143098 734 143298 856
rect 143466 734 143666 856
rect 143834 734 144034 856
rect 144202 734 144402 856
rect 144570 734 144770 856
rect 144938 734 145138 856
rect 145306 734 145506 856
rect 145674 734 145874 856
rect 146042 734 146242 856
rect 146410 734 146610 856
rect 146778 734 146978 856
rect 147146 734 147346 856
rect 147514 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148450 856
rect 148618 734 148726 856
rect 148894 734 149094 856
rect 149262 734 149462 856
rect 149630 734 149830 856
rect 149998 734 150198 856
rect 150366 734 150566 856
rect 150734 734 150934 856
rect 151102 734 151302 856
rect 151470 734 151670 856
rect 151838 734 152038 856
rect 152206 734 152406 856
rect 152574 734 152774 856
rect 152942 734 153142 856
rect 153310 734 153510 856
rect 153678 734 153878 856
rect 154046 734 154246 856
rect 154414 734 154614 856
rect 154782 734 154982 856
rect 155150 734 155350 856
rect 155518 734 155718 856
rect 155886 734 156086 856
rect 156254 734 156454 856
rect 156622 734 156730 856
rect 156898 734 157098 856
rect 157266 734 157466 856
rect 157634 734 157834 856
rect 158002 734 158202 856
rect 158370 734 158570 856
rect 158738 734 158938 856
rect 159106 734 159306 856
rect 159474 734 159674 856
rect 159842 734 160042 856
rect 160210 734 160410 856
rect 160578 734 160778 856
rect 160946 734 161146 856
rect 161314 734 161514 856
rect 161682 734 161882 856
rect 162050 734 162250 856
rect 162418 734 162618 856
rect 162786 734 162986 856
rect 163154 734 163354 856
rect 163522 734 163722 856
rect 163890 734 164090 856
rect 164258 734 164366 856
rect 164534 734 164734 856
rect 164902 734 165102 856
rect 165270 734 165470 856
rect 165638 734 165838 856
rect 166006 734 166206 856
rect 166374 734 166574 856
rect 166742 734 166942 856
rect 167110 734 167310 856
rect 167478 734 167678 856
rect 167846 734 168046 856
rect 168214 734 168414 856
rect 168582 734 168782 856
rect 168950 734 169150 856
rect 169318 734 169518 856
rect 169686 734 169886 856
rect 170054 734 170254 856
rect 170422 734 170622 856
rect 170790 734 170990 856
rect 171158 734 171358 856
rect 171526 734 171726 856
rect 171894 734 172094 856
rect 172262 734 172370 856
rect 172538 734 172738 856
rect 172906 734 173106 856
rect 173274 734 173474 856
rect 173642 734 173842 856
rect 174010 734 174210 856
rect 174378 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175314 856
rect 175482 734 175682 856
rect 175850 734 176050 856
rect 176218 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178186 856
<< metal3 >>
rect 179200 115608 180000 115728
rect 0 113296 800 113416
rect 179200 107040 180000 107160
rect 0 99968 800 100088
rect 179200 98472 180000 98592
rect 179200 89904 180000 90024
rect 0 86640 800 86760
rect 179200 81336 180000 81456
rect 0 73312 800 73432
rect 179200 72768 180000 72888
rect 179200 64200 180000 64320
rect 0 59984 800 60104
rect 179200 55632 180000 55752
rect 179200 47064 180000 47184
rect 0 46656 800 46776
rect 179200 38496 180000 38616
rect 0 33328 800 33448
rect 179200 29928 180000 30048
rect 179200 21360 180000 21480
rect 0 20000 800 20120
rect 179200 12792 180000 12912
rect 0 6672 800 6792
rect 179200 4224 180000 4344
<< obsm3 >>
rect 800 115808 179200 117741
rect 800 115528 179120 115808
rect 800 113496 179200 115528
rect 880 113216 179200 113496
rect 800 107240 179200 113216
rect 800 106960 179120 107240
rect 800 100168 179200 106960
rect 880 99888 179200 100168
rect 800 98672 179200 99888
rect 800 98392 179120 98672
rect 800 90104 179200 98392
rect 800 89824 179120 90104
rect 800 86840 179200 89824
rect 880 86560 179200 86840
rect 800 81536 179200 86560
rect 800 81256 179120 81536
rect 800 73512 179200 81256
rect 880 73232 179200 73512
rect 800 72968 179200 73232
rect 800 72688 179120 72968
rect 800 64400 179200 72688
rect 800 64120 179120 64400
rect 800 60184 179200 64120
rect 880 59904 179200 60184
rect 800 55832 179200 59904
rect 800 55552 179120 55832
rect 800 47264 179200 55552
rect 800 46984 179120 47264
rect 800 46856 179200 46984
rect 880 46576 179200 46856
rect 800 38696 179200 46576
rect 800 38416 179120 38696
rect 800 33528 179200 38416
rect 880 33248 179200 33528
rect 800 30128 179200 33248
rect 800 29848 179120 30128
rect 800 21560 179200 29848
rect 800 21280 179120 21560
rect 800 20200 179200 21280
rect 880 19920 179200 20200
rect 800 12992 179200 19920
rect 800 12712 179120 12992
rect 800 6872 179200 12712
rect 880 6592 179200 6872
rect 800 4424 179200 6592
rect 800 4144 179120 4424
rect 800 2143 179200 4144
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 88011 5067 96173 117741
<< labels >>
rlabel metal3 s 0 6672 800 6792 6 active
port 1 nsew signal input
rlabel metal2 s 173254 119200 173310 120000 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 179200 47064 180000 47184 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal3 s 179200 55632 180000 55752 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 0 73312 800 73432 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal3 s 179200 64200 180000 64320 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 0 86640 800 86760 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 179200 12792 180000 12912 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal3 s 179200 72768 180000 72888 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal3 s 179200 81336 180000 81456 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal3 s 179200 89904 180000 90024 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 179200 98472 180000 98592 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal3 s 0 99968 800 100088 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal3 s 0 113296 800 113416 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal3 s 179200 107040 180000 107160 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 179200 115608 180000 115728 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 179200 21360 180000 21480 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 0 33328 800 33448 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 179200 29928 180000 30048 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 0 46656 800 46776 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 179200 38496 180000 38616 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 45742 119200 45798 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 50250 119200 50306 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 54758 119200 54814 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 59266 119200 59322 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 63682 119200 63738 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 68190 119200 68246 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 72698 119200 72754 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 77206 119200 77262 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 81714 119200 81770 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 86222 119200 86278 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 95238 119200 95294 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 99746 119200 99802 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 104254 119200 104310 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 113270 119200 113326 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 117778 119200 117834 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 122194 119200 122250 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 126702 119200 126758 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 131210 119200 131266 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 135718 119200 135774 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 140226 119200 140282 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 144734 119200 144790 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 149242 119200 149298 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 153750 119200 153806 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 158258 119200 158314 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 162766 119200 162822 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 167274 119200 167330 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 14186 119200 14242 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18694 119200 18750 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 23202 119200 23258 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 27710 119200 27766 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 32218 119200 32274 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 36726 119200 36782 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 41234 119200 41290 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 47214 119200 47270 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 51722 119200 51778 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 56230 119200 56286 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 65246 119200 65302 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 69754 119200 69810 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 78770 119200 78826 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 83186 119200 83242 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 87694 119200 87750 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6734 119200 6790 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 92202 119200 92258 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 96710 119200 96766 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 101218 119200 101274 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 105726 119200 105782 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 110234 119200 110290 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 114742 119200 114798 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 119250 119200 119306 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 123758 119200 123814 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 128266 119200 128322 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 11242 119200 11298 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 137282 119200 137338 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 141698 119200 141754 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 146206 119200 146262 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 150714 119200 150770 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 155222 119200 155278 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 159730 119200 159786 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 168746 119200 168802 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15750 119200 15806 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 20258 119200 20314 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24674 119200 24730 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 29182 119200 29238 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 33690 119200 33746 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 38198 119200 38254 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 42706 119200 42762 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 48686 119200 48742 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 53194 119200 53250 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 57702 119200 57758 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 62210 119200 62266 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 66718 119200 66774 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 71226 119200 71282 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 80242 119200 80298 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 84750 119200 84806 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 89258 119200 89314 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 8206 119200 8262 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 93766 119200 93822 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 98274 119200 98330 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 102690 119200 102746 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 111706 119200 111762 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 116214 119200 116270 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 120722 119200 120778 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 125230 119200 125286 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 129738 119200 129794 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 134246 119200 134302 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12714 119200 12770 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 138754 119200 138810 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 143262 119200 143318 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 147770 119200 147826 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 152278 119200 152334 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 156786 119200 156842 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 161202 119200 161258 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 165710 119200 165766 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 170218 119200 170274 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21730 119200 21786 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 26238 119200 26294 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 35254 119200 35310 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 39762 119200 39818 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 44178 119200 44234 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 158994 0 159050 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 166630 0 166686 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 168838 0 168894 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 172150 0 172206 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 174266 0 174322 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 126242 0 126298 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal2 s 171782 119200 171838 120000 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 179200 4224 180000 4344 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 174726 119200 174782 120000 6 user_irq[1]
port 531 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7555378
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_decap_3.magic.gds
string GDS_START 297990
<< end >>

