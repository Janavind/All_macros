magic
tech sky130A
magscale 1 2
timestamp 1653957317
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118176
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9678 119200 9734 120000
rect 11150 119200 11206 120000
rect 12622 119200 12678 120000
rect 14094 119200 14150 120000
rect 15566 119200 15622 120000
rect 17038 119200 17094 120000
rect 18602 119200 18658 120000
rect 20074 119200 20130 120000
rect 21546 119200 21602 120000
rect 23018 119200 23074 120000
rect 24490 119200 24546 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30470 119200 30526 120000
rect 31942 119200 31998 120000
rect 33414 119200 33470 120000
rect 34886 119200 34942 120000
rect 36450 119200 36506 120000
rect 37922 119200 37978 120000
rect 39394 119200 39450 120000
rect 40866 119200 40922 120000
rect 42338 119200 42394 120000
rect 43902 119200 43958 120000
rect 45374 119200 45430 120000
rect 46846 119200 46902 120000
rect 48318 119200 48374 120000
rect 49790 119200 49846 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54298 119200 54354 120000
rect 55770 119200 55826 120000
rect 57242 119200 57298 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63222 119200 63278 120000
rect 64694 119200 64750 120000
rect 66166 119200 66222 120000
rect 67638 119200 67694 120000
rect 69110 119200 69166 120000
rect 70674 119200 70730 120000
rect 72146 119200 72202 120000
rect 73618 119200 73674 120000
rect 75090 119200 75146 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79598 119200 79654 120000
rect 81070 119200 81126 120000
rect 82542 119200 82598 120000
rect 84014 119200 84070 120000
rect 85486 119200 85542 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89994 119200 90050 120000
rect 91466 119200 91522 120000
rect 92938 119200 92994 120000
rect 94410 119200 94466 120000
rect 95974 119200 96030 120000
rect 97446 119200 97502 120000
rect 98918 119200 98974 120000
rect 100390 119200 100446 120000
rect 101862 119200 101918 120000
rect 103334 119200 103390 120000
rect 104898 119200 104954 120000
rect 106370 119200 106426 120000
rect 107842 119200 107898 120000
rect 109314 119200 109370 120000
rect 110786 119200 110842 120000
rect 112350 119200 112406 120000
rect 113822 119200 113878 120000
rect 115294 119200 115350 120000
rect 116766 119200 116822 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122746 119200 122802 120000
rect 124218 119200 124274 120000
rect 125690 119200 125746 120000
rect 127162 119200 127218 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131670 119200 131726 120000
rect 133142 119200 133198 120000
rect 134614 119200 134670 120000
rect 136086 119200 136142 120000
rect 137558 119200 137614 120000
rect 139122 119200 139178 120000
rect 140594 119200 140650 120000
rect 142066 119200 142122 120000
rect 143538 119200 143594 120000
rect 145010 119200 145066 120000
rect 146574 119200 146630 120000
rect 148046 119200 148102 120000
rect 149518 119200 149574 120000
rect 150990 119200 151046 120000
rect 152462 119200 152518 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 156970 119200 157026 120000
rect 158442 119200 158498 120000
rect 159914 119200 159970 120000
rect 161386 119200 161442 120000
rect 162858 119200 162914 120000
rect 164422 119200 164478 120000
rect 165894 119200 165950 120000
rect 167366 119200 167422 120000
rect 168838 119200 168894 120000
rect 170310 119200 170366 120000
rect 171782 119200 171838 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61842 0 61898 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64050 0 64106 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68742 0 68798 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84198 0 84254 800
rect 84474 0 84530 800
rect 84842 0 84898 800
rect 85210 0 85266 800
rect 85578 0 85634 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87786 0 87842 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92386 0 92442 800
rect 92754 0 92810 800
rect 93122 0 93178 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95330 0 95386 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97814 0 97870 800
rect 98182 0 98238 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99286 0 99342 800
rect 99654 0 99710 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112902 0 112958 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115018 0 115074 800
rect 115386 0 115442 800
rect 115754 0 115810 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122654 0 122710 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125874 0 125930 800
rect 126242 0 126298 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131578 0 131634 800
rect 131946 0 132002 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136270 0 136326 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137742 0 137798 800
rect 138018 0 138074 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141330 0 141386 800
rect 141698 0 141754 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146666 0 146722 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152094 0 152150 800
rect 152462 0 152518 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153474 0 153530 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159638 0 159694 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160742 0 160798 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 164974 0 165030 800
rect 165342 0 165398 800
rect 165710 0 165766 800
rect 166078 0 166134 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167918 0 167974 800
rect 168286 0 168342 800
rect 168654 0 168710 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 170034 0 170090 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171138 0 171194 800
rect 171506 0 171562 800
rect 171874 0 171930 800
rect 172242 0 172298 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6586 119354
rect 6754 119144 8058 119354
rect 8226 119144 9622 119354
rect 9790 119144 11094 119354
rect 11262 119144 12566 119354
rect 12734 119144 14038 119354
rect 14206 119144 15510 119354
rect 15678 119144 16982 119354
rect 17150 119144 18546 119354
rect 18714 119144 20018 119354
rect 20186 119144 21490 119354
rect 21658 119144 22962 119354
rect 23130 119144 24434 119354
rect 24602 119144 25906 119354
rect 26074 119144 27470 119354
rect 27638 119144 28942 119354
rect 29110 119144 30414 119354
rect 30582 119144 31886 119354
rect 32054 119144 33358 119354
rect 33526 119144 34830 119354
rect 34998 119144 36394 119354
rect 36562 119144 37866 119354
rect 38034 119144 39338 119354
rect 39506 119144 40810 119354
rect 40978 119144 42282 119354
rect 42450 119144 43846 119354
rect 44014 119144 45318 119354
rect 45486 119144 46790 119354
rect 46958 119144 48262 119354
rect 48430 119144 49734 119354
rect 49902 119144 51206 119354
rect 51374 119144 52770 119354
rect 52938 119144 54242 119354
rect 54410 119144 55714 119354
rect 55882 119144 57186 119354
rect 57354 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61694 119354
rect 61862 119144 63166 119354
rect 63334 119144 64638 119354
rect 64806 119144 66110 119354
rect 66278 119144 67582 119354
rect 67750 119144 69054 119354
rect 69222 119144 70618 119354
rect 70786 119144 72090 119354
rect 72258 119144 73562 119354
rect 73730 119144 75034 119354
rect 75202 119144 76506 119354
rect 76674 119144 78070 119354
rect 78238 119144 79542 119354
rect 79710 119144 81014 119354
rect 81182 119144 82486 119354
rect 82654 119144 83958 119354
rect 84126 119144 85430 119354
rect 85598 119144 86994 119354
rect 87162 119144 88466 119354
rect 88634 119144 89938 119354
rect 90106 119144 91410 119354
rect 91578 119144 92882 119354
rect 93050 119144 94354 119354
rect 94522 119144 95918 119354
rect 96086 119144 97390 119354
rect 97558 119144 98862 119354
rect 99030 119144 100334 119354
rect 100502 119144 101806 119354
rect 101974 119144 103278 119354
rect 103446 119144 104842 119354
rect 105010 119144 106314 119354
rect 106482 119144 107786 119354
rect 107954 119144 109258 119354
rect 109426 119144 110730 119354
rect 110898 119144 112294 119354
rect 112462 119144 113766 119354
rect 113934 119144 115238 119354
rect 115406 119144 116710 119354
rect 116878 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121218 119354
rect 121386 119144 122690 119354
rect 122858 119144 124162 119354
rect 124330 119144 125634 119354
rect 125802 119144 127106 119354
rect 127274 119144 128578 119354
rect 128746 119144 130142 119354
rect 130310 119144 131614 119354
rect 131782 119144 133086 119354
rect 133254 119144 134558 119354
rect 134726 119144 136030 119354
rect 136198 119144 137502 119354
rect 137670 119144 139066 119354
rect 139234 119144 140538 119354
rect 140706 119144 142010 119354
rect 142178 119144 143482 119354
rect 143650 119144 144954 119354
rect 145122 119144 146518 119354
rect 146686 119144 147990 119354
rect 148158 119144 149462 119354
rect 149630 119144 150934 119354
rect 151102 119144 152406 119354
rect 152574 119144 153878 119354
rect 154046 119144 155442 119354
rect 155610 119144 156914 119354
rect 157082 119144 158386 119354
rect 158554 119144 159858 119354
rect 160026 119144 161330 119354
rect 161498 119144 162802 119354
rect 162970 119144 164366 119354
rect 164534 119144 165838 119354
rect 166006 119144 167310 119354
rect 167478 119144 168782 119354
rect 168950 119144 170254 119354
rect 170422 119144 171726 119354
rect 171894 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 3918 856
rect 4086 734 4286 856
rect 4454 734 4654 856
rect 4822 734 5022 856
rect 5190 734 5390 856
rect 5558 734 5758 856
rect 5926 734 6126 856
rect 6294 734 6494 856
rect 6662 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7874 856
rect 8042 734 8242 856
rect 8410 734 8610 856
rect 8778 734 8978 856
rect 9146 734 9346 856
rect 9514 734 9714 856
rect 9882 734 10082 856
rect 10250 734 10450 856
rect 10618 734 10818 856
rect 10986 734 11186 856
rect 11354 734 11462 856
rect 11630 734 11830 856
rect 11998 734 12198 856
rect 12366 734 12566 856
rect 12734 734 12934 856
rect 13102 734 13302 856
rect 13470 734 13670 856
rect 13838 734 14038 856
rect 14206 734 14406 856
rect 14574 734 14774 856
rect 14942 734 15142 856
rect 15310 734 15418 856
rect 15586 734 15786 856
rect 15954 734 16154 856
rect 16322 734 16522 856
rect 16690 734 16890 856
rect 17058 734 17258 856
rect 17426 734 17626 856
rect 17794 734 17994 856
rect 18162 734 18362 856
rect 18530 734 18730 856
rect 18898 734 19098 856
rect 19266 734 19374 856
rect 19542 734 19742 856
rect 19910 734 20110 856
rect 20278 734 20478 856
rect 20646 734 20846 856
rect 21014 734 21214 856
rect 21382 734 21582 856
rect 21750 734 21950 856
rect 22118 734 22318 856
rect 22486 734 22686 856
rect 22854 734 22962 856
rect 23130 734 23330 856
rect 23498 734 23698 856
rect 23866 734 24066 856
rect 24234 734 24434 856
rect 24602 734 24802 856
rect 24970 734 25170 856
rect 25338 734 25538 856
rect 25706 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 26918 856
rect 27086 734 27286 856
rect 27454 734 27654 856
rect 27822 734 28022 856
rect 28190 734 28390 856
rect 28558 734 28758 856
rect 28926 734 29126 856
rect 29294 734 29494 856
rect 29662 734 29862 856
rect 30030 734 30230 856
rect 30398 734 30598 856
rect 30766 734 30874 856
rect 31042 734 31242 856
rect 31410 734 31610 856
rect 31778 734 31978 856
rect 32146 734 32346 856
rect 32514 734 32714 856
rect 32882 734 33082 856
rect 33250 734 33450 856
rect 33618 734 33818 856
rect 33986 734 34186 856
rect 34354 734 34462 856
rect 34630 734 34830 856
rect 34998 734 35198 856
rect 35366 734 35566 856
rect 35734 734 35934 856
rect 36102 734 36302 856
rect 36470 734 36670 856
rect 36838 734 37038 856
rect 37206 734 37406 856
rect 37574 734 37774 856
rect 37942 734 38142 856
rect 38310 734 38418 856
rect 38586 734 38786 856
rect 38954 734 39154 856
rect 39322 734 39522 856
rect 39690 734 39890 856
rect 40058 734 40258 856
rect 40426 734 40626 856
rect 40794 734 40994 856
rect 41162 734 41362 856
rect 41530 734 41730 856
rect 41898 734 42098 856
rect 42266 734 42374 856
rect 42542 734 42742 856
rect 42910 734 43110 856
rect 43278 734 43478 856
rect 43646 734 43846 856
rect 44014 734 44214 856
rect 44382 734 44582 856
rect 44750 734 44950 856
rect 45118 734 45318 856
rect 45486 734 45686 856
rect 45854 734 45962 856
rect 46130 734 46330 856
rect 46498 734 46698 856
rect 46866 734 47066 856
rect 47234 734 47434 856
rect 47602 734 47802 856
rect 47970 734 48170 856
rect 48338 734 48538 856
rect 48706 734 48906 856
rect 49074 734 49274 856
rect 49442 734 49642 856
rect 49810 734 49918 856
rect 50086 734 50286 856
rect 50454 734 50654 856
rect 50822 734 51022 856
rect 51190 734 51390 856
rect 51558 734 51758 856
rect 51926 734 52126 856
rect 52294 734 52494 856
rect 52662 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53874 856
rect 54042 734 54242 856
rect 54410 734 54610 856
rect 54778 734 54978 856
rect 55146 734 55346 856
rect 55514 734 55714 856
rect 55882 734 56082 856
rect 56250 734 56450 856
rect 56618 734 56818 856
rect 56986 734 57186 856
rect 57354 734 57462 856
rect 57630 734 57830 856
rect 57998 734 58198 856
rect 58366 734 58566 856
rect 58734 734 58934 856
rect 59102 734 59302 856
rect 59470 734 59670 856
rect 59838 734 60038 856
rect 60206 734 60406 856
rect 60574 734 60774 856
rect 60942 734 61142 856
rect 61310 734 61418 856
rect 61586 734 61786 856
rect 61954 734 62154 856
rect 62322 734 62522 856
rect 62690 734 62890 856
rect 63058 734 63258 856
rect 63426 734 63626 856
rect 63794 734 63994 856
rect 64162 734 64362 856
rect 64530 734 64730 856
rect 64898 734 65098 856
rect 65266 734 65374 856
rect 65542 734 65742 856
rect 65910 734 66110 856
rect 66278 734 66478 856
rect 66646 734 66846 856
rect 67014 734 67214 856
rect 67382 734 67582 856
rect 67750 734 67950 856
rect 68118 734 68318 856
rect 68486 734 68686 856
rect 68854 734 68962 856
rect 69130 734 69330 856
rect 69498 734 69698 856
rect 69866 734 70066 856
rect 70234 734 70434 856
rect 70602 734 70802 856
rect 70970 734 71170 856
rect 71338 734 71538 856
rect 71706 734 71906 856
rect 72074 734 72274 856
rect 72442 734 72642 856
rect 72810 734 72918 856
rect 73086 734 73286 856
rect 73454 734 73654 856
rect 73822 734 74022 856
rect 74190 734 74390 856
rect 74558 734 74758 856
rect 74926 734 75126 856
rect 75294 734 75494 856
rect 75662 734 75862 856
rect 76030 734 76230 856
rect 76398 734 76598 856
rect 76766 734 76874 856
rect 77042 734 77242 856
rect 77410 734 77610 856
rect 77778 734 77978 856
rect 78146 734 78346 856
rect 78514 734 78714 856
rect 78882 734 79082 856
rect 79250 734 79450 856
rect 79618 734 79818 856
rect 79986 734 80186 856
rect 80354 734 80462 856
rect 80630 734 80830 856
rect 80998 734 81198 856
rect 81366 734 81566 856
rect 81734 734 81934 856
rect 82102 734 82302 856
rect 82470 734 82670 856
rect 82838 734 83038 856
rect 83206 734 83406 856
rect 83574 734 83774 856
rect 83942 734 84142 856
rect 84310 734 84418 856
rect 84586 734 84786 856
rect 84954 734 85154 856
rect 85322 734 85522 856
rect 85690 734 85890 856
rect 86058 734 86258 856
rect 86426 734 86626 856
rect 86794 734 86994 856
rect 87162 734 87362 856
rect 87530 734 87730 856
rect 87898 734 88098 856
rect 88266 734 88374 856
rect 88542 734 88742 856
rect 88910 734 89110 856
rect 89278 734 89478 856
rect 89646 734 89846 856
rect 90014 734 90214 856
rect 90382 734 90582 856
rect 90750 734 90950 856
rect 91118 734 91318 856
rect 91486 734 91686 856
rect 91854 734 91962 856
rect 92130 734 92330 856
rect 92498 734 92698 856
rect 92866 734 93066 856
rect 93234 734 93434 856
rect 93602 734 93802 856
rect 93970 734 94170 856
rect 94338 734 94538 856
rect 94706 734 94906 856
rect 95074 734 95274 856
rect 95442 734 95642 856
rect 95810 734 95918 856
rect 96086 734 96286 856
rect 96454 734 96654 856
rect 96822 734 97022 856
rect 97190 734 97390 856
rect 97558 734 97758 856
rect 97926 734 98126 856
rect 98294 734 98494 856
rect 98662 734 98862 856
rect 99030 734 99230 856
rect 99398 734 99598 856
rect 99766 734 99874 856
rect 100042 734 100242 856
rect 100410 734 100610 856
rect 100778 734 100978 856
rect 101146 734 101346 856
rect 101514 734 101714 856
rect 101882 734 102082 856
rect 102250 734 102450 856
rect 102618 734 102818 856
rect 102986 734 103186 856
rect 103354 734 103462 856
rect 103630 734 103830 856
rect 103998 734 104198 856
rect 104366 734 104566 856
rect 104734 734 104934 856
rect 105102 734 105302 856
rect 105470 734 105670 856
rect 105838 734 106038 856
rect 106206 734 106406 856
rect 106574 734 106774 856
rect 106942 734 107142 856
rect 107310 734 107418 856
rect 107586 734 107786 856
rect 107954 734 108154 856
rect 108322 734 108522 856
rect 108690 734 108890 856
rect 109058 734 109258 856
rect 109426 734 109626 856
rect 109794 734 109994 856
rect 110162 734 110362 856
rect 110530 734 110730 856
rect 110898 734 111098 856
rect 111266 734 111374 856
rect 111542 734 111742 856
rect 111910 734 112110 856
rect 112278 734 112478 856
rect 112646 734 112846 856
rect 113014 734 113214 856
rect 113382 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114318 856
rect 114486 734 114686 856
rect 114854 734 114962 856
rect 115130 734 115330 856
rect 115498 734 115698 856
rect 115866 734 116066 856
rect 116234 734 116434 856
rect 116602 734 116802 856
rect 116970 734 117170 856
rect 117338 734 117538 856
rect 117706 734 117906 856
rect 118074 734 118274 856
rect 118442 734 118642 856
rect 118810 734 118918 856
rect 119086 734 119286 856
rect 119454 734 119654 856
rect 119822 734 120022 856
rect 120190 734 120390 856
rect 120558 734 120758 856
rect 120926 734 121126 856
rect 121294 734 121494 856
rect 121662 734 121862 856
rect 122030 734 122230 856
rect 122398 734 122598 856
rect 122766 734 122874 856
rect 123042 734 123242 856
rect 123410 734 123610 856
rect 123778 734 123978 856
rect 124146 734 124346 856
rect 124514 734 124714 856
rect 124882 734 125082 856
rect 125250 734 125450 856
rect 125618 734 125818 856
rect 125986 734 126186 856
rect 126354 734 126462 856
rect 126630 734 126830 856
rect 126998 734 127198 856
rect 127366 734 127566 856
rect 127734 734 127934 856
rect 128102 734 128302 856
rect 128470 734 128670 856
rect 128838 734 129038 856
rect 129206 734 129406 856
rect 129574 734 129774 856
rect 129942 734 130142 856
rect 130310 734 130418 856
rect 130586 734 130786 856
rect 130954 734 131154 856
rect 131322 734 131522 856
rect 131690 734 131890 856
rect 132058 734 132258 856
rect 132426 734 132626 856
rect 132794 734 132994 856
rect 133162 734 133362 856
rect 133530 734 133730 856
rect 133898 734 134098 856
rect 134266 734 134374 856
rect 134542 734 134742 856
rect 134910 734 135110 856
rect 135278 734 135478 856
rect 135646 734 135846 856
rect 136014 734 136214 856
rect 136382 734 136582 856
rect 136750 734 136950 856
rect 137118 734 137318 856
rect 137486 734 137686 856
rect 137854 734 137962 856
rect 138130 734 138330 856
rect 138498 734 138698 856
rect 138866 734 139066 856
rect 139234 734 139434 856
rect 139602 734 139802 856
rect 139970 734 140170 856
rect 140338 734 140538 856
rect 140706 734 140906 856
rect 141074 734 141274 856
rect 141442 734 141642 856
rect 141810 734 141918 856
rect 142086 734 142286 856
rect 142454 734 142654 856
rect 142822 734 143022 856
rect 143190 734 143390 856
rect 143558 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144494 856
rect 144662 734 144862 856
rect 145030 734 145230 856
rect 145398 734 145598 856
rect 145766 734 145874 856
rect 146042 734 146242 856
rect 146410 734 146610 856
rect 146778 734 146978 856
rect 147146 734 147346 856
rect 147514 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148450 856
rect 148618 734 148818 856
rect 148986 734 149186 856
rect 149354 734 149462 856
rect 149630 734 149830 856
rect 149998 734 150198 856
rect 150366 734 150566 856
rect 150734 734 150934 856
rect 151102 734 151302 856
rect 151470 734 151670 856
rect 151838 734 152038 856
rect 152206 734 152406 856
rect 152574 734 152774 856
rect 152942 734 153142 856
rect 153310 734 153418 856
rect 153586 734 153786 856
rect 153954 734 154154 856
rect 154322 734 154522 856
rect 154690 734 154890 856
rect 155058 734 155258 856
rect 155426 734 155626 856
rect 155794 734 155994 856
rect 156162 734 156362 856
rect 156530 734 156730 856
rect 156898 734 157098 856
rect 157266 734 157374 856
rect 157542 734 157742 856
rect 157910 734 158110 856
rect 158278 734 158478 856
rect 158646 734 158846 856
rect 159014 734 159214 856
rect 159382 734 159582 856
rect 159750 734 159950 856
rect 160118 734 160318 856
rect 160486 734 160686 856
rect 160854 734 160962 856
rect 161130 734 161330 856
rect 161498 734 161698 856
rect 161866 734 162066 856
rect 162234 734 162434 856
rect 162602 734 162802 856
rect 162970 734 163170 856
rect 163338 734 163538 856
rect 163706 734 163906 856
rect 164074 734 164274 856
rect 164442 734 164642 856
rect 164810 734 164918 856
rect 165086 734 165286 856
rect 165454 734 165654 856
rect 165822 734 166022 856
rect 166190 734 166390 856
rect 166558 734 166758 856
rect 166926 734 167126 856
rect 167294 734 167494 856
rect 167662 734 167862 856
rect 168030 734 168230 856
rect 168398 734 168598 856
rect 168766 734 168874 856
rect 169042 734 169242 856
rect 169410 734 169610 856
rect 169778 734 169978 856
rect 170146 734 170346 856
rect 170514 734 170714 856
rect 170882 734 171082 856
rect 171250 734 171450 856
rect 171618 734 171818 856
rect 171986 734 172186 856
rect 172354 734 172462 856
rect 172630 734 172830 856
rect 172998 734 173198 856
rect 173366 734 173566 856
rect 173734 734 173934 856
rect 174102 734 174302 856
rect 174470 734 174670 856
rect 174838 734 175038 856
rect 175206 734 175406 856
rect 175574 734 175774 856
rect 175942 734 176142 856
rect 176310 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178186 856
<< metal3 >>
rect 179200 112344 180000 112464
rect 0 111392 800 111512
rect 179200 97384 180000 97504
rect 0 94256 800 94376
rect 179200 82424 180000 82544
rect 0 77120 800 77240
rect 179200 67464 180000 67584
rect 0 59984 800 60104
rect 179200 52368 180000 52488
rect 0 42848 800 42968
rect 179200 37408 180000 37528
rect 0 25712 800 25832
rect 179200 22448 180000 22568
rect 0 8576 800 8696
rect 179200 7488 180000 7608
<< obsm3 >>
rect 4208 112544 179200 117537
rect 4208 112264 179120 112544
rect 4208 97584 179200 112264
rect 4208 97304 179120 97584
rect 4208 82624 179200 97304
rect 4208 82344 179120 82624
rect 4208 67664 179200 82344
rect 4208 67384 179120 67664
rect 4208 52568 179200 67384
rect 4208 52288 179120 52568
rect 4208 37608 179200 52288
rect 4208 37328 179120 37608
rect 4208 22648 179200 37328
rect 4208 22368 179120 22648
rect 4208 7688 179200 22368
rect 4208 7408 179120 7688
rect 4208 2143 179200 7408
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 77155 112915 80165 117197
<< labels >>
rlabel metal2 s 176198 0 176254 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 42848 800 42968 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 179200 67464 180000 67584 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 77120 800 77240 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 179200 82424 180000 82544 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 94256 800 94376 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 176474 0 176530 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 111392 800 111512 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 179200 97384 180000 97504 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 179200 112344 180000 112464 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 176842 0 176898 800 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 0 8576 800 8696 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 179200 37408 180000 37528 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 179200 52368 180000 52488 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 171782 119200 171838 120000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 0 25712 800 25832 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 45374 119200 45430 120000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 49790 119200 49846 120000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 54298 119200 54354 120000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 58714 119200 58770 120000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 63222 119200 63278 120000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 67638 119200 67694 120000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 81070 119200 81126 120000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 85486 119200 85542 120000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 89994 119200 90050 120000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 94410 119200 94466 120000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 98918 119200 98974 120000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 103334 119200 103390 120000 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 107842 119200 107898 120000 6 io_in[24]
port 46 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 116766 119200 116822 120000 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 121274 119200 121330 120000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 125690 119200 125746 120000 6 io_in[28]
port 50 nsew signal input
rlabel metal2 s 130198 119200 130254 120000 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 io_in[32]
port 55 nsew signal input
rlabel metal2 s 148046 119200 148102 120000 6 io_in[33]
port 56 nsew signal input
rlabel metal2 s 152462 119200 152518 120000 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 156970 119200 157026 120000 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 161386 119200 161442 120000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 165894 119200 165950 120000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 14094 119200 14150 120000 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 18602 119200 18658 120000 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 23018 119200 23074 120000 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 27526 119200 27582 120000 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 31942 119200 31998 120000 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 36450 119200 36506 120000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 40866 119200 40922 120000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 46846 119200 46902 120000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 69110 119200 69166 120000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 73618 119200 73674 120000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 95974 119200 96030 120000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 100390 119200 100446 120000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 104898 119200 104954 120000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal2 s 109314 119200 109370 120000 6 io_oeb[24]
port 84 nsew signal output
rlabel metal2 s 113822 119200 113878 120000 6 io_oeb[25]
port 85 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 122746 119200 122802 120000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 127162 119200 127218 120000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal2 s 131670 119200 131726 120000 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 11150 119200 11206 120000 6 io_oeb[2]
port 90 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 140594 119200 140650 120000 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 145010 119200 145066 120000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal2 s 149518 119200 149574 120000 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 158442 119200 158498 120000 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 162858 119200 162914 120000 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 15566 119200 15622 120000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 33414 119200 33470 120000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 37922 119200 37978 120000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 42338 119200 42394 120000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 48318 119200 48374 120000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 57242 119200 57298 120000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 61750 119200 61806 120000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 66166 119200 66222 120000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 84014 119200 84070 120000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 92938 119200 92994 120000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 101862 119200 101918 120000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_out[23]
port 121 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 128634 119200 128690 120000 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 133142 119200 133198 120000 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 12622 119200 12678 120000 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 137558 119200 137614 120000 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 142066 119200 142122 120000 6 io_out[31]
port 130 nsew signal output
rlabel metal2 s 146574 119200 146630 120000 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 150990 119200 151046 120000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 159914 119200 159970 120000 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 164422 119200 164478 120000 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 168838 119200 168894 120000 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 17038 119200 17094 120000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 21546 119200 21602 120000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 43902 119200 43958 120000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 131946 0 132002 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 154946 0 155002 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 157154 0 157210 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 158166 0 158222 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 63314 0 63370 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 144182 0 144238 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 170310 119200 170366 120000 6 user_clock2
port 528 nsew signal input
rlabel metal3 s 179200 7488 180000 7608 6 user_irq[0]
port 529 nsew signal output
rlabel metal3 s 179200 22448 180000 22568 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 532 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 533 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 533 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7624250
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_four.magic.gds
string GDS_START 217786
<< end >>

