VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.190 1421.780 1114.510 1421.840 ;
        RECT 2898.990 1421.780 2899.310 1421.840 ;
        RECT 1114.190 1421.640 2899.310 1421.780 ;
        RECT 1114.190 1421.580 1114.510 1421.640 ;
        RECT 2898.990 1421.580 2899.310 1421.640 ;
      LAYER via ;
        RECT 1114.220 1421.580 1114.480 1421.840 ;
        RECT 2899.020 1421.580 2899.280 1421.840 ;
      LAYER met2 ;
        RECT 2899.010 1426.795 2899.290 1427.165 ;
        RECT 2899.080 1421.870 2899.220 1426.795 ;
        RECT 1114.220 1421.550 1114.480 1421.870 ;
        RECT 2899.020 1421.550 2899.280 1421.870 ;
        RECT 1114.280 492.845 1114.420 1421.550 ;
        RECT 1114.210 492.475 1114.490 492.845 ;
      LAYER via2 ;
        RECT 2899.010 1426.840 2899.290 1427.120 ;
        RECT 1114.210 492.520 1114.490 492.800 ;
      LAYER met3 ;
        RECT 2898.985 1427.130 2899.315 1427.145 ;
        RECT 2917.600 1427.130 2924.800 1427.580 ;
        RECT 2898.985 1426.830 2924.800 1427.130 ;
        RECT 2898.985 1426.815 2899.315 1426.830 ;
        RECT 2917.600 1426.380 2924.800 1426.830 ;
        RECT 1114.185 492.810 1114.515 492.825 ;
        RECT 1098.790 492.510 1114.515 492.810 ;
        RECT 1098.790 490.400 1099.090 492.510 ;
        RECT 1114.185 492.495 1114.515 492.510 ;
        RECT 1096.000 489.800 1100.000 490.400 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1048.410 1010.720 1048.730 1010.780 ;
        RECT 2228.770 1010.720 2229.090 1010.780 ;
        RECT 1048.410 1010.580 2229.090 1010.720 ;
        RECT 1048.410 1010.520 1048.730 1010.580 ;
        RECT 2228.770 1010.520 2229.090 1010.580 ;
      LAYER via ;
        RECT 1048.440 1010.520 1048.700 1010.780 ;
        RECT 2228.800 1010.520 2229.060 1010.780 ;
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
        RECT 2230.700 3512.170 2230.840 3517.600 ;
        RECT 2228.860 3512.030 2230.840 3512.170 ;
        RECT 2228.860 1010.810 2229.000 3512.030 ;
        RECT 1048.440 1010.490 1048.700 1010.810 ;
        RECT 2228.800 1010.490 2229.060 1010.810 ;
        RECT 1046.490 999.330 1046.770 1000.000 ;
        RECT 1048.500 999.330 1048.640 1010.490 ;
        RECT 1046.490 999.190 1048.640 999.330 ;
        RECT 1046.490 996.000 1046.770 999.190 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.310 1011.060 1055.630 1011.120 ;
        RECT 1904.470 1011.060 1904.790 1011.120 ;
        RECT 1055.310 1010.920 1904.790 1011.060 ;
        RECT 1055.310 1010.860 1055.630 1010.920 ;
        RECT 1904.470 1010.860 1904.790 1010.920 ;
      LAYER via ;
        RECT 1055.340 1010.860 1055.600 1011.120 ;
        RECT 1904.500 1010.860 1904.760 1011.120 ;
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
        RECT 1905.940 3512.170 1906.080 3517.600 ;
        RECT 1904.560 3512.030 1906.080 3512.170 ;
        RECT 1904.560 1011.150 1904.700 3512.030 ;
        RECT 1055.340 1010.830 1055.600 1011.150 ;
        RECT 1904.500 1010.830 1904.760 1011.150 ;
        RECT 1053.850 999.330 1054.130 1000.000 ;
        RECT 1055.400 999.330 1055.540 1010.830 ;
        RECT 1053.850 999.190 1055.540 999.330 ;
        RECT 1053.850 996.000 1054.130 999.190 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 909.030 998.140 909.350 998.200 ;
        RECT 869.330 998.000 909.350 998.140 ;
        RECT 191.430 997.800 191.750 997.860 ;
        RECT 191.430 997.660 276.070 997.800 ;
        RECT 191.430 997.600 191.750 997.660 ;
        RECT 275.930 997.120 276.070 997.660 ;
        RECT 469.130 997.660 517.570 997.800 ;
        RECT 469.130 997.120 469.270 997.660 ;
        RECT 275.930 996.980 469.270 997.120 ;
        RECT 517.430 997.120 517.570 997.660 ;
        RECT 869.330 997.120 869.470 998.000 ;
        RECT 909.030 997.940 909.350 998.000 ;
        RECT 909.030 997.460 909.350 997.520 ;
        RECT 909.030 997.320 917.770 997.460 ;
        RECT 909.030 997.260 909.350 997.320 ;
        RECT 517.430 996.980 869.470 997.120 ;
        RECT 917.630 997.120 917.770 997.320 ;
        RECT 1580.170 997.120 1580.490 997.180 ;
        RECT 917.630 996.980 1580.490 997.120 ;
        RECT 1580.170 996.920 1580.490 996.980 ;
      LAYER via ;
        RECT 191.460 997.600 191.720 997.860 ;
        RECT 909.060 997.940 909.320 998.200 ;
        RECT 909.060 997.260 909.320 997.520 ;
        RECT 1580.200 996.920 1580.460 997.180 ;
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
        RECT 1581.640 3512.170 1581.780 3517.600 ;
        RECT 1580.260 3512.030 1581.780 3512.170 ;
        RECT 909.060 997.910 909.320 998.230 ;
        RECT 191.460 997.570 191.720 997.890 ;
        RECT 191.520 702.965 191.660 997.570 ;
        RECT 909.120 997.550 909.260 997.910 ;
        RECT 909.060 997.230 909.320 997.550 ;
        RECT 1580.260 997.210 1580.400 3512.030 ;
        RECT 1580.200 996.890 1580.460 997.210 ;
        RECT 191.450 702.595 191.730 702.965 ;
      LAYER via2 ;
        RECT 191.450 702.640 191.730 702.920 ;
      LAYER met3 ;
        RECT 191.425 702.930 191.755 702.945 ;
        RECT 191.425 702.630 201.170 702.930 ;
        RECT 191.425 702.615 191.755 702.630 ;
        RECT 200.870 700.520 201.170 702.630 ;
        RECT 200.000 699.920 204.000 700.520 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1097.170 393.620 1097.490 393.680 ;
        RECT 1255.870 393.620 1256.190 393.680 ;
        RECT 1097.170 393.480 1256.190 393.620 ;
        RECT 1097.170 393.420 1097.490 393.480 ;
        RECT 1255.870 393.420 1256.190 393.480 ;
      LAYER via ;
        RECT 1097.200 393.420 1097.460 393.680 ;
        RECT 1255.900 393.420 1256.160 393.680 ;
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
        RECT 1257.340 3512.170 1257.480 3517.600 ;
        RECT 1255.960 3512.030 1257.480 3512.170 ;
        RECT 1097.090 400.180 1097.370 404.000 ;
        RECT 1097.090 400.000 1097.400 400.180 ;
        RECT 1097.260 393.710 1097.400 400.000 ;
        RECT 1255.960 393.710 1256.100 3512.030 ;
        RECT 1097.200 393.390 1097.460 393.710 ;
        RECT 1255.900 393.390 1256.160 393.710 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 997.460 931.890 997.520 ;
        RECT 1111.890 997.460 1112.210 997.520 ;
        RECT 931.570 997.320 1112.210 997.460 ;
        RECT 931.570 997.260 931.890 997.320 ;
        RECT 1111.890 997.260 1112.210 997.320 ;
      LAYER via ;
        RECT 931.600 997.260 931.860 997.520 ;
        RECT 1111.920 997.260 1112.180 997.520 ;
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
        RECT 932.580 3415.570 932.720 3517.600 ;
        RECT 932.120 3415.430 932.720 3415.570 ;
        RECT 932.120 1048.870 932.260 3415.430 ;
        RECT 931.660 1048.730 932.260 1048.870 ;
        RECT 931.660 997.550 931.800 1048.730 ;
        RECT 931.600 997.230 931.860 997.550 ;
        RECT 1111.920 997.230 1112.180 997.550 ;
        RECT 1111.980 731.525 1112.120 997.230 ;
        RECT 1111.910 731.155 1112.190 731.525 ;
      LAYER via2 ;
        RECT 1111.910 731.200 1112.190 731.480 ;
      LAYER met3 ;
        RECT 1111.885 731.490 1112.215 731.505 ;
        RECT 1098.790 731.190 1112.215 731.490 ;
        RECT 1098.790 730.440 1099.090 731.190 ;
        RECT 1111.885 731.175 1112.215 731.190 ;
        RECT 1096.000 729.840 1100.000 730.440 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.810 3504.280 193.130 3504.340 ;
        RECT 608.190 3504.280 608.510 3504.340 ;
        RECT 192.810 3504.140 608.510 3504.280 ;
        RECT 192.810 3504.080 193.130 3504.140 ;
        RECT 608.190 3504.080 608.510 3504.140 ;
      LAYER via ;
        RECT 192.840 3504.080 193.100 3504.340 ;
        RECT 608.220 3504.080 608.480 3504.340 ;
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
        RECT 608.280 3504.370 608.420 3517.600 ;
        RECT 192.840 3504.050 193.100 3504.370 ;
        RECT 608.220 3504.050 608.480 3504.370 ;
        RECT 192.900 785.245 193.040 3504.050 ;
        RECT 192.830 784.875 193.110 785.245 ;
      LAYER via2 ;
        RECT 192.830 784.920 193.110 785.200 ;
      LAYER met3 ;
        RECT 200.000 785.600 204.000 786.200 ;
        RECT 192.805 785.210 193.135 785.225 ;
        RECT 200.870 785.210 201.170 785.600 ;
        RECT 192.805 784.910 201.170 785.210 ;
        RECT 192.805 784.895 193.135 784.910 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.350 3501.900 192.670 3501.960 ;
        RECT 283.890 3501.900 284.210 3501.960 ;
        RECT 192.350 3501.760 284.210 3501.900 ;
        RECT 192.350 3501.700 192.670 3501.760 ;
        RECT 283.890 3501.700 284.210 3501.760 ;
      LAYER via ;
        RECT 192.380 3501.700 192.640 3501.960 ;
        RECT 283.920 3501.700 284.180 3501.960 ;
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
        RECT 283.980 3501.990 284.120 3517.600 ;
        RECT 192.380 3501.670 192.640 3501.990 ;
        RECT 283.920 3501.670 284.180 3501.990 ;
        RECT 192.440 874.325 192.580 3501.670 ;
        RECT 192.370 873.955 192.650 874.325 ;
      LAYER via2 ;
        RECT 192.370 874.000 192.650 874.280 ;
      LAYER met3 ;
        RECT 192.345 874.290 192.675 874.305 ;
        RECT 192.345 873.990 201.170 874.290 ;
        RECT 192.345 873.975 192.675 873.990 ;
        RECT 200.870 871.880 201.170 873.990 ;
        RECT 200.000 871.280 204.000 871.880 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 3485.240 16.950 3485.300 ;
        RECT 1110.970 3485.240 1111.290 3485.300 ;
        RECT 16.630 3485.100 1111.290 3485.240 ;
        RECT 16.630 3485.040 16.950 3485.100 ;
        RECT 1110.970 3485.040 1111.290 3485.100 ;
      LAYER via ;
        RECT 16.660 3485.040 16.920 3485.300 ;
        RECT 1111.000 3485.040 1111.260 3485.300 ;
      LAYER met2 ;
        RECT 16.650 3486.515 16.930 3486.885 ;
        RECT 16.720 3485.330 16.860 3486.515 ;
        RECT 16.660 3485.010 16.920 3485.330 ;
        RECT 1111.000 3485.010 1111.260 3485.330 ;
        RECT 1111.060 792.725 1111.200 3485.010 ;
        RECT 1110.990 792.355 1111.270 792.725 ;
      LAYER via2 ;
        RECT 16.650 3486.560 16.930 3486.840 ;
        RECT 1110.990 792.400 1111.270 792.680 ;
      LAYER met3 ;
        RECT -4.800 3486.850 2.400 3487.300 ;
        RECT 16.625 3486.850 16.955 3486.865 ;
        RECT -4.800 3486.550 16.955 3486.850 ;
        RECT -4.800 3486.100 2.400 3486.550 ;
        RECT 16.625 3486.535 16.955 3486.550 ;
        RECT 1110.965 792.690 1111.295 792.705 ;
        RECT 1098.790 792.390 1111.295 792.690 ;
        RECT 1098.790 790.280 1099.090 792.390 ;
        RECT 1110.965 792.375 1111.295 792.390 ;
        RECT 1096.000 789.680 1100.000 790.280 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 3222.420 16.030 3222.480 ;
        RECT 948.590 3222.420 948.910 3222.480 ;
        RECT 15.710 3222.280 948.910 3222.420 ;
        RECT 15.710 3222.220 16.030 3222.280 ;
        RECT 948.590 3222.220 948.910 3222.280 ;
        RECT 948.590 1013.780 948.910 1013.840 ;
        RECT 1058.990 1013.780 1059.310 1013.840 ;
        RECT 948.590 1013.640 1059.310 1013.780 ;
        RECT 948.590 1013.580 948.910 1013.640 ;
        RECT 1058.990 1013.580 1059.310 1013.640 ;
      LAYER via ;
        RECT 15.740 3222.220 16.000 3222.480 ;
        RECT 948.620 3222.220 948.880 3222.480 ;
        RECT 948.620 1013.580 948.880 1013.840 ;
        RECT 1059.020 1013.580 1059.280 1013.840 ;
      LAYER met2 ;
        RECT 15.730 3225.395 16.010 3225.765 ;
        RECT 15.800 3222.510 15.940 3225.395 ;
        RECT 15.740 3222.190 16.000 3222.510 ;
        RECT 948.620 3222.190 948.880 3222.510 ;
        RECT 948.680 1013.870 948.820 3222.190 ;
        RECT 948.620 1013.550 948.880 1013.870 ;
        RECT 1059.020 1013.550 1059.280 1013.870 ;
        RECT 1059.080 999.330 1059.220 1013.550 ;
        RECT 1060.750 999.330 1061.030 1000.000 ;
        RECT 1059.080 999.190 1061.030 999.330 ;
        RECT 1060.750 996.000 1061.030 999.190 ;
      LAYER via2 ;
        RECT 15.730 3225.440 16.010 3225.720 ;
      LAYER met3 ;
        RECT -4.800 3225.730 2.400 3226.180 ;
        RECT 15.705 3225.730 16.035 3225.745 ;
        RECT -4.800 3225.430 16.035 3225.730 ;
        RECT -4.800 3224.980 2.400 3225.430 ;
        RECT 15.705 3225.415 16.035 3225.430 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2960.280 16.030 2960.340 ;
        RECT 914.090 2960.280 914.410 2960.340 ;
        RECT 15.710 2960.140 914.410 2960.280 ;
        RECT 15.710 2960.080 16.030 2960.140 ;
        RECT 914.090 2960.080 914.410 2960.140 ;
        RECT 914.090 1013.440 914.410 1013.500 ;
        RECT 1066.350 1013.440 1066.670 1013.500 ;
        RECT 914.090 1013.300 1066.670 1013.440 ;
        RECT 914.090 1013.240 914.410 1013.300 ;
        RECT 1066.350 1013.240 1066.670 1013.300 ;
      LAYER via ;
        RECT 15.740 2960.080 16.000 2960.340 ;
        RECT 914.120 2960.080 914.380 2960.340 ;
        RECT 914.120 1013.240 914.380 1013.500 ;
        RECT 1066.380 1013.240 1066.640 1013.500 ;
      LAYER met2 ;
        RECT 15.730 2964.955 16.010 2965.325 ;
        RECT 15.800 2960.370 15.940 2964.955 ;
        RECT 15.740 2960.050 16.000 2960.370 ;
        RECT 914.120 2960.050 914.380 2960.370 ;
        RECT 914.180 1013.530 914.320 2960.050 ;
        RECT 914.120 1013.210 914.380 1013.530 ;
        RECT 1066.380 1013.210 1066.640 1013.530 ;
        RECT 1066.440 999.330 1066.580 1013.210 ;
        RECT 1067.650 999.330 1067.930 1000.000 ;
        RECT 1066.440 999.190 1067.930 999.330 ;
        RECT 1067.650 996.000 1067.930 999.190 ;
      LAYER via2 ;
        RECT 15.730 2965.000 16.010 2965.280 ;
      LAYER met3 ;
        RECT -4.800 2965.290 2.400 2965.740 ;
        RECT 15.705 2965.290 16.035 2965.305 ;
        RECT -4.800 2964.990 16.035 2965.290 ;
        RECT -4.800 2964.540 2.400 2964.990 ;
        RECT 15.705 2964.975 16.035 2964.990 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.470 1690.720 1007.790 1690.780 ;
        RECT 2900.830 1690.720 2901.150 1690.780 ;
        RECT 1007.470 1690.580 2901.150 1690.720 ;
        RECT 1007.470 1690.520 1007.790 1690.580 ;
        RECT 2900.830 1690.520 2901.150 1690.580 ;
      LAYER via ;
        RECT 1007.500 1690.520 1007.760 1690.780 ;
        RECT 2900.860 1690.520 2901.120 1690.780 ;
      LAYER met2 ;
        RECT 2900.850 1692.675 2901.130 1693.045 ;
        RECT 2900.920 1690.810 2901.060 1692.675 ;
        RECT 1007.500 1690.490 1007.760 1690.810 ;
        RECT 2900.860 1690.490 2901.120 1690.810 ;
        RECT 1007.560 1048.870 1007.700 1690.490 ;
        RECT 1007.560 1048.730 1009.080 1048.870 ;
        RECT 1008.940 999.330 1009.080 1048.730 ;
        RECT 1011.070 999.330 1011.350 1000.000 ;
        RECT 1008.940 999.190 1011.350 999.330 ;
        RECT 1011.070 996.000 1011.350 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1692.720 2901.130 1693.000 ;
      LAYER met3 ;
        RECT 2900.825 1693.010 2901.155 1693.025 ;
        RECT 2917.600 1693.010 2924.800 1693.460 ;
        RECT 2900.825 1692.710 2924.800 1693.010 ;
        RECT 2900.825 1692.695 2901.155 1692.710 ;
        RECT 2917.600 1692.260 2924.800 1692.710 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2698.140 16.490 2698.200 ;
        RECT 920.990 2698.140 921.310 2698.200 ;
        RECT 16.170 2698.000 921.310 2698.140 ;
        RECT 16.170 2697.940 16.490 2698.000 ;
        RECT 920.990 2697.940 921.310 2698.000 ;
        RECT 920.990 1013.100 921.310 1013.160 ;
        RECT 1073.710 1013.100 1074.030 1013.160 ;
        RECT 920.990 1012.960 1074.030 1013.100 ;
        RECT 920.990 1012.900 921.310 1012.960 ;
        RECT 1073.710 1012.900 1074.030 1012.960 ;
      LAYER via ;
        RECT 16.200 2697.940 16.460 2698.200 ;
        RECT 921.020 2697.940 921.280 2698.200 ;
        RECT 921.020 1012.900 921.280 1013.160 ;
        RECT 1073.740 1012.900 1074.000 1013.160 ;
      LAYER met2 ;
        RECT 16.190 2703.835 16.470 2704.205 ;
        RECT 16.260 2698.230 16.400 2703.835 ;
        RECT 16.200 2697.910 16.460 2698.230 ;
        RECT 921.020 2697.910 921.280 2698.230 ;
        RECT 921.080 1013.190 921.220 2697.910 ;
        RECT 921.020 1012.870 921.280 1013.190 ;
        RECT 1073.740 1012.870 1074.000 1013.190 ;
        RECT 1073.800 999.330 1073.940 1012.870 ;
        RECT 1075.010 999.330 1075.290 1000.000 ;
        RECT 1073.800 999.190 1075.290 999.330 ;
        RECT 1075.010 996.000 1075.290 999.190 ;
      LAYER via2 ;
        RECT 16.190 2703.880 16.470 2704.160 ;
      LAYER met3 ;
        RECT -4.800 2704.170 2.400 2704.620 ;
        RECT 16.165 2704.170 16.495 2704.185 ;
        RECT -4.800 2703.870 16.495 2704.170 ;
        RECT -4.800 2703.420 2.400 2703.870 ;
        RECT 16.165 2703.855 16.495 2703.870 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2442.800 17.410 2442.860 ;
        RECT 1097.630 2442.800 1097.950 2442.860 ;
        RECT 17.090 2442.660 1097.950 2442.800 ;
        RECT 17.090 2442.600 17.410 2442.660 ;
        RECT 1097.630 2442.600 1097.950 2442.660 ;
      LAYER via ;
        RECT 17.120 2442.600 17.380 2442.860 ;
        RECT 1097.660 2442.600 1097.920 2442.860 ;
      LAYER met2 ;
        RECT 17.110 2443.395 17.390 2443.765 ;
        RECT 17.180 2442.890 17.320 2443.395 ;
        RECT 17.120 2442.570 17.380 2442.890 ;
        RECT 1097.660 2442.570 1097.920 2442.890 ;
        RECT 1097.720 403.650 1097.860 2442.570 ;
        RECT 1098.930 403.650 1099.210 404.000 ;
        RECT 1097.720 403.510 1099.210 403.650 ;
        RECT 1098.930 400.000 1099.210 403.510 ;
      LAYER via2 ;
        RECT 17.110 2443.440 17.390 2443.720 ;
      LAYER met3 ;
        RECT -4.800 2443.730 2.400 2444.180 ;
        RECT 17.085 2443.730 17.415 2443.745 ;
        RECT -4.800 2443.430 17.415 2443.730 ;
        RECT -4.800 2442.980 2.400 2443.430 ;
        RECT 17.085 2443.415 17.415 2443.430 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2180.660 17.870 2180.720 ;
        RECT 1111.430 2180.660 1111.750 2180.720 ;
        RECT 17.550 2180.520 1111.750 2180.660 ;
        RECT 17.550 2180.460 17.870 2180.520 ;
        RECT 1111.430 2180.460 1111.750 2180.520 ;
      LAYER via ;
        RECT 17.580 2180.460 17.840 2180.720 ;
        RECT 1111.460 2180.460 1111.720 2180.720 ;
      LAYER met2 ;
        RECT 17.570 2182.955 17.850 2183.325 ;
        RECT 17.640 2180.750 17.780 2182.955 ;
        RECT 17.580 2180.430 17.840 2180.750 ;
        RECT 1111.460 2180.430 1111.720 2180.750 ;
        RECT 1111.520 852.565 1111.660 2180.430 ;
        RECT 1111.450 852.195 1111.730 852.565 ;
      LAYER via2 ;
        RECT 17.570 2183.000 17.850 2183.280 ;
        RECT 1111.450 852.240 1111.730 852.520 ;
      LAYER met3 ;
        RECT -4.800 2183.290 2.400 2183.740 ;
        RECT 17.545 2183.290 17.875 2183.305 ;
        RECT -4.800 2182.990 17.875 2183.290 ;
        RECT -4.800 2182.540 2.400 2182.990 ;
        RECT 17.545 2182.975 17.875 2182.990 ;
        RECT 1111.425 852.530 1111.755 852.545 ;
        RECT 1098.790 852.230 1111.755 852.530 ;
        RECT 1098.790 850.120 1099.090 852.230 ;
        RECT 1111.425 852.215 1111.755 852.230 ;
        RECT 1096.000 849.520 1100.000 850.120 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 959.040 17.410 959.100 ;
        RECT 190.050 959.040 190.370 959.100 ;
        RECT 17.090 958.900 190.370 959.040 ;
        RECT 17.090 958.840 17.410 958.900 ;
        RECT 190.050 958.840 190.370 958.900 ;
      LAYER via ;
        RECT 17.120 958.840 17.380 959.100 ;
        RECT 190.080 958.840 190.340 959.100 ;
      LAYER met2 ;
        RECT 17.110 1921.835 17.390 1922.205 ;
        RECT 17.180 959.130 17.320 1921.835 ;
        RECT 17.120 958.810 17.380 959.130 ;
        RECT 190.080 958.810 190.340 959.130 ;
        RECT 190.140 958.645 190.280 958.810 ;
        RECT 190.070 958.275 190.350 958.645 ;
      LAYER via2 ;
        RECT 17.110 1921.880 17.390 1922.160 ;
        RECT 190.070 958.320 190.350 958.600 ;
      LAYER met3 ;
        RECT -4.800 1922.170 2.400 1922.620 ;
        RECT 17.085 1922.170 17.415 1922.185 ;
        RECT -4.800 1921.870 17.415 1922.170 ;
        RECT -4.800 1921.420 2.400 1921.870 ;
        RECT 17.085 1921.855 17.415 1921.870 ;
        RECT 190.045 958.610 190.375 958.625 ;
        RECT 190.045 958.310 202.090 958.610 ;
        RECT 190.045 958.295 190.375 958.310 ;
        RECT 201.790 957.560 202.090 958.310 ;
        RECT 200.000 956.960 204.000 957.560 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1656.380 16.490 1656.440 ;
        RECT 927.890 1656.380 928.210 1656.440 ;
        RECT 16.170 1656.240 928.210 1656.380 ;
        RECT 16.170 1656.180 16.490 1656.240 ;
        RECT 927.890 1656.180 928.210 1656.240 ;
        RECT 927.890 1012.080 928.210 1012.140 ;
        RECT 1080.150 1012.080 1080.470 1012.140 ;
        RECT 927.890 1011.940 1080.470 1012.080 ;
        RECT 927.890 1011.880 928.210 1011.940 ;
        RECT 1080.150 1011.880 1080.470 1011.940 ;
      LAYER via ;
        RECT 16.200 1656.180 16.460 1656.440 ;
        RECT 927.920 1656.180 928.180 1656.440 ;
        RECT 927.920 1011.880 928.180 1012.140 ;
        RECT 1080.180 1011.880 1080.440 1012.140 ;
      LAYER met2 ;
        RECT 16.190 1661.395 16.470 1661.765 ;
        RECT 16.260 1656.470 16.400 1661.395 ;
        RECT 16.200 1656.150 16.460 1656.470 ;
        RECT 927.920 1656.150 928.180 1656.470 ;
        RECT 927.980 1012.170 928.120 1656.150 ;
        RECT 927.920 1011.850 928.180 1012.170 ;
        RECT 1080.180 1011.850 1080.440 1012.170 ;
        RECT 1080.240 999.330 1080.380 1011.850 ;
        RECT 1081.910 999.330 1082.190 1000.000 ;
        RECT 1080.240 999.190 1082.190 999.330 ;
        RECT 1081.910 996.000 1082.190 999.190 ;
      LAYER via2 ;
        RECT 16.190 1661.440 16.470 1661.720 ;
      LAYER met3 ;
        RECT -4.800 1661.730 2.400 1662.180 ;
        RECT 16.165 1661.730 16.495 1661.745 ;
        RECT -4.800 1661.430 16.495 1661.730 ;
        RECT -4.800 1660.980 2.400 1661.430 ;
        RECT 16.165 1661.415 16.495 1661.430 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1393.900 16.490 1393.960 ;
        RECT 934.790 1393.900 935.110 1393.960 ;
        RECT 16.170 1393.760 935.110 1393.900 ;
        RECT 16.170 1393.700 16.490 1393.760 ;
        RECT 934.790 1393.700 935.110 1393.760 ;
        RECT 934.790 1012.420 935.110 1012.480 ;
        RECT 1087.510 1012.420 1087.830 1012.480 ;
        RECT 934.790 1012.280 1087.830 1012.420 ;
        RECT 934.790 1012.220 935.110 1012.280 ;
        RECT 1087.510 1012.220 1087.830 1012.280 ;
      LAYER via ;
        RECT 16.200 1393.700 16.460 1393.960 ;
        RECT 934.820 1393.700 935.080 1393.960 ;
        RECT 934.820 1012.220 935.080 1012.480 ;
        RECT 1087.540 1012.220 1087.800 1012.480 ;
      LAYER met2 ;
        RECT 16.190 1400.275 16.470 1400.645 ;
        RECT 16.260 1393.990 16.400 1400.275 ;
        RECT 16.200 1393.670 16.460 1393.990 ;
        RECT 934.820 1393.670 935.080 1393.990 ;
        RECT 934.880 1012.510 935.020 1393.670 ;
        RECT 934.820 1012.190 935.080 1012.510 ;
        RECT 1087.540 1012.190 1087.800 1012.510 ;
        RECT 1087.600 999.330 1087.740 1012.190 ;
        RECT 1089.270 999.330 1089.550 1000.000 ;
        RECT 1087.600 999.190 1089.550 999.330 ;
        RECT 1089.270 996.000 1089.550 999.190 ;
      LAYER via2 ;
        RECT 16.190 1400.320 16.470 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.165 1400.610 16.495 1400.625 ;
        RECT -4.800 1400.310 16.495 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.165 1400.295 16.495 1400.310 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1138.900 17.870 1138.960 ;
        RECT 941.690 1138.900 942.010 1138.960 ;
        RECT 17.550 1138.760 942.010 1138.900 ;
        RECT 17.550 1138.700 17.870 1138.760 ;
        RECT 941.690 1138.700 942.010 1138.760 ;
        RECT 941.690 1012.760 942.010 1012.820 ;
        RECT 1094.870 1012.760 1095.190 1012.820 ;
        RECT 941.690 1012.620 1095.190 1012.760 ;
        RECT 941.690 1012.560 942.010 1012.620 ;
        RECT 1094.870 1012.560 1095.190 1012.620 ;
      LAYER via ;
        RECT 17.580 1138.700 17.840 1138.960 ;
        RECT 941.720 1138.700 941.980 1138.960 ;
        RECT 941.720 1012.560 941.980 1012.820 ;
        RECT 1094.900 1012.560 1095.160 1012.820 ;
      LAYER met2 ;
        RECT 17.570 1139.835 17.850 1140.205 ;
        RECT 17.640 1138.990 17.780 1139.835 ;
        RECT 17.580 1138.670 17.840 1138.990 ;
        RECT 941.720 1138.670 941.980 1138.990 ;
        RECT 941.780 1012.850 941.920 1138.670 ;
        RECT 941.720 1012.530 941.980 1012.850 ;
        RECT 1094.900 1012.530 1095.160 1012.850 ;
        RECT 1094.960 999.330 1095.100 1012.530 ;
        RECT 1096.170 999.330 1096.450 1000.000 ;
        RECT 1094.960 999.190 1096.450 999.330 ;
        RECT 1096.170 996.000 1096.450 999.190 ;
      LAYER via2 ;
        RECT 17.570 1139.880 17.850 1140.160 ;
      LAYER met3 ;
        RECT -4.800 1140.170 2.400 1140.620 ;
        RECT 17.545 1140.170 17.875 1140.185 ;
        RECT -4.800 1139.870 17.875 1140.170 ;
        RECT -4.800 1139.420 2.400 1139.870 ;
        RECT 17.545 1139.855 17.875 1139.870 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 199.710 998.140 200.030 998.200 ;
        RECT 272.390 998.140 272.710 998.200 ;
        RECT 199.710 998.000 272.710 998.140 ;
        RECT 199.710 997.940 200.030 998.000 ;
        RECT 272.390 997.940 272.710 998.000 ;
        RECT 490.890 998.140 491.210 998.200 ;
        RECT 503.770 998.140 504.090 998.200 ;
        RECT 490.890 998.000 504.090 998.140 ;
        RECT 490.890 997.940 491.210 998.000 ;
        RECT 503.770 997.940 504.090 998.000 ;
        RECT 272.390 997.260 272.710 997.520 ;
        RECT 490.890 997.260 491.210 997.520 ;
        RECT 503.770 997.260 504.090 997.520 ;
        RECT 272.480 996.780 272.620 997.260 ;
        RECT 490.980 996.780 491.120 997.260 ;
        RECT 272.480 996.640 296.770 996.780 ;
        RECT 199.710 996.100 200.030 996.160 ;
        RECT 131.030 995.960 200.030 996.100 ;
        RECT 15.710 995.080 16.030 995.140 ;
        RECT 131.030 995.080 131.170 995.960 ;
        RECT 199.710 995.900 200.030 995.960 ;
        RECT 15.710 994.940 131.170 995.080 ;
        RECT 296.630 995.080 296.770 996.640 ;
        RECT 427.730 996.640 469.270 996.780 ;
        RECT 427.730 995.080 427.870 996.640 ;
        RECT 469.130 996.440 469.270 996.640 ;
        RECT 469.820 996.640 491.120 996.780 ;
        RECT 469.820 996.440 469.960 996.640 ;
        RECT 469.130 996.300 469.960 996.440 ;
        RECT 503.860 996.440 504.000 997.260 ;
        RECT 503.860 996.300 517.570 996.440 ;
        RECT 296.630 994.940 427.870 995.080 ;
        RECT 15.710 994.880 16.030 994.940 ;
        RECT 517.430 994.740 517.570 996.300 ;
        RECT 738.230 996.300 745.270 996.440 ;
        RECT 738.230 995.760 738.370 996.300 ;
        RECT 745.130 996.100 745.270 996.300 ;
        RECT 752.030 996.300 759.070 996.440 ;
        RECT 752.030 996.100 752.170 996.300 ;
        RECT 745.130 995.960 752.170 996.100 ;
        RECT 717.530 995.620 724.570 995.760 ;
        RECT 586.430 994.940 587.260 995.080 ;
        RECT 586.430 994.740 586.570 994.940 ;
        RECT 517.430 994.600 586.570 994.740 ;
        RECT 587.120 994.740 587.260 994.940 ;
        RECT 655.430 994.940 656.260 995.080 ;
        RECT 655.430 994.740 655.570 994.940 ;
        RECT 587.120 994.600 655.570 994.740 ;
        RECT 656.120 994.740 656.260 994.940 ;
        RECT 717.530 994.740 717.670 995.620 ;
        RECT 724.430 995.420 724.570 995.620 ;
        RECT 731.330 995.620 738.370 995.760 ;
        RECT 731.330 995.420 731.470 995.620 ;
        RECT 724.430 995.280 731.470 995.420 ;
        RECT 758.930 995.420 759.070 996.300 ;
        RECT 841.730 996.300 848.770 996.440 ;
        RECT 793.430 995.620 800.470 995.760 ;
        RECT 758.930 995.280 765.970 995.420 ;
        RECT 765.830 995.080 765.970 995.280 ;
        RECT 772.730 995.280 786.670 995.420 ;
        RECT 772.730 995.080 772.870 995.280 ;
        RECT 765.830 994.940 772.870 995.080 ;
        RECT 786.530 995.080 786.670 995.280 ;
        RECT 793.430 995.080 793.570 995.620 ;
        RECT 800.330 995.420 800.470 995.620 ;
        RECT 814.130 995.620 821.170 995.760 ;
        RECT 800.330 995.280 807.370 995.420 ;
        RECT 786.530 994.940 793.570 995.080 ;
        RECT 807.230 995.080 807.370 995.280 ;
        RECT 814.130 995.080 814.270 995.620 ;
        RECT 821.030 995.420 821.170 995.620 ;
        RECT 841.730 995.420 841.870 996.300 ;
        RECT 848.630 995.760 848.770 996.300 ;
        RECT 848.630 995.620 862.570 995.760 ;
        RECT 821.030 995.280 841.870 995.420 ;
        RECT 807.230 994.940 814.270 995.080 ;
        RECT 656.120 994.600 717.670 994.740 ;
        RECT 862.430 994.740 862.570 995.620 ;
        RECT 1112.350 995.080 1112.670 995.140 ;
        RECT 869.330 994.940 889.020 995.080 ;
        RECT 869.330 994.740 869.470 994.940 ;
        RECT 862.430 994.600 869.470 994.740 ;
        RECT 888.880 994.740 889.020 994.940 ;
        RECT 917.630 994.940 1112.670 995.080 ;
        RECT 917.630 994.740 917.770 994.940 ;
        RECT 1112.350 994.880 1112.670 994.940 ;
        RECT 888.880 994.600 917.770 994.740 ;
      LAYER via ;
        RECT 199.740 997.940 200.000 998.200 ;
        RECT 272.420 997.940 272.680 998.200 ;
        RECT 490.920 997.940 491.180 998.200 ;
        RECT 503.800 997.940 504.060 998.200 ;
        RECT 272.420 997.260 272.680 997.520 ;
        RECT 490.920 997.260 491.180 997.520 ;
        RECT 503.800 997.260 504.060 997.520 ;
        RECT 15.740 994.880 16.000 995.140 ;
        RECT 199.740 995.900 200.000 996.160 ;
        RECT 1112.380 994.880 1112.640 995.140 ;
      LAYER met2 ;
        RECT 199.740 997.910 200.000 998.230 ;
        RECT 272.420 997.910 272.680 998.230 ;
        RECT 490.920 997.910 491.180 998.230 ;
        RECT 503.800 997.910 504.060 998.230 ;
        RECT 199.800 996.190 199.940 997.910 ;
        RECT 272.480 997.550 272.620 997.910 ;
        RECT 490.980 997.550 491.120 997.910 ;
        RECT 503.860 997.550 504.000 997.910 ;
        RECT 272.420 997.230 272.680 997.550 ;
        RECT 490.920 997.230 491.180 997.550 ;
        RECT 503.800 997.230 504.060 997.550 ;
        RECT 199.740 995.870 200.000 996.190 ;
        RECT 15.740 994.850 16.000 995.170 ;
        RECT 1112.380 994.850 1112.640 995.170 ;
        RECT 15.800 879.765 15.940 994.850 ;
        RECT 1112.440 909.005 1112.580 994.850 ;
        RECT 1112.370 908.635 1112.650 909.005 ;
        RECT 15.730 879.395 16.010 879.765 ;
      LAYER via2 ;
        RECT 1112.370 908.680 1112.650 908.960 ;
        RECT 15.730 879.440 16.010 879.720 ;
      LAYER met3 ;
        RECT 1096.000 909.360 1100.000 909.960 ;
        RECT 1098.790 908.970 1099.090 909.360 ;
        RECT 1112.345 908.970 1112.675 908.985 ;
        RECT 1098.790 908.670 1112.675 908.970 ;
        RECT 1112.345 908.655 1112.675 908.670 ;
        RECT -4.800 879.730 2.400 880.180 ;
        RECT 15.705 879.730 16.035 879.745 ;
        RECT -4.800 879.430 16.035 879.730 ;
        RECT -4.800 878.980 2.400 879.430 ;
        RECT 15.705 879.415 16.035 879.430 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 989.555 20.610 989.925 ;
        RECT 1097.190 989.555 1097.470 989.925 ;
        RECT 20.400 618.645 20.540 989.555 ;
        RECT 1097.260 972.245 1097.400 989.555 ;
        RECT 1097.190 971.875 1097.470 972.245 ;
        RECT 20.330 618.275 20.610 618.645 ;
      LAYER via2 ;
        RECT 20.330 989.600 20.610 989.880 ;
        RECT 1097.190 989.600 1097.470 989.880 ;
        RECT 1097.190 971.920 1097.470 972.200 ;
        RECT 20.330 618.320 20.610 618.600 ;
      LAYER met3 ;
        RECT 20.305 989.890 20.635 989.905 ;
        RECT 1097.165 989.890 1097.495 989.905 ;
        RECT 20.305 989.590 1097.495 989.890 ;
        RECT 20.305 989.575 20.635 989.590 ;
        RECT 1097.165 989.575 1097.495 989.590 ;
        RECT 1097.165 972.210 1097.495 972.225 ;
        RECT 1096.950 971.895 1097.495 972.210 ;
        RECT 1096.950 969.800 1097.250 971.895 ;
        RECT 1096.000 969.200 1100.000 969.800 ;
        RECT -4.800 618.610 2.400 619.060 ;
        RECT 20.305 618.610 20.635 618.625 ;
        RECT -4.800 618.310 20.635 618.610 ;
        RECT -4.800 617.860 2.400 618.310 ;
        RECT 20.305 618.295 20.635 618.310 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.650 989.980 1114.970 990.040 ;
        RECT 2902.210 989.980 2902.530 990.040 ;
        RECT 1114.650 989.840 2902.530 989.980 ;
        RECT 1114.650 989.780 1114.970 989.840 ;
        RECT 2902.210 989.780 2902.530 989.840 ;
      LAYER via ;
        RECT 1114.680 989.780 1114.940 990.040 ;
        RECT 2902.240 989.780 2902.500 990.040 ;
      LAYER met2 ;
        RECT 2902.230 1958.555 2902.510 1958.925 ;
        RECT 2902.300 990.070 2902.440 1958.555 ;
        RECT 1114.680 989.750 1114.940 990.070 ;
        RECT 2902.240 989.750 2902.500 990.070 ;
        RECT 1114.740 611.845 1114.880 989.750 ;
        RECT 1114.670 611.475 1114.950 611.845 ;
      LAYER via2 ;
        RECT 2902.230 1958.600 2902.510 1958.880 ;
        RECT 1114.670 611.520 1114.950 611.800 ;
      LAYER met3 ;
        RECT 2902.205 1958.890 2902.535 1958.905 ;
        RECT 2917.600 1958.890 2924.800 1959.340 ;
        RECT 2902.205 1958.590 2924.800 1958.890 ;
        RECT 2902.205 1958.575 2902.535 1958.590 ;
        RECT 2917.600 1958.140 2924.800 1958.590 ;
        RECT 1114.645 611.810 1114.975 611.825 ;
        RECT 1098.790 611.510 1114.975 611.810 ;
        RECT 1098.790 610.080 1099.090 611.510 ;
        RECT 1114.645 611.495 1114.975 611.510 ;
        RECT 1096.000 609.480 1100.000 610.080 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.270 2222.140 1021.590 2222.200 ;
        RECT 2900.830 2222.140 2901.150 2222.200 ;
        RECT 1021.270 2222.000 2901.150 2222.140 ;
        RECT 1021.270 2221.940 1021.590 2222.000 ;
        RECT 2900.830 2221.940 2901.150 2222.000 ;
      LAYER via ;
        RECT 1021.300 2221.940 1021.560 2222.200 ;
        RECT 2900.860 2221.940 2901.120 2222.200 ;
      LAYER met2 ;
        RECT 2900.850 2223.755 2901.130 2224.125 ;
        RECT 2900.920 2222.230 2901.060 2223.755 ;
        RECT 1021.300 2221.910 1021.560 2222.230 ;
        RECT 2900.860 2221.910 2901.120 2222.230 ;
        RECT 1021.360 1048.870 1021.500 2221.910 ;
        RECT 1021.360 1048.730 1023.800 1048.870 ;
        RECT 1023.660 999.330 1023.800 1048.730 ;
        RECT 1025.330 999.330 1025.610 1000.000 ;
        RECT 1023.660 999.190 1025.610 999.330 ;
        RECT 1025.330 996.000 1025.610 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2223.800 2901.130 2224.080 ;
      LAYER met3 ;
        RECT 2900.825 2224.090 2901.155 2224.105 ;
        RECT 2917.600 2224.090 2924.800 2224.540 ;
        RECT 2900.825 2223.790 2924.800 2224.090 ;
        RECT 2900.825 2223.775 2901.155 2223.790 ;
        RECT 2917.600 2223.340 2924.800 2223.790 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 676.160 1117.730 676.220 ;
        RECT 2901.750 676.160 2902.070 676.220 ;
        RECT 1117.410 676.020 2902.070 676.160 ;
        RECT 1117.410 675.960 1117.730 676.020 ;
        RECT 2901.750 675.960 2902.070 676.020 ;
      LAYER via ;
        RECT 1117.440 675.960 1117.700 676.220 ;
        RECT 2901.780 675.960 2902.040 676.220 ;
      LAYER met2 ;
        RECT 2901.770 2489.635 2902.050 2490.005 ;
        RECT 2901.840 676.250 2901.980 2489.635 ;
        RECT 1117.440 675.930 1117.700 676.250 ;
        RECT 2901.780 675.930 2902.040 676.250 ;
        RECT 1117.500 672.365 1117.640 675.930 ;
        RECT 1117.430 671.995 1117.710 672.365 ;
      LAYER via2 ;
        RECT 2901.770 2489.680 2902.050 2489.960 ;
        RECT 1117.430 672.040 1117.710 672.320 ;
      LAYER met3 ;
        RECT 2901.745 2489.970 2902.075 2489.985 ;
        RECT 2917.600 2489.970 2924.800 2490.420 ;
        RECT 2901.745 2489.670 2924.800 2489.970 ;
        RECT 2901.745 2489.655 2902.075 2489.670 ;
        RECT 2917.600 2489.220 2924.800 2489.670 ;
        RECT 1117.405 672.330 1117.735 672.345 ;
        RECT 1098.790 672.030 1117.735 672.330 ;
        RECT 1098.790 669.920 1099.090 672.030 ;
        RECT 1117.405 672.015 1117.735 672.030 ;
        RECT 1096.000 669.320 1100.000 669.920 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.170 2753.220 1028.490 2753.280 ;
        RECT 2898.990 2753.220 2899.310 2753.280 ;
        RECT 1028.170 2753.080 2899.310 2753.220 ;
        RECT 1028.170 2753.020 1028.490 2753.080 ;
        RECT 2898.990 2753.020 2899.310 2753.080 ;
      LAYER via ;
        RECT 1028.200 2753.020 1028.460 2753.280 ;
        RECT 2899.020 2753.020 2899.280 2753.280 ;
      LAYER met2 ;
        RECT 2899.010 2755.515 2899.290 2755.885 ;
        RECT 2899.080 2753.310 2899.220 2755.515 ;
        RECT 1028.200 2752.990 1028.460 2753.310 ;
        RECT 2899.020 2752.990 2899.280 2753.310 ;
        RECT 1028.260 1048.870 1028.400 2752.990 ;
        RECT 1028.260 1048.730 1030.240 1048.870 ;
        RECT 1030.100 999.330 1030.240 1048.730 ;
        RECT 1032.230 999.330 1032.510 1000.000 ;
        RECT 1030.100 999.190 1032.510 999.330 ;
        RECT 1032.230 996.000 1032.510 999.190 ;
      LAYER via2 ;
        RECT 2899.010 2755.560 2899.290 2755.840 ;
      LAYER met3 ;
        RECT 2898.985 2755.850 2899.315 2755.865 ;
        RECT 2917.600 2755.850 2924.800 2756.300 ;
        RECT 2898.985 2755.550 2924.800 2755.850 ;
        RECT 2898.985 2755.535 2899.315 2755.550 ;
        RECT 2917.600 2755.100 2924.800 2755.550 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 191.890 3015.700 192.210 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 191.890 3015.560 2901.150 3015.700 ;
        RECT 191.890 3015.500 192.210 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 191.920 3015.500 192.180 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 191.920 3015.470 192.180 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 191.980 617.285 192.120 3015.470 ;
        RECT 191.910 616.915 192.190 617.285 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 191.910 616.960 192.190 617.240 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 191.885 617.250 192.215 617.265 ;
        RECT 191.885 616.950 201.170 617.250 ;
        RECT 191.885 616.935 192.215 616.950 ;
        RECT 200.870 614.840 201.170 616.950 ;
        RECT 200.000 614.240 204.000 614.840 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1093.490 393.280 1093.810 393.340 ;
        RECT 2901.290 393.280 2901.610 393.340 ;
        RECT 1093.490 393.140 2901.610 393.280 ;
        RECT 1093.490 393.080 1093.810 393.140 ;
        RECT 2901.290 393.080 2901.610 393.140 ;
      LAYER via ;
        RECT 1093.520 393.080 1093.780 393.340 ;
        RECT 2901.320 393.080 2901.580 393.340 ;
      LAYER met2 ;
        RECT 2901.310 3286.595 2901.590 3286.965 ;
        RECT 1093.410 400.180 1093.690 404.000 ;
        RECT 1093.410 400.000 1093.720 400.180 ;
        RECT 1093.580 393.370 1093.720 400.000 ;
        RECT 2901.380 393.370 2901.520 3286.595 ;
        RECT 1093.520 393.050 1093.780 393.370 ;
        RECT 2901.320 393.050 2901.580 393.370 ;
      LAYER via2 ;
        RECT 2901.310 3286.640 2901.590 3286.920 ;
      LAYER met3 ;
        RECT 2901.285 3286.930 2901.615 3286.945 ;
        RECT 2917.600 3286.930 2924.800 3287.380 ;
        RECT 2901.285 3286.630 2924.800 3286.930 ;
        RECT 2901.285 3286.615 2901.615 3286.630 ;
        RECT 2917.600 3286.180 2924.800 3286.630 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
        RECT 2879.300 3512.170 2879.440 3517.600 ;
        RECT 2877.460 3512.030 2879.440 3512.170 ;
        RECT 2877.460 1011.005 2877.600 3512.030 ;
        RECT 1041.070 1010.635 1041.350 1011.005 ;
        RECT 2877.390 1010.635 2877.670 1011.005 ;
        RECT 1039.590 999.330 1039.870 1000.000 ;
        RECT 1041.140 999.330 1041.280 1010.635 ;
        RECT 1039.590 999.190 1041.280 999.330 ;
        RECT 1039.590 996.000 1039.870 999.190 ;
      LAYER via2 ;
        RECT 1041.070 1010.680 1041.350 1010.960 ;
        RECT 2877.390 1010.680 2877.670 1010.960 ;
      LAYER met3 ;
        RECT 1041.045 1010.970 1041.375 1010.985 ;
        RECT 2877.365 1010.970 2877.695 1010.985 ;
        RECT 1041.045 1010.670 2877.695 1010.970 ;
        RECT 1041.045 1010.655 1041.375 1010.670 ;
        RECT 2877.365 1010.655 2877.695 1010.670 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1095.330 392.940 1095.650 393.000 ;
        RECT 2553.070 392.940 2553.390 393.000 ;
        RECT 1095.330 392.800 2553.390 392.940 ;
        RECT 1095.330 392.740 1095.650 392.800 ;
        RECT 2553.070 392.740 2553.390 392.800 ;
      LAYER via ;
        RECT 1095.360 392.740 1095.620 393.000 ;
        RECT 2553.100 392.740 2553.360 393.000 ;
      LAYER met2 ;
        RECT 2553.160 3517.910 2554.220 3518.050 ;
        RECT 1095.250 400.180 1095.530 404.000 ;
        RECT 1095.250 400.000 1095.560 400.180 ;
        RECT 1095.420 393.030 1095.560 400.000 ;
        RECT 2553.160 393.030 2553.300 3517.910 ;
        RECT 2554.080 3517.370 2554.220 3517.910 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
        RECT 2555.000 3517.370 2555.140 3517.600 ;
        RECT 2554.080 3517.230 2555.140 3517.370 ;
        RECT 1095.360 392.710 1095.620 393.030 ;
        RECT 2553.100 392.710 2553.360 393.030 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.170 99.860 200.490 99.920 ;
        RECT 2901.290 99.860 2901.610 99.920 ;
        RECT 200.170 99.720 2901.610 99.860 ;
        RECT 200.170 99.660 200.490 99.720 ;
        RECT 2901.290 99.660 2901.610 99.720 ;
      LAYER via ;
        RECT 200.200 99.660 200.460 99.920 ;
        RECT 2901.320 99.660 2901.580 99.920 ;
      LAYER met2 ;
        RECT 203.310 996.610 203.590 1000.000 ;
        RECT 200.260 996.470 203.590 996.610 ;
        RECT 200.260 99.950 200.400 996.470 ;
        RECT 203.310 996.000 203.590 996.470 ;
        RECT 200.200 99.630 200.460 99.950 ;
        RECT 2901.320 99.630 2901.580 99.950 ;
        RECT 2901.380 33.165 2901.520 99.630 ;
        RECT 2901.310 32.795 2901.590 33.165 ;
      LAYER via2 ;
        RECT 2901.310 32.840 2901.590 33.120 ;
      LAYER met3 ;
        RECT 2901.285 33.130 2901.615 33.145 ;
        RECT 2917.600 33.130 2924.800 33.580 ;
        RECT 2901.285 32.830 2924.800 33.130 ;
        RECT 2901.285 32.815 2901.615 32.830 ;
        RECT 2917.600 32.380 2924.800 32.830 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 2284.020 414.390 2284.080 ;
        RECT 2900.830 2284.020 2901.150 2284.080 ;
        RECT 414.070 2283.880 2901.150 2284.020 ;
        RECT 414.070 2283.820 414.390 2283.880 ;
        RECT 2900.830 2283.820 2901.150 2283.880 ;
      LAYER via ;
        RECT 414.100 2283.820 414.360 2284.080 ;
        RECT 2900.860 2283.820 2901.120 2284.080 ;
      LAYER met2 ;
        RECT 2900.850 2290.395 2901.130 2290.765 ;
        RECT 2900.920 2284.110 2901.060 2290.395 ;
        RECT 414.100 2283.790 414.360 2284.110 ;
        RECT 2900.860 2283.790 2901.120 2284.110 ;
        RECT 414.160 999.330 414.300 2283.790 ;
        RECT 415.830 999.330 416.110 1000.000 ;
        RECT 414.160 999.190 416.110 999.330 ;
        RECT 415.830 996.000 416.110 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2290.440 2901.130 2290.720 ;
      LAYER met3 ;
        RECT 2900.825 2290.730 2901.155 2290.745 ;
        RECT 2917.600 2290.730 2924.800 2291.180 ;
        RECT 2900.825 2290.430 2924.800 2290.730 ;
        RECT 2900.825 2290.415 2901.155 2290.430 ;
        RECT 2917.600 2289.980 2924.800 2290.430 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 2553.300 435.090 2553.360 ;
        RECT 2900.830 2553.300 2901.150 2553.360 ;
        RECT 434.770 2553.160 2901.150 2553.300 ;
        RECT 434.770 2553.100 435.090 2553.160 ;
        RECT 2900.830 2553.100 2901.150 2553.160 ;
      LAYER via ;
        RECT 434.800 2553.100 435.060 2553.360 ;
        RECT 2900.860 2553.100 2901.120 2553.360 ;
      LAYER met2 ;
        RECT 2900.850 2556.275 2901.130 2556.645 ;
        RECT 2900.920 2553.390 2901.060 2556.275 ;
        RECT 434.800 2553.070 435.060 2553.390 ;
        RECT 2900.860 2553.070 2901.120 2553.390 ;
        RECT 434.860 999.330 435.000 2553.070 ;
        RECT 436.990 999.330 437.270 1000.000 ;
        RECT 434.860 999.190 437.270 999.330 ;
        RECT 436.990 996.000 437.270 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2556.320 2901.130 2556.600 ;
      LAYER met3 ;
        RECT 2900.825 2556.610 2901.155 2556.625 ;
        RECT 2917.600 2556.610 2924.800 2557.060 ;
        RECT 2900.825 2556.310 2924.800 2556.610 ;
        RECT 2900.825 2556.295 2901.155 2556.310 ;
        RECT 2917.600 2555.860 2924.800 2556.310 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 2815.440 455.790 2815.500 ;
        RECT 2900.830 2815.440 2901.150 2815.500 ;
        RECT 455.470 2815.300 2901.150 2815.440 ;
        RECT 455.470 2815.240 455.790 2815.300 ;
        RECT 2900.830 2815.240 2901.150 2815.300 ;
      LAYER via ;
        RECT 455.500 2815.240 455.760 2815.500 ;
        RECT 2900.860 2815.240 2901.120 2815.500 ;
      LAYER met2 ;
        RECT 2900.850 2821.475 2901.130 2821.845 ;
        RECT 2900.920 2815.530 2901.060 2821.475 ;
        RECT 455.500 2815.210 455.760 2815.530 ;
        RECT 2900.860 2815.210 2901.120 2815.530 ;
        RECT 455.560 1048.870 455.700 2815.210 ;
        RECT 455.560 1048.730 456.160 1048.870 ;
        RECT 456.020 999.330 456.160 1048.730 ;
        RECT 458.150 999.330 458.430 1000.000 ;
        RECT 456.020 999.190 458.430 999.330 ;
        RECT 458.150 996.000 458.430 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2821.520 2901.130 2821.800 ;
      LAYER met3 ;
        RECT 2900.825 2821.810 2901.155 2821.825 ;
        RECT 2917.600 2821.810 2924.800 2822.260 ;
        RECT 2900.825 2821.510 2924.800 2821.810 ;
        RECT 2900.825 2821.495 2901.155 2821.510 ;
        RECT 2917.600 2821.060 2924.800 2821.510 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 3084.380 476.490 3084.440 ;
        RECT 2900.830 3084.380 2901.150 3084.440 ;
        RECT 476.170 3084.240 2901.150 3084.380 ;
        RECT 476.170 3084.180 476.490 3084.240 ;
        RECT 2900.830 3084.180 2901.150 3084.240 ;
      LAYER via ;
        RECT 476.200 3084.180 476.460 3084.440 ;
        RECT 2900.860 3084.180 2901.120 3084.440 ;
      LAYER met2 ;
        RECT 2900.850 3087.355 2901.130 3087.725 ;
        RECT 2900.920 3084.470 2901.060 3087.355 ;
        RECT 476.200 3084.150 476.460 3084.470 ;
        RECT 2900.860 3084.150 2901.120 3084.470 ;
        RECT 476.260 1048.870 476.400 3084.150 ;
        RECT 476.260 1048.730 477.320 1048.870 ;
        RECT 477.180 999.330 477.320 1048.730 ;
        RECT 479.310 999.330 479.590 1000.000 ;
        RECT 477.180 999.190 479.590 999.330 ;
        RECT 479.310 996.000 479.590 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3087.400 2901.130 3087.680 ;
      LAYER met3 ;
        RECT 2900.825 3087.690 2901.155 3087.705 ;
        RECT 2917.600 3087.690 2924.800 3088.140 ;
        RECT 2900.825 3087.390 2924.800 3087.690 ;
        RECT 2900.825 3087.375 2901.155 3087.390 ;
        RECT 2917.600 3086.940 2924.800 3087.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 3353.660 497.190 3353.720 ;
        RECT 2900.830 3353.660 2901.150 3353.720 ;
        RECT 496.870 3353.520 2901.150 3353.660 ;
        RECT 496.870 3353.460 497.190 3353.520 ;
        RECT 2900.830 3353.460 2901.150 3353.520 ;
      LAYER via ;
        RECT 496.900 3353.460 497.160 3353.720 ;
        RECT 2900.860 3353.460 2901.120 3353.720 ;
      LAYER met2 ;
        RECT 496.900 3353.430 497.160 3353.750 ;
        RECT 2900.860 3353.605 2901.120 3353.750 ;
        RECT 496.960 1048.870 497.100 3353.430 ;
        RECT 2900.850 3353.235 2901.130 3353.605 ;
        RECT 496.960 1048.730 499.400 1048.870 ;
        RECT 499.260 999.330 499.400 1048.730 ;
        RECT 500.930 999.330 501.210 1000.000 ;
        RECT 499.260 999.190 501.210 999.330 ;
        RECT 500.930 996.000 501.210 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3353.280 2901.130 3353.560 ;
      LAYER met3 ;
        RECT 2900.825 3353.570 2901.155 3353.585 ;
        RECT 2917.600 3353.570 2924.800 3354.020 ;
        RECT 2900.825 3353.270 2924.800 3353.570 ;
        RECT 2900.825 3353.255 2901.155 3353.270 ;
        RECT 2917.600 3352.820 2924.800 3353.270 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.330 1017.860 520.650 1017.920 ;
        RECT 2794.570 1017.860 2794.890 1017.920 ;
        RECT 520.330 1017.720 2794.890 1017.860 ;
        RECT 520.330 1017.660 520.650 1017.720 ;
        RECT 2794.570 1017.660 2794.890 1017.720 ;
      LAYER via ;
        RECT 520.360 1017.660 520.620 1017.920 ;
        RECT 2794.600 1017.660 2794.860 1017.920 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3512.170 2798.480 3517.600 ;
        RECT 2794.660 3512.030 2798.480 3512.170 ;
        RECT 2794.660 1017.950 2794.800 3512.030 ;
        RECT 520.360 1017.630 520.620 1017.950 ;
        RECT 2794.600 1017.630 2794.860 1017.950 ;
        RECT 520.420 999.330 520.560 1017.630 ;
        RECT 522.090 999.330 522.370 1000.000 ;
        RECT 520.420 999.190 522.370 999.330 ;
        RECT 522.090 996.000 522.370 999.190 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.490 1018.200 541.810 1018.260 ;
        RECT 2470.270 1018.200 2470.590 1018.260 ;
        RECT 541.490 1018.060 2470.590 1018.200 ;
        RECT 541.490 1018.000 541.810 1018.060 ;
        RECT 2470.270 1018.000 2470.590 1018.060 ;
      LAYER via ;
        RECT 541.520 1018.000 541.780 1018.260 ;
        RECT 2470.300 1018.000 2470.560 1018.260 ;
      LAYER met2 ;
        RECT 2470.360 3517.910 2473.260 3518.050 ;
        RECT 2470.360 1018.290 2470.500 3517.910 ;
        RECT 2473.120 3517.370 2473.260 3517.910 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2473.120 3517.230 2474.180 3517.370 ;
        RECT 541.520 1017.970 541.780 1018.290 ;
        RECT 2470.300 1017.970 2470.560 1018.290 ;
        RECT 541.580 999.330 541.720 1017.970 ;
        RECT 543.250 999.330 543.530 1000.000 ;
        RECT 541.580 999.190 543.530 999.330 ;
        RECT 543.250 996.000 543.530 999.190 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 562.650 1018.540 562.970 1018.600 ;
        RECT 2145.970 1018.540 2146.290 1018.600 ;
        RECT 562.650 1018.400 2146.290 1018.540 ;
        RECT 562.650 1018.340 562.970 1018.400 ;
        RECT 2145.970 1018.340 2146.290 1018.400 ;
      LAYER via ;
        RECT 562.680 1018.340 562.940 1018.600 ;
        RECT 2146.000 1018.340 2146.260 1018.600 ;
      LAYER met2 ;
        RECT 2146.060 3517.910 2148.500 3518.050 ;
        RECT 2146.060 1018.630 2146.200 3517.910 ;
        RECT 2148.360 3517.370 2148.500 3517.910 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2148.360 3517.230 2149.420 3517.370 ;
        RECT 562.680 1018.310 562.940 1018.630 ;
        RECT 2146.000 1018.310 2146.260 1018.630 ;
        RECT 562.740 999.330 562.880 1018.310 ;
        RECT 564.410 999.330 564.690 1000.000 ;
        RECT 562.740 999.190 564.690 999.330 ;
        RECT 564.410 996.000 564.690 999.190 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 583.810 1018.880 584.130 1018.940 ;
        RECT 1821.670 1018.880 1821.990 1018.940 ;
        RECT 583.810 1018.740 1821.990 1018.880 ;
        RECT 583.810 1018.680 584.130 1018.740 ;
        RECT 1821.670 1018.680 1821.990 1018.740 ;
      LAYER via ;
        RECT 583.840 1018.680 584.100 1018.940 ;
        RECT 1821.700 1018.680 1821.960 1018.940 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3512.170 1825.120 3517.600 ;
        RECT 1821.760 3512.030 1825.120 3512.170 ;
        RECT 1821.760 1018.970 1821.900 3512.030 ;
        RECT 583.840 1018.650 584.100 1018.970 ;
        RECT 1821.700 1018.650 1821.960 1018.970 ;
        RECT 583.900 999.330 584.040 1018.650 ;
        RECT 586.030 999.330 586.310 1000.000 ;
        RECT 583.900 999.190 586.310 999.330 ;
        RECT 586.030 996.000 586.310 999.190 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1102.320 3505.500 1104.760 3505.640 ;
        RECT 1095.330 3504.960 1095.650 3505.020 ;
        RECT 1102.320 3504.960 1102.460 3505.500 ;
        RECT 1095.330 3504.820 1102.460 3504.960 ;
        RECT 1095.330 3504.760 1095.650 3504.820 ;
        RECT 1104.620 3504.620 1104.760 3505.500 ;
        RECT 1500.590 3504.620 1500.910 3504.680 ;
        RECT 1104.620 3504.480 1500.910 3504.620 ;
        RECT 1500.590 3504.420 1500.910 3504.480 ;
        RECT 1093.490 3498.500 1093.810 3498.560 ;
        RECT 1095.330 3498.500 1095.650 3498.560 ;
        RECT 1093.490 3498.360 1095.650 3498.500 ;
        RECT 1093.490 3498.300 1093.810 3498.360 ;
        RECT 1095.330 3498.300 1095.650 3498.360 ;
        RECT 607.730 1020.580 608.050 1020.640 ;
        RECT 1093.490 1020.580 1093.810 1020.640 ;
        RECT 607.730 1020.440 1093.810 1020.580 ;
        RECT 607.730 1020.380 608.050 1020.440 ;
        RECT 1093.490 1020.380 1093.810 1020.440 ;
      LAYER via ;
        RECT 1095.360 3504.760 1095.620 3505.020 ;
        RECT 1500.620 3504.420 1500.880 3504.680 ;
        RECT 1093.520 3498.300 1093.780 3498.560 ;
        RECT 1095.360 3498.300 1095.620 3498.560 ;
        RECT 607.760 1020.380 608.020 1020.640 ;
        RECT 1093.520 1020.380 1093.780 1020.640 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1095.360 3504.730 1095.620 3505.050 ;
        RECT 1095.420 3498.590 1095.560 3504.730 ;
        RECT 1500.680 3504.710 1500.820 3517.600 ;
        RECT 1500.620 3504.390 1500.880 3504.710 ;
        RECT 1093.520 3498.270 1093.780 3498.590 ;
        RECT 1095.360 3498.270 1095.620 3498.590 ;
        RECT 1093.580 1020.670 1093.720 3498.270 ;
        RECT 607.760 1020.350 608.020 1020.670 ;
        RECT 1093.520 1020.350 1093.780 1020.670 ;
        RECT 607.190 999.330 607.470 1000.000 ;
        RECT 607.820 999.330 607.960 1020.350 ;
        RECT 607.190 999.190 607.960 999.330 ;
        RECT 607.190 996.000 607.470 999.190 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 225.930 1001.200 226.250 1001.260 ;
        RECT 2903.590 1001.200 2903.910 1001.260 ;
        RECT 225.930 1001.060 2903.910 1001.200 ;
        RECT 225.930 1001.000 226.250 1001.060 ;
        RECT 2903.590 1001.000 2903.910 1001.060 ;
      LAYER via ;
        RECT 225.960 1001.000 226.220 1001.260 ;
        RECT 2903.620 1001.000 2903.880 1001.260 ;
      LAYER met2 ;
        RECT 225.960 1000.970 226.220 1001.290 ;
        RECT 2903.620 1000.970 2903.880 1001.290 ;
        RECT 224.470 999.330 224.750 1000.000 ;
        RECT 226.020 999.330 226.160 1000.970 ;
        RECT 224.470 999.190 226.160 999.330 ;
        RECT 224.470 996.000 224.750 999.190 ;
        RECT 2903.680 231.725 2903.820 1000.970 ;
        RECT 2903.610 231.355 2903.890 231.725 ;
      LAYER via2 ;
        RECT 2903.610 231.400 2903.890 231.680 ;
      LAYER met3 ;
        RECT 2903.585 231.690 2903.915 231.705 ;
        RECT 2917.600 231.690 2924.800 232.140 ;
        RECT 2903.585 231.390 2924.800 231.690 ;
        RECT 2903.585 231.375 2903.915 231.390 ;
        RECT 2917.600 230.940 2924.800 231.390 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1102.690 3504.760 1103.010 3505.020 ;
        RECT 1104.990 3504.960 1105.310 3505.020 ;
        RECT 1175.830 3504.960 1176.150 3505.020 ;
        RECT 1104.990 3504.820 1176.150 3504.960 ;
        RECT 1104.990 3504.760 1105.310 3504.820 ;
        RECT 1175.830 3504.760 1176.150 3504.820 ;
        RECT 1093.950 3504.620 1094.270 3504.680 ;
        RECT 1102.780 3504.620 1102.920 3504.760 ;
        RECT 1093.950 3504.480 1102.920 3504.620 ;
        RECT 1093.950 3504.420 1094.270 3504.480 ;
        RECT 627.970 1021.260 628.290 1021.320 ;
        RECT 1093.950 1021.260 1094.270 1021.320 ;
        RECT 627.970 1021.120 1094.270 1021.260 ;
        RECT 627.970 1021.060 628.290 1021.120 ;
        RECT 1093.950 1021.060 1094.270 1021.120 ;
      LAYER via ;
        RECT 1102.720 3504.760 1102.980 3505.020 ;
        RECT 1105.020 3504.760 1105.280 3505.020 ;
        RECT 1175.860 3504.760 1176.120 3505.020 ;
        RECT 1093.980 3504.420 1094.240 3504.680 ;
        RECT 628.000 1021.060 628.260 1021.320 ;
        RECT 1093.980 1021.060 1094.240 1021.320 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3505.050 1176.060 3517.600 ;
        RECT 1102.720 3504.960 1102.980 3505.050 ;
        RECT 1105.020 3504.960 1105.280 3505.050 ;
        RECT 1102.720 3504.820 1105.280 3504.960 ;
        RECT 1102.720 3504.730 1102.980 3504.820 ;
        RECT 1105.020 3504.730 1105.280 3504.820 ;
        RECT 1175.860 3504.730 1176.120 3505.050 ;
        RECT 1093.980 3504.390 1094.240 3504.710 ;
        RECT 1094.040 1021.350 1094.180 3504.390 ;
        RECT 628.000 1021.030 628.260 1021.350 ;
        RECT 1093.980 1021.030 1094.240 1021.350 ;
        RECT 628.060 999.330 628.200 1021.030 ;
        RECT 628.350 999.330 628.630 1000.000 ;
        RECT 628.060 999.190 628.630 999.330 ;
        RECT 628.350 996.000 628.630 999.190 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 1016.840 648.990 1016.900 ;
        RECT 848.770 1016.840 849.090 1016.900 ;
        RECT 648.670 1016.700 849.090 1016.840 ;
        RECT 648.670 1016.640 648.990 1016.700 ;
        RECT 848.770 1016.640 849.090 1016.700 ;
      LAYER via ;
        RECT 648.700 1016.640 648.960 1016.900 ;
        RECT 848.800 1016.640 849.060 1016.900 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3512.170 851.760 3517.600 ;
        RECT 848.860 3512.030 851.760 3512.170 ;
        RECT 848.860 1016.930 849.000 3512.030 ;
        RECT 648.700 1016.610 648.960 1016.930 ;
        RECT 848.800 1016.610 849.060 1016.930 ;
        RECT 648.760 999.330 648.900 1016.610 ;
        RECT 649.510 999.330 649.790 1000.000 ;
        RECT 648.760 999.190 649.790 999.330 ;
        RECT 649.510 996.000 649.790 999.190 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 1016.500 525.250 1016.560 ;
        RECT 669.370 1016.500 669.690 1016.560 ;
        RECT 524.930 1016.360 669.690 1016.500 ;
        RECT 524.930 1016.300 525.250 1016.360 ;
        RECT 669.370 1016.300 669.690 1016.360 ;
      LAYER via ;
        RECT 524.960 1016.300 525.220 1016.560 ;
        RECT 669.400 1016.300 669.660 1016.560 ;
      LAYER met2 ;
        RECT 525.020 3517.910 526.540 3518.050 ;
        RECT 525.020 1016.590 525.160 3517.910 ;
        RECT 526.400 3517.370 526.540 3517.910 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3517.370 527.460 3517.600 ;
        RECT 526.400 3517.230 527.460 3517.370 ;
        RECT 524.960 1016.270 525.220 1016.590 ;
        RECT 669.400 1016.270 669.660 1016.590 ;
        RECT 669.460 999.330 669.600 1016.270 ;
        RECT 671.130 999.330 671.410 1000.000 ;
        RECT 669.460 999.190 671.410 999.330 ;
        RECT 671.130 996.000 671.410 999.190 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.920 202.790 3502.980 ;
        RECT 224.090 3502.920 224.410 3502.980 ;
        RECT 202.470 3502.780 224.410 3502.920 ;
        RECT 202.470 3502.720 202.790 3502.780 ;
        RECT 224.090 3502.720 224.410 3502.780 ;
        RECT 224.090 1020.920 224.410 1020.980 ;
        RECT 690.530 1020.920 690.850 1020.980 ;
        RECT 224.090 1020.780 690.850 1020.920 ;
        RECT 224.090 1020.720 224.410 1020.780 ;
        RECT 690.530 1020.720 690.850 1020.780 ;
      LAYER via ;
        RECT 202.500 3502.720 202.760 3502.980 ;
        RECT 224.120 3502.720 224.380 3502.980 ;
        RECT 224.120 1020.720 224.380 1020.980 ;
        RECT 690.560 1020.720 690.820 1020.980 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3503.010 202.700 3517.600 ;
        RECT 202.500 3502.690 202.760 3503.010 ;
        RECT 224.120 3502.690 224.380 3503.010 ;
        RECT 224.180 1021.010 224.320 3502.690 ;
        RECT 224.120 1020.690 224.380 1021.010 ;
        RECT 690.560 1020.690 690.820 1021.010 ;
        RECT 690.620 999.330 690.760 1020.690 ;
        RECT 692.290 999.330 692.570 1000.000 ;
        RECT 690.620 999.190 692.570 999.330 ;
        RECT 692.290 996.000 692.570 999.190 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3415.880 17.410 3415.940 ;
        RECT 224.550 3415.880 224.870 3415.940 ;
        RECT 17.090 3415.740 224.870 3415.880 ;
        RECT 17.090 3415.680 17.410 3415.740 ;
        RECT 224.550 3415.680 224.870 3415.740 ;
        RECT 224.550 1020.240 224.870 1020.300 ;
        RECT 711.690 1020.240 712.010 1020.300 ;
        RECT 224.550 1020.100 712.010 1020.240 ;
        RECT 224.550 1020.040 224.870 1020.100 ;
        RECT 711.690 1020.040 712.010 1020.100 ;
      LAYER via ;
        RECT 17.120 3415.680 17.380 3415.940 ;
        RECT 224.580 3415.680 224.840 3415.940 ;
        RECT 224.580 1020.040 224.840 1020.300 ;
        RECT 711.720 1020.040 711.980 1020.300 ;
      LAYER met2 ;
        RECT 17.110 3421.235 17.390 3421.605 ;
        RECT 17.180 3415.970 17.320 3421.235 ;
        RECT 17.120 3415.650 17.380 3415.970 ;
        RECT 224.580 3415.650 224.840 3415.970 ;
        RECT 224.640 1020.330 224.780 3415.650 ;
        RECT 224.580 1020.010 224.840 1020.330 ;
        RECT 711.720 1020.010 711.980 1020.330 ;
        RECT 711.780 999.330 711.920 1020.010 ;
        RECT 713.450 999.330 713.730 1000.000 ;
        RECT 711.780 999.190 713.730 999.330 ;
        RECT 713.450 996.000 713.730 999.190 ;
      LAYER via2 ;
        RECT 17.110 3421.280 17.390 3421.560 ;
      LAYER met3 ;
        RECT -4.800 3421.570 2.400 3422.020 ;
        RECT 17.085 3421.570 17.415 3421.585 ;
        RECT -4.800 3421.270 17.415 3421.570 ;
        RECT -4.800 3420.820 2.400 3421.270 ;
        RECT 17.085 3421.255 17.415 3421.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3160.540 17.410 3160.600 ;
        RECT 225.010 3160.540 225.330 3160.600 ;
        RECT 17.090 3160.400 225.330 3160.540 ;
        RECT 17.090 3160.340 17.410 3160.400 ;
        RECT 225.010 3160.340 225.330 3160.400 ;
        RECT 225.010 1019.560 225.330 1019.620 ;
        RECT 732.850 1019.560 733.170 1019.620 ;
        RECT 225.010 1019.420 733.170 1019.560 ;
        RECT 225.010 1019.360 225.330 1019.420 ;
        RECT 732.850 1019.360 733.170 1019.420 ;
      LAYER via ;
        RECT 17.120 3160.340 17.380 3160.600 ;
        RECT 225.040 3160.340 225.300 3160.600 ;
        RECT 225.040 1019.360 225.300 1019.620 ;
        RECT 732.880 1019.360 733.140 1019.620 ;
      LAYER met2 ;
        RECT 17.120 3160.485 17.380 3160.630 ;
        RECT 17.110 3160.115 17.390 3160.485 ;
        RECT 225.040 3160.310 225.300 3160.630 ;
        RECT 225.100 1019.650 225.240 3160.310 ;
        RECT 225.040 1019.330 225.300 1019.650 ;
        RECT 732.880 1019.330 733.140 1019.650 ;
        RECT 732.940 999.330 733.080 1019.330 ;
        RECT 734.610 999.330 734.890 1000.000 ;
        RECT 732.940 999.190 734.890 999.330 ;
        RECT 734.610 996.000 734.890 999.190 ;
      LAYER via2 ;
        RECT 17.110 3160.160 17.390 3160.440 ;
      LAYER met3 ;
        RECT -4.800 3160.450 2.400 3160.900 ;
        RECT 17.085 3160.450 17.415 3160.465 ;
        RECT -4.800 3160.150 17.415 3160.450 ;
        RECT -4.800 3159.700 2.400 3160.150 ;
        RECT 17.085 3160.135 17.415 3160.150 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2898.400 16.950 2898.460 ;
        RECT 225.470 2898.400 225.790 2898.460 ;
        RECT 16.630 2898.260 225.790 2898.400 ;
        RECT 16.630 2898.200 16.950 2898.260 ;
        RECT 225.470 2898.200 225.790 2898.260 ;
        RECT 225.470 1019.220 225.790 1019.280 ;
        RECT 754.470 1019.220 754.790 1019.280 ;
        RECT 225.470 1019.080 754.790 1019.220 ;
        RECT 225.470 1019.020 225.790 1019.080 ;
        RECT 754.470 1019.020 754.790 1019.080 ;
      LAYER via ;
        RECT 16.660 2898.200 16.920 2898.460 ;
        RECT 225.500 2898.200 225.760 2898.460 ;
        RECT 225.500 1019.020 225.760 1019.280 ;
        RECT 754.500 1019.020 754.760 1019.280 ;
      LAYER met2 ;
        RECT 16.650 2899.675 16.930 2900.045 ;
        RECT 16.720 2898.490 16.860 2899.675 ;
        RECT 16.660 2898.170 16.920 2898.490 ;
        RECT 225.500 2898.170 225.760 2898.490 ;
        RECT 225.560 1019.310 225.700 2898.170 ;
        RECT 225.500 1018.990 225.760 1019.310 ;
        RECT 754.500 1018.990 754.760 1019.310 ;
        RECT 754.560 999.330 754.700 1018.990 ;
        RECT 755.770 999.330 756.050 1000.000 ;
        RECT 754.560 999.190 756.050 999.330 ;
        RECT 755.770 996.000 756.050 999.190 ;
      LAYER via2 ;
        RECT 16.650 2899.720 16.930 2900.000 ;
      LAYER met3 ;
        RECT -4.800 2900.010 2.400 2900.460 ;
        RECT 16.625 2900.010 16.955 2900.025 ;
        RECT -4.800 2899.710 16.955 2900.010 ;
        RECT -4.800 2899.260 2.400 2899.710 ;
        RECT 16.625 2899.695 16.955 2899.710 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2635.920 17.410 2635.980 ;
        RECT 772.870 2635.920 773.190 2635.980 ;
        RECT 17.090 2635.780 773.190 2635.920 ;
        RECT 17.090 2635.720 17.410 2635.780 ;
        RECT 772.870 2635.720 773.190 2635.780 ;
      LAYER via ;
        RECT 17.120 2635.720 17.380 2635.980 ;
        RECT 772.900 2635.720 773.160 2635.980 ;
      LAYER met2 ;
        RECT 17.110 2639.235 17.390 2639.605 ;
        RECT 17.180 2636.010 17.320 2639.235 ;
        RECT 17.120 2635.690 17.380 2636.010 ;
        RECT 772.900 2635.690 773.160 2636.010 ;
        RECT 772.960 1048.870 773.100 2635.690 ;
        RECT 772.960 1048.730 775.400 1048.870 ;
        RECT 775.260 999.330 775.400 1048.730 ;
        RECT 777.390 999.330 777.670 1000.000 ;
        RECT 775.260 999.190 777.670 999.330 ;
        RECT 777.390 996.000 777.670 999.190 ;
      LAYER via2 ;
        RECT 17.110 2639.280 17.390 2639.560 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 17.085 2639.570 17.415 2639.585 ;
        RECT -4.800 2639.270 17.415 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 17.085 2639.255 17.415 2639.270 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2373.780 17.410 2373.840 ;
        RECT 793.570 2373.780 793.890 2373.840 ;
        RECT 17.090 2373.640 793.890 2373.780 ;
        RECT 17.090 2373.580 17.410 2373.640 ;
        RECT 793.570 2373.580 793.890 2373.640 ;
      LAYER via ;
        RECT 17.120 2373.580 17.380 2373.840 ;
        RECT 793.600 2373.580 793.860 2373.840 ;
      LAYER met2 ;
        RECT 17.110 2378.115 17.390 2378.485 ;
        RECT 17.180 2373.870 17.320 2378.115 ;
        RECT 17.120 2373.550 17.380 2373.870 ;
        RECT 793.600 2373.550 793.860 2373.870 ;
        RECT 793.660 1048.870 793.800 2373.550 ;
        RECT 793.660 1048.730 796.560 1048.870 ;
        RECT 796.420 999.330 796.560 1048.730 ;
        RECT 798.550 999.330 798.830 1000.000 ;
        RECT 796.420 999.190 798.830 999.330 ;
        RECT 798.550 996.000 798.830 999.190 ;
      LAYER via2 ;
        RECT 17.110 2378.160 17.390 2378.440 ;
      LAYER met3 ;
        RECT -4.800 2378.450 2.400 2378.900 ;
        RECT 17.085 2378.450 17.415 2378.465 ;
        RECT -4.800 2378.150 17.415 2378.450 ;
        RECT -4.800 2377.700 2.400 2378.150 ;
        RECT 17.085 2378.135 17.415 2378.150 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2111.640 17.410 2111.700 ;
        RECT 814.270 2111.640 814.590 2111.700 ;
        RECT 17.090 2111.500 814.590 2111.640 ;
        RECT 17.090 2111.440 17.410 2111.500 ;
        RECT 814.270 2111.440 814.590 2111.500 ;
      LAYER via ;
        RECT 17.120 2111.440 17.380 2111.700 ;
        RECT 814.300 2111.440 814.560 2111.700 ;
      LAYER met2 ;
        RECT 17.110 2117.675 17.390 2118.045 ;
        RECT 17.180 2111.730 17.320 2117.675 ;
        RECT 17.120 2111.410 17.380 2111.730 ;
        RECT 814.300 2111.410 814.560 2111.730 ;
        RECT 814.360 1048.870 814.500 2111.410 ;
        RECT 814.360 1048.730 817.720 1048.870 ;
        RECT 817.580 999.330 817.720 1048.730 ;
        RECT 819.710 999.330 819.990 1000.000 ;
        RECT 817.580 999.190 819.990 999.330 ;
        RECT 819.710 996.000 819.990 999.190 ;
      LAYER via2 ;
        RECT 17.110 2117.720 17.390 2118.000 ;
      LAYER met3 ;
        RECT -4.800 2118.010 2.400 2118.460 ;
        RECT 17.085 2118.010 17.415 2118.025 ;
        RECT -4.800 2117.710 17.415 2118.010 ;
        RECT -4.800 2117.260 2.400 2117.710 ;
        RECT 17.085 2117.695 17.415 2117.710 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 247.090 1001.880 247.410 1001.940 ;
        RECT 2900.830 1001.880 2901.150 1001.940 ;
        RECT 247.090 1001.740 2901.150 1001.880 ;
        RECT 247.090 1001.680 247.410 1001.740 ;
        RECT 2900.830 1001.680 2901.150 1001.740 ;
      LAYER via ;
        RECT 247.120 1001.680 247.380 1001.940 ;
        RECT 2900.860 1001.680 2901.120 1001.940 ;
      LAYER met2 ;
        RECT 247.120 1001.650 247.380 1001.970 ;
        RECT 2900.860 1001.650 2901.120 1001.970 ;
        RECT 245.630 999.330 245.910 1000.000 ;
        RECT 247.180 999.330 247.320 1001.650 ;
        RECT 245.630 999.190 247.320 999.330 ;
        RECT 245.630 996.000 245.910 999.190 ;
        RECT 2900.920 430.965 2901.060 1001.650 ;
        RECT 2900.850 430.595 2901.130 430.965 ;
      LAYER via2 ;
        RECT 2900.850 430.640 2901.130 430.920 ;
      LAYER met3 ;
        RECT 2900.825 430.930 2901.155 430.945 ;
        RECT 2917.600 430.930 2924.800 431.380 ;
        RECT 2900.825 430.630 2924.800 430.930 ;
        RECT 2900.825 430.615 2901.155 430.630 ;
        RECT 2917.600 430.180 2924.800 430.630 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1856.300 17.870 1856.360 ;
        RECT 834.970 1856.300 835.290 1856.360 ;
        RECT 17.550 1856.160 835.290 1856.300 ;
        RECT 17.550 1856.100 17.870 1856.160 ;
        RECT 834.970 1856.100 835.290 1856.160 ;
      LAYER via ;
        RECT 17.580 1856.100 17.840 1856.360 ;
        RECT 835.000 1856.100 835.260 1856.360 ;
      LAYER met2 ;
        RECT 17.570 1856.555 17.850 1856.925 ;
        RECT 17.640 1856.390 17.780 1856.555 ;
        RECT 17.580 1856.070 17.840 1856.390 ;
        RECT 835.000 1856.070 835.260 1856.390 ;
        RECT 835.060 1048.870 835.200 1856.070 ;
        RECT 835.060 1048.730 838.880 1048.870 ;
        RECT 838.740 999.330 838.880 1048.730 ;
        RECT 840.870 999.330 841.150 1000.000 ;
        RECT 838.740 999.190 841.150 999.330 ;
        RECT 840.870 996.000 841.150 999.190 ;
      LAYER via2 ;
        RECT 17.570 1856.600 17.850 1856.880 ;
      LAYER met3 ;
        RECT -4.800 1856.890 2.400 1857.340 ;
        RECT 17.545 1856.890 17.875 1856.905 ;
        RECT -4.800 1856.590 17.875 1856.890 ;
        RECT -4.800 1856.140 2.400 1856.590 ;
        RECT 17.545 1856.575 17.875 1856.590 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1594.160 16.950 1594.220 ;
        RECT 862.570 1594.160 862.890 1594.220 ;
        RECT 16.630 1594.020 862.890 1594.160 ;
        RECT 16.630 1593.960 16.950 1594.020 ;
        RECT 862.570 1593.960 862.890 1594.020 ;
      LAYER via ;
        RECT 16.660 1593.960 16.920 1594.220 ;
        RECT 862.600 1593.960 862.860 1594.220 ;
      LAYER met2 ;
        RECT 16.650 1596.115 16.930 1596.485 ;
        RECT 16.720 1594.250 16.860 1596.115 ;
        RECT 16.660 1593.930 16.920 1594.250 ;
        RECT 862.600 1593.930 862.860 1594.250 ;
        RECT 862.660 1048.870 862.800 1593.930 ;
        RECT 862.660 1048.730 863.260 1048.870 ;
        RECT 862.490 999.330 862.770 1000.000 ;
        RECT 863.120 999.330 863.260 1048.730 ;
        RECT 862.490 999.190 863.260 999.330 ;
        RECT 862.490 996.000 862.770 999.190 ;
      LAYER via2 ;
        RECT 16.650 1596.160 16.930 1596.440 ;
      LAYER met3 ;
        RECT -4.800 1596.450 2.400 1596.900 ;
        RECT 16.625 1596.450 16.955 1596.465 ;
        RECT -4.800 1596.150 16.955 1596.450 ;
        RECT -4.800 1595.700 2.400 1596.150 ;
        RECT 16.625 1596.135 16.955 1596.150 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1332.020 15.570 1332.080 ;
        RECT 883.270 1332.020 883.590 1332.080 ;
        RECT 15.250 1331.880 883.590 1332.020 ;
        RECT 15.250 1331.820 15.570 1331.880 ;
        RECT 883.270 1331.820 883.590 1331.880 ;
      LAYER via ;
        RECT 15.280 1331.820 15.540 1332.080 ;
        RECT 883.300 1331.820 883.560 1332.080 ;
      LAYER met2 ;
        RECT 15.270 1335.675 15.550 1336.045 ;
        RECT 15.340 1332.110 15.480 1335.675 ;
        RECT 15.280 1331.790 15.540 1332.110 ;
        RECT 883.300 1331.790 883.560 1332.110 ;
        RECT 883.360 999.330 883.500 1331.790 ;
        RECT 883.650 999.330 883.930 1000.000 ;
        RECT 883.360 999.190 883.930 999.330 ;
        RECT 883.650 996.000 883.930 999.190 ;
      LAYER via2 ;
        RECT 15.270 1335.720 15.550 1336.000 ;
      LAYER met3 ;
        RECT -4.800 1336.010 2.400 1336.460 ;
        RECT 15.245 1336.010 15.575 1336.025 ;
        RECT -4.800 1335.710 15.575 1336.010 ;
        RECT -4.800 1335.260 2.400 1335.710 ;
        RECT 15.245 1335.695 15.575 1335.710 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1069.880 16.030 1069.940 ;
        RECT 900.290 1069.880 900.610 1069.940 ;
        RECT 15.710 1069.740 900.610 1069.880 ;
        RECT 15.710 1069.680 16.030 1069.740 ;
        RECT 900.290 1069.680 900.610 1069.740 ;
        RECT 900.290 1012.760 900.610 1012.820 ;
        RECT 903.970 1012.760 904.290 1012.820 ;
        RECT 900.290 1012.620 904.290 1012.760 ;
        RECT 900.290 1012.560 900.610 1012.620 ;
        RECT 903.970 1012.560 904.290 1012.620 ;
      LAYER via ;
        RECT 15.740 1069.680 16.000 1069.940 ;
        RECT 900.320 1069.680 900.580 1069.940 ;
        RECT 900.320 1012.560 900.580 1012.820 ;
        RECT 904.000 1012.560 904.260 1012.820 ;
      LAYER met2 ;
        RECT 15.730 1074.555 16.010 1074.925 ;
        RECT 15.800 1069.970 15.940 1074.555 ;
        RECT 15.740 1069.650 16.000 1069.970 ;
        RECT 900.320 1069.650 900.580 1069.970 ;
        RECT 900.380 1012.850 900.520 1069.650 ;
        RECT 900.320 1012.530 900.580 1012.850 ;
        RECT 904.000 1012.530 904.260 1012.850 ;
        RECT 904.060 999.330 904.200 1012.530 ;
        RECT 904.810 999.330 905.090 1000.000 ;
        RECT 904.060 999.190 905.090 999.330 ;
        RECT 904.810 996.000 905.090 999.190 ;
      LAYER via2 ;
        RECT 15.730 1074.600 16.010 1074.880 ;
      LAYER met3 ;
        RECT -4.800 1074.890 2.400 1075.340 ;
        RECT 15.705 1074.890 16.035 1074.905 ;
        RECT -4.800 1074.590 16.035 1074.890 ;
        RECT -4.800 1074.140 2.400 1074.590 ;
        RECT 15.705 1074.575 16.035 1074.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1004.260 16.490 1004.320 ;
        RECT 924.670 1004.260 924.990 1004.320 ;
        RECT 16.170 1004.120 924.990 1004.260 ;
        RECT 16.170 1004.060 16.490 1004.120 ;
        RECT 924.670 1004.060 924.990 1004.120 ;
      LAYER via ;
        RECT 16.200 1004.060 16.460 1004.320 ;
        RECT 924.700 1004.060 924.960 1004.320 ;
      LAYER met2 ;
        RECT 16.200 1004.030 16.460 1004.350 ;
        RECT 924.700 1004.030 924.960 1004.350 ;
        RECT 16.260 814.485 16.400 1004.030 ;
        RECT 924.760 999.330 924.900 1004.030 ;
        RECT 925.970 999.330 926.250 1000.000 ;
        RECT 924.760 999.190 926.250 999.330 ;
        RECT 925.970 996.000 926.250 999.190 ;
        RECT 16.190 814.115 16.470 814.485 ;
      LAYER via2 ;
        RECT 16.190 814.160 16.470 814.440 ;
      LAYER met3 ;
        RECT -4.800 814.450 2.400 814.900 ;
        RECT 16.165 814.450 16.495 814.465 ;
        RECT -4.800 814.150 16.495 814.450 ;
        RECT -4.800 813.700 2.400 814.150 ;
        RECT 16.165 814.135 16.495 814.150 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.850 1008.340 20.170 1008.400 ;
        RECT 945.830 1008.340 946.150 1008.400 ;
        RECT 19.850 1008.200 946.150 1008.340 ;
        RECT 19.850 1008.140 20.170 1008.200 ;
        RECT 945.830 1008.140 946.150 1008.200 ;
      LAYER via ;
        RECT 19.880 1008.140 20.140 1008.400 ;
        RECT 945.860 1008.140 946.120 1008.400 ;
      LAYER met2 ;
        RECT 19.880 1008.110 20.140 1008.430 ;
        RECT 945.860 1008.110 946.120 1008.430 ;
        RECT 19.940 553.365 20.080 1008.110 ;
        RECT 945.920 999.330 946.060 1008.110 ;
        RECT 947.130 999.330 947.410 1000.000 ;
        RECT 945.920 999.190 947.410 999.330 ;
        RECT 947.130 996.000 947.410 999.190 ;
        RECT 19.870 552.995 20.150 553.365 ;
      LAYER via2 ;
        RECT 19.870 553.040 20.150 553.320 ;
      LAYER met3 ;
        RECT -4.800 553.330 2.400 553.780 ;
        RECT 19.845 553.330 20.175 553.345 ;
        RECT -4.800 553.030 20.175 553.330 ;
        RECT -4.800 552.580 2.400 553.030 ;
        RECT 19.845 553.015 20.175 553.030 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 1003.240 18.790 1003.300 ;
        RECT 967.450 1003.240 967.770 1003.300 ;
        RECT 18.470 1003.100 967.770 1003.240 ;
        RECT 18.470 1003.040 18.790 1003.100 ;
        RECT 967.450 1003.040 967.770 1003.100 ;
      LAYER via ;
        RECT 18.500 1003.040 18.760 1003.300 ;
        RECT 967.480 1003.040 967.740 1003.300 ;
      LAYER met2 ;
        RECT 18.500 1003.010 18.760 1003.330 ;
        RECT 967.480 1003.010 967.740 1003.330 ;
        RECT 18.560 358.205 18.700 1003.010 ;
        RECT 967.540 999.330 967.680 1003.010 ;
        RECT 968.750 999.330 969.030 1000.000 ;
        RECT 967.540 999.190 969.030 999.330 ;
        RECT 968.750 996.000 969.030 999.190 ;
        RECT 18.490 357.835 18.770 358.205 ;
      LAYER via2 ;
        RECT 18.490 357.880 18.770 358.160 ;
      LAYER met3 ;
        RECT -4.800 358.170 2.400 358.620 ;
        RECT 18.465 358.170 18.795 358.185 ;
        RECT -4.800 357.870 18.795 358.170 ;
        RECT -4.800 357.420 2.400 357.870 ;
        RECT 18.465 357.855 18.795 357.870 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 1001.115 988.450 1001.485 ;
        RECT 988.240 999.330 988.380 1001.115 ;
        RECT 989.910 999.330 990.190 1000.000 ;
        RECT 988.240 999.190 990.190 999.330 ;
        RECT 989.910 996.000 990.190 999.190 ;
      LAYER via2 ;
        RECT 988.170 1001.160 988.450 1001.440 ;
      LAYER met3 ;
        RECT 17.750 1001.450 18.130 1001.460 ;
        RECT 988.145 1001.450 988.475 1001.465 ;
        RECT 17.750 1001.150 988.475 1001.450 ;
        RECT 17.750 1001.140 18.130 1001.150 ;
        RECT 988.145 1001.135 988.475 1001.150 ;
        RECT -4.800 162.330 2.400 162.780 ;
        RECT 17.750 162.330 18.130 162.340 ;
        RECT -4.800 162.030 18.130 162.330 ;
        RECT -4.800 161.580 2.400 162.030 ;
        RECT 17.750 162.020 18.130 162.030 ;
      LAYER via3 ;
        RECT 17.780 1001.140 18.100 1001.460 ;
        RECT 17.780 162.020 18.100 162.340 ;
      LAYER met4 ;
        RECT 17.775 1001.135 18.105 1001.465 ;
        RECT 17.790 162.345 18.090 1001.135 ;
        RECT 17.775 162.015 18.105 162.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 268.250 1009.360 268.570 1009.420 ;
        RECT 1100.850 1009.360 1101.170 1009.420 ;
        RECT 268.250 1009.220 1101.170 1009.360 ;
        RECT 268.250 1009.160 268.570 1009.220 ;
        RECT 1100.850 1009.160 1101.170 1009.220 ;
        RECT 1100.850 634.680 1101.170 634.740 ;
        RECT 2899.910 634.680 2900.230 634.740 ;
        RECT 1100.850 634.540 2900.230 634.680 ;
        RECT 1100.850 634.480 1101.170 634.540 ;
        RECT 2899.910 634.480 2900.230 634.540 ;
      LAYER via ;
        RECT 268.280 1009.160 268.540 1009.420 ;
        RECT 1100.880 1009.160 1101.140 1009.420 ;
        RECT 1100.880 634.480 1101.140 634.740 ;
        RECT 2899.940 634.480 2900.200 634.740 ;
      LAYER met2 ;
        RECT 268.280 1009.130 268.540 1009.450 ;
        RECT 1100.880 1009.130 1101.140 1009.450 ;
        RECT 266.790 999.330 267.070 1000.000 ;
        RECT 268.340 999.330 268.480 1009.130 ;
        RECT 266.790 999.190 268.480 999.330 ;
        RECT 266.790 996.000 267.070 999.190 ;
        RECT 1100.940 634.770 1101.080 1009.130 ;
        RECT 1100.880 634.450 1101.140 634.770 ;
        RECT 2899.940 634.450 2900.200 634.770 ;
        RECT 2900.000 630.205 2900.140 634.450 ;
        RECT 2899.930 629.835 2900.210 630.205 ;
      LAYER via2 ;
        RECT 2899.930 629.880 2900.210 630.160 ;
      LAYER met3 ;
        RECT 2899.905 630.170 2900.235 630.185 ;
        RECT 2917.600 630.170 2924.800 630.620 ;
        RECT 2899.905 629.870 2924.800 630.170 ;
        RECT 2899.905 629.855 2900.235 629.870 ;
        RECT 2917.600 629.420 2924.800 629.870 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.950 1010.380 289.270 1010.440 ;
        RECT 1102.230 1010.380 1102.550 1010.440 ;
        RECT 288.950 1010.240 1102.550 1010.380 ;
        RECT 288.950 1010.180 289.270 1010.240 ;
        RECT 1102.230 1010.180 1102.550 1010.240 ;
        RECT 1102.230 834.940 1102.550 835.000 ;
        RECT 2899.910 834.940 2900.230 835.000 ;
        RECT 1102.230 834.800 2900.230 834.940 ;
        RECT 1102.230 834.740 1102.550 834.800 ;
        RECT 2899.910 834.740 2900.230 834.800 ;
      LAYER via ;
        RECT 288.980 1010.180 289.240 1010.440 ;
        RECT 1102.260 1010.180 1102.520 1010.440 ;
        RECT 1102.260 834.740 1102.520 835.000 ;
        RECT 2899.940 834.740 2900.200 835.000 ;
      LAYER met2 ;
        RECT 288.980 1010.150 289.240 1010.470 ;
        RECT 1102.260 1010.150 1102.520 1010.470 ;
        RECT 287.950 999.330 288.230 1000.000 ;
        RECT 289.040 999.330 289.180 1010.150 ;
        RECT 287.950 999.190 289.180 999.330 ;
        RECT 287.950 996.000 288.230 999.190 ;
        RECT 1102.320 835.030 1102.460 1010.150 ;
        RECT 1102.260 834.710 1102.520 835.030 ;
        RECT 2899.940 834.710 2900.200 835.030 ;
        RECT 2900.000 829.445 2900.140 834.710 ;
        RECT 2899.930 829.075 2900.210 829.445 ;
      LAYER via2 ;
        RECT 2899.930 829.120 2900.210 829.400 ;
      LAYER met3 ;
        RECT 2899.905 829.410 2900.235 829.425 ;
        RECT 2917.600 829.410 2924.800 829.860 ;
        RECT 2899.905 829.110 2924.800 829.410 ;
        RECT 2899.905 829.095 2900.235 829.110 ;
        RECT 2917.600 828.660 2924.800 829.110 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 307.810 1028.400 308.130 1028.460 ;
        RECT 2900.830 1028.400 2901.150 1028.460 ;
        RECT 307.810 1028.260 2901.150 1028.400 ;
        RECT 307.810 1028.200 308.130 1028.260 ;
        RECT 2900.830 1028.200 2901.150 1028.260 ;
      LAYER via ;
        RECT 307.840 1028.200 308.100 1028.460 ;
        RECT 2900.860 1028.200 2901.120 1028.460 ;
      LAYER met2 ;
        RECT 307.840 1028.170 308.100 1028.490 ;
        RECT 2900.850 1028.315 2901.130 1028.685 ;
        RECT 2900.860 1028.170 2901.120 1028.315 ;
        RECT 307.900 999.330 308.040 1028.170 ;
        RECT 309.570 999.330 309.850 1000.000 ;
        RECT 307.900 999.190 309.850 999.330 ;
        RECT 309.570 996.000 309.850 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1028.360 2901.130 1028.640 ;
      LAYER met3 ;
        RECT 2900.825 1028.650 2901.155 1028.665 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2900.825 1028.350 2924.800 1028.650 ;
        RECT 2900.825 1028.335 2901.155 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 1221.520 324.690 1221.580 ;
        RECT 2900.830 1221.520 2901.150 1221.580 ;
        RECT 324.370 1221.380 2901.150 1221.520 ;
        RECT 324.370 1221.320 324.690 1221.380 ;
        RECT 2900.830 1221.320 2901.150 1221.380 ;
      LAYER via ;
        RECT 324.400 1221.320 324.660 1221.580 ;
        RECT 2900.860 1221.320 2901.120 1221.580 ;
      LAYER met2 ;
        RECT 2900.850 1227.555 2901.130 1227.925 ;
        RECT 2900.920 1221.610 2901.060 1227.555 ;
        RECT 324.400 1221.290 324.660 1221.610 ;
        RECT 2900.860 1221.290 2901.120 1221.610 ;
        RECT 324.460 1048.870 324.600 1221.290 ;
        RECT 324.460 1048.730 329.200 1048.870 ;
        RECT 329.060 999.330 329.200 1048.730 ;
        RECT 330.730 999.330 331.010 1000.000 ;
        RECT 329.060 999.190 331.010 999.330 ;
        RECT 330.730 996.000 331.010 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1227.600 2901.130 1227.880 ;
      LAYER met3 ;
        RECT 2900.825 1227.890 2901.155 1227.905 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2900.825 1227.590 2924.800 1227.890 ;
        RECT 2900.825 1227.575 2901.155 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.970 1490.800 352.290 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 351.970 1490.660 2901.150 1490.800 ;
        RECT 351.970 1490.600 352.290 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 352.000 1490.600 352.260 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1493.435 2901.130 1493.805 ;
        RECT 2900.920 1490.890 2901.060 1493.435 ;
        RECT 352.000 1490.570 352.260 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 352.060 1048.870 352.200 1490.570 ;
        RECT 352.060 1048.730 352.660 1048.870 ;
        RECT 351.890 999.330 352.170 1000.000 ;
        RECT 352.520 999.330 352.660 1048.730 ;
        RECT 351.890 999.190 352.660 999.330 ;
        RECT 351.890 996.000 352.170 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1493.480 2901.130 1493.760 ;
      LAYER met3 ;
        RECT 2900.825 1493.770 2901.155 1493.785 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2900.825 1493.470 2924.800 1493.770 ;
        RECT 2900.825 1493.455 2901.155 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 1759.740 372.990 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 372.670 1759.600 2901.150 1759.740 ;
        RECT 372.670 1759.540 372.990 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
      LAYER via ;
        RECT 372.700 1759.540 372.960 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
      LAYER met2 ;
        RECT 372.700 1759.510 372.960 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 372.760 999.330 372.900 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 373.050 999.330 373.330 1000.000 ;
        RECT 372.760 999.190 373.330 999.330 ;
        RECT 373.050 996.000 373.330 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.370 2021.880 393.690 2021.940 ;
        RECT 2899.910 2021.880 2900.230 2021.940 ;
        RECT 393.370 2021.740 2900.230 2021.880 ;
        RECT 393.370 2021.680 393.690 2021.740 ;
        RECT 2899.910 2021.680 2900.230 2021.740 ;
      LAYER via ;
        RECT 393.400 2021.680 393.660 2021.940 ;
        RECT 2899.940 2021.680 2900.200 2021.940 ;
      LAYER met2 ;
        RECT 2899.930 2024.515 2900.210 2024.885 ;
        RECT 2900.000 2021.970 2900.140 2024.515 ;
        RECT 393.400 2021.650 393.660 2021.970 ;
        RECT 2899.940 2021.650 2900.200 2021.970 ;
        RECT 393.460 999.330 393.600 2021.650 ;
        RECT 394.670 999.330 394.950 1000.000 ;
        RECT 393.460 999.190 394.950 999.330 ;
        RECT 394.670 996.000 394.950 999.190 ;
      LAYER via2 ;
        RECT 2899.930 2024.560 2900.210 2024.840 ;
      LAYER met3 ;
        RECT 2899.905 2024.850 2900.235 2024.865 ;
        RECT 2917.600 2024.850 2924.800 2025.300 ;
        RECT 2899.905 2024.550 2924.800 2024.850 ;
        RECT 2899.905 2024.535 2900.235 2024.550 ;
        RECT 2917.600 2024.100 2924.800 2024.550 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 212.130 1000.860 212.450 1000.920 ;
        RECT 2903.130 1000.860 2903.450 1000.920 ;
        RECT 212.130 1000.720 2903.450 1000.860 ;
        RECT 212.130 1000.660 212.450 1000.720 ;
        RECT 2903.130 1000.660 2903.450 1000.720 ;
      LAYER via ;
        RECT 212.160 1000.660 212.420 1000.920 ;
        RECT 2903.160 1000.660 2903.420 1000.920 ;
      LAYER met2 ;
        RECT 212.160 1000.630 212.420 1000.950 ;
        RECT 2903.160 1000.630 2903.420 1000.950 ;
        RECT 210.210 999.330 210.490 1000.000 ;
        RECT 212.220 999.330 212.360 1000.630 ;
        RECT 210.210 999.190 212.360 999.330 ;
        RECT 210.210 996.000 210.490 999.190 ;
        RECT 2903.220 165.765 2903.360 1000.630 ;
        RECT 2903.150 165.395 2903.430 165.765 ;
      LAYER via2 ;
        RECT 2903.150 165.440 2903.430 165.720 ;
      LAYER met3 ;
        RECT 2903.125 165.730 2903.455 165.745 ;
        RECT 2917.600 165.730 2924.800 166.180 ;
        RECT 2903.125 165.430 2924.800 165.730 ;
        RECT 2903.125 165.415 2903.455 165.430 ;
        RECT 2917.600 164.980 2924.800 165.430 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 2422.060 421.290 2422.120 ;
        RECT 2900.830 2422.060 2901.150 2422.120 ;
        RECT 420.970 2421.920 2901.150 2422.060 ;
        RECT 420.970 2421.860 421.290 2421.920 ;
        RECT 2900.830 2421.860 2901.150 2421.920 ;
      LAYER via ;
        RECT 421.000 2421.860 421.260 2422.120 ;
        RECT 2900.860 2421.860 2901.120 2422.120 ;
      LAYER met2 ;
        RECT 2900.850 2422.995 2901.130 2423.365 ;
        RECT 2900.920 2422.150 2901.060 2422.995 ;
        RECT 421.000 2421.830 421.260 2422.150 ;
        RECT 2900.860 2421.830 2901.120 2422.150 ;
        RECT 421.060 999.330 421.200 2421.830 ;
        RECT 422.730 999.330 423.010 1000.000 ;
        RECT 421.060 999.190 423.010 999.330 ;
        RECT 422.730 996.000 423.010 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2423.040 2901.130 2423.320 ;
      LAYER met3 ;
        RECT 2900.825 2423.330 2901.155 2423.345 ;
        RECT 2917.600 2423.330 2924.800 2423.780 ;
        RECT 2900.825 2423.030 2924.800 2423.330 ;
        RECT 2900.825 2423.015 2901.155 2423.030 ;
        RECT 2917.600 2422.580 2924.800 2423.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 2684.200 441.990 2684.260 ;
        RECT 2899.450 2684.200 2899.770 2684.260 ;
        RECT 441.670 2684.060 2899.770 2684.200 ;
        RECT 441.670 2684.000 441.990 2684.060 ;
        RECT 2899.450 2684.000 2899.770 2684.060 ;
      LAYER via ;
        RECT 441.700 2684.000 441.960 2684.260 ;
        RECT 2899.480 2684.000 2899.740 2684.260 ;
      LAYER met2 ;
        RECT 2899.470 2688.875 2899.750 2689.245 ;
        RECT 2899.540 2684.290 2899.680 2688.875 ;
        RECT 441.700 2683.970 441.960 2684.290 ;
        RECT 2899.480 2683.970 2899.740 2684.290 ;
        RECT 441.760 1048.870 441.900 2683.970 ;
        RECT 441.760 1048.730 442.360 1048.870 ;
        RECT 442.220 999.330 442.360 1048.730 ;
        RECT 443.890 999.330 444.170 1000.000 ;
        RECT 442.220 999.190 444.170 999.330 ;
        RECT 443.890 996.000 444.170 999.190 ;
      LAYER via2 ;
        RECT 2899.470 2688.920 2899.750 2689.200 ;
      LAYER met3 ;
        RECT 2899.445 2689.210 2899.775 2689.225 ;
        RECT 2917.600 2689.210 2924.800 2689.660 ;
        RECT 2899.445 2688.910 2924.800 2689.210 ;
        RECT 2899.445 2688.895 2899.775 2688.910 ;
        RECT 2917.600 2688.460 2924.800 2688.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 2953.480 462.690 2953.540 ;
        RECT 2900.830 2953.480 2901.150 2953.540 ;
        RECT 462.370 2953.340 2901.150 2953.480 ;
        RECT 462.370 2953.280 462.690 2953.340 ;
        RECT 2900.830 2953.280 2901.150 2953.340 ;
      LAYER via ;
        RECT 462.400 2953.280 462.660 2953.540 ;
        RECT 2900.860 2953.280 2901.120 2953.540 ;
      LAYER met2 ;
        RECT 2900.850 2954.755 2901.130 2955.125 ;
        RECT 2900.920 2953.570 2901.060 2954.755 ;
        RECT 462.400 2953.250 462.660 2953.570 ;
        RECT 2900.860 2953.250 2901.120 2953.570 ;
        RECT 462.460 1048.870 462.600 2953.250 ;
        RECT 462.460 1048.730 463.520 1048.870 ;
        RECT 463.380 999.330 463.520 1048.730 ;
        RECT 465.510 999.330 465.790 1000.000 ;
        RECT 463.380 999.190 465.790 999.330 ;
        RECT 465.510 996.000 465.790 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2954.800 2901.130 2955.080 ;
      LAYER met3 ;
        RECT 2900.825 2955.090 2901.155 2955.105 ;
        RECT 2917.600 2955.090 2924.800 2955.540 ;
        RECT 2900.825 2954.790 2924.800 2955.090 ;
        RECT 2900.825 2954.775 2901.155 2954.790 ;
        RECT 2917.600 2954.340 2924.800 2954.790 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 3215.620 483.390 3215.680 ;
        RECT 2900.830 3215.620 2901.150 3215.680 ;
        RECT 483.070 3215.480 2901.150 3215.620 ;
        RECT 483.070 3215.420 483.390 3215.480 ;
        RECT 2900.830 3215.420 2901.150 3215.480 ;
      LAYER via ;
        RECT 483.100 3215.420 483.360 3215.680 ;
        RECT 2900.860 3215.420 2901.120 3215.680 ;
      LAYER met2 ;
        RECT 2900.850 3219.955 2901.130 3220.325 ;
        RECT 2900.920 3215.710 2901.060 3219.955 ;
        RECT 483.100 3215.390 483.360 3215.710 ;
        RECT 2900.860 3215.390 2901.120 3215.710 ;
        RECT 483.160 1048.870 483.300 3215.390 ;
        RECT 483.160 1048.730 484.680 1048.870 ;
        RECT 484.540 999.330 484.680 1048.730 ;
        RECT 486.670 999.330 486.950 1000.000 ;
        RECT 484.540 999.190 486.950 999.330 ;
        RECT 486.670 996.000 486.950 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3220.000 2901.130 3220.280 ;
      LAYER met3 ;
        RECT 2900.825 3220.290 2901.155 3220.305 ;
        RECT 2917.600 3220.290 2924.800 3220.740 ;
        RECT 2900.825 3219.990 2924.800 3220.290 ;
        RECT 2900.825 3219.975 2901.155 3219.990 ;
        RECT 2917.600 3219.540 2924.800 3219.990 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 3484.900 504.090 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 503.770 3484.760 2901.150 3484.900 ;
        RECT 503.770 3484.700 504.090 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 503.800 3484.700 504.060 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3485.835 2901.130 3486.205 ;
        RECT 2900.920 3484.990 2901.060 3485.835 ;
        RECT 503.800 3484.670 504.060 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 503.860 1048.870 504.000 3484.670 ;
        RECT 503.860 1048.730 505.840 1048.870 ;
        RECT 505.700 999.330 505.840 1048.730 ;
        RECT 507.830 999.330 508.110 1000.000 ;
        RECT 505.700 999.190 508.110 999.330 ;
        RECT 507.830 996.000 508.110 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3485.880 2901.130 3486.160 ;
      LAYER met3 ;
        RECT 2900.825 3486.170 2901.155 3486.185 ;
        RECT 2917.600 3486.170 2924.800 3486.620 ;
        RECT 2900.825 3485.870 2924.800 3486.170 ;
        RECT 2900.825 3485.855 2901.155 3485.870 ;
        RECT 2917.600 3485.420 2924.800 3485.870 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 3501.900 524.790 3501.960 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 524.470 3501.760 2636.190 3501.900 ;
        RECT 524.470 3501.700 524.790 3501.760 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
      LAYER via ;
        RECT 524.500 3501.700 524.760 3501.960 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.990 2636.100 3517.600 ;
        RECT 524.500 3501.670 524.760 3501.990 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 524.560 1000.570 524.700 3501.670 ;
        RECT 524.560 1000.430 527.000 1000.570 ;
        RECT 526.860 999.330 527.000 1000.430 ;
        RECT 528.990 999.330 529.270 1000.000 ;
        RECT 526.860 999.190 529.270 999.330 ;
        RECT 528.990 996.000 529.270 999.190 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 3502.580 545.490 3502.640 ;
        RECT 2311.570 3502.580 2311.890 3502.640 ;
        RECT 545.170 3502.440 2311.890 3502.580 ;
        RECT 545.170 3502.380 545.490 3502.440 ;
        RECT 2311.570 3502.380 2311.890 3502.440 ;
      LAYER via ;
        RECT 545.200 3502.380 545.460 3502.640 ;
        RECT 2311.600 3502.380 2311.860 3502.640 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3502.670 2311.800 3517.600 ;
        RECT 545.200 3502.350 545.460 3502.670 ;
        RECT 2311.600 3502.350 2311.860 3502.670 ;
        RECT 545.260 1048.870 545.400 3502.350 ;
        RECT 545.260 1048.730 549.080 1048.870 ;
        RECT 548.940 999.330 549.080 1048.730 ;
        RECT 550.610 999.330 550.890 1000.000 ;
        RECT 548.940 999.190 550.890 999.330 ;
        RECT 550.610 996.000 550.890 999.190 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 3503.260 566.190 3503.320 ;
        RECT 1987.270 3503.260 1987.590 3503.320 ;
        RECT 565.870 3503.120 1987.590 3503.260 ;
        RECT 565.870 3503.060 566.190 3503.120 ;
        RECT 1987.270 3503.060 1987.590 3503.120 ;
      LAYER via ;
        RECT 565.900 3503.060 566.160 3503.320 ;
        RECT 1987.300 3503.060 1987.560 3503.320 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3503.350 1987.500 3517.600 ;
        RECT 565.900 3503.030 566.160 3503.350 ;
        RECT 1987.300 3503.030 1987.560 3503.350 ;
        RECT 565.960 1048.870 566.100 3503.030 ;
        RECT 565.960 1048.730 570.240 1048.870 ;
        RECT 570.100 999.330 570.240 1048.730 ;
        RECT 571.770 999.330 572.050 1000.000 ;
        RECT 570.100 999.190 572.050 999.330 ;
        RECT 571.770 996.000 572.050 999.190 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 3503.940 586.890 3504.000 ;
        RECT 1662.510 3503.940 1662.830 3504.000 ;
        RECT 586.570 3503.800 1662.830 3503.940 ;
        RECT 586.570 3503.740 586.890 3503.800 ;
        RECT 1662.510 3503.740 1662.830 3503.800 ;
      LAYER via ;
        RECT 586.600 3503.740 586.860 3504.000 ;
        RECT 1662.540 3503.740 1662.800 3504.000 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3504.030 1662.740 3517.600 ;
        RECT 586.600 3503.710 586.860 3504.030 ;
        RECT 1662.540 3503.710 1662.800 3504.030 ;
        RECT 586.660 1048.870 586.800 3503.710 ;
        RECT 586.660 1048.730 591.400 1048.870 ;
        RECT 591.260 999.330 591.400 1048.730 ;
        RECT 592.930 999.330 593.210 1000.000 ;
        RECT 591.260 999.190 593.210 999.330 ;
        RECT 592.930 996.000 593.210 999.190 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 969.750 3501.220 970.070 3501.280 ;
        RECT 1338.210 3501.220 1338.530 3501.280 ;
        RECT 969.750 3501.080 1338.530 3501.220 ;
        RECT 969.750 3501.020 970.070 3501.080 ;
        RECT 1338.210 3501.020 1338.530 3501.080 ;
        RECT 614.630 1017.520 614.950 1017.580 ;
        RECT 969.750 1017.520 970.070 1017.580 ;
        RECT 614.630 1017.380 970.070 1017.520 ;
        RECT 614.630 1017.320 614.950 1017.380 ;
        RECT 969.750 1017.320 970.070 1017.380 ;
      LAYER via ;
        RECT 969.780 3501.020 970.040 3501.280 ;
        RECT 1338.240 3501.020 1338.500 3501.280 ;
        RECT 614.660 1017.320 614.920 1017.580 ;
        RECT 969.780 1017.320 970.040 1017.580 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3501.310 1338.440 3517.600 ;
        RECT 969.780 3500.990 970.040 3501.310 ;
        RECT 1338.240 3500.990 1338.500 3501.310 ;
        RECT 969.840 1017.610 969.980 3500.990 ;
        RECT 614.660 1017.290 614.920 1017.610 ;
        RECT 969.780 1017.290 970.040 1017.610 ;
        RECT 614.090 999.330 614.370 1000.000 ;
        RECT 614.720 999.330 614.860 1017.290 ;
        RECT 614.090 999.190 614.860 999.330 ;
        RECT 614.090 996.000 614.370 999.190 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 233.290 1001.540 233.610 1001.600 ;
        RECT 2904.510 1001.540 2904.830 1001.600 ;
        RECT 233.290 1001.400 2904.830 1001.540 ;
        RECT 233.290 1001.340 233.610 1001.400 ;
        RECT 2904.510 1001.340 2904.830 1001.400 ;
      LAYER via ;
        RECT 233.320 1001.340 233.580 1001.600 ;
        RECT 2904.540 1001.340 2904.800 1001.600 ;
      LAYER met2 ;
        RECT 233.320 1001.310 233.580 1001.630 ;
        RECT 2904.540 1001.310 2904.800 1001.630 ;
        RECT 231.370 999.330 231.650 1000.000 ;
        RECT 233.380 999.330 233.520 1001.310 ;
        RECT 231.370 999.190 233.520 999.330 ;
        RECT 231.370 996.000 231.650 999.190 ;
        RECT 2904.600 365.005 2904.740 1001.310 ;
        RECT 2904.530 364.635 2904.810 365.005 ;
      LAYER via2 ;
        RECT 2904.530 364.680 2904.810 364.960 ;
      LAYER met3 ;
        RECT 2904.505 364.970 2904.835 364.985 ;
        RECT 2917.600 364.970 2924.800 365.420 ;
        RECT 2904.505 364.670 2924.800 364.970 ;
        RECT 2904.505 364.655 2904.835 364.670 ;
        RECT 2917.600 364.220 2924.800 364.670 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 969.290 3498.500 969.610 3498.560 ;
        RECT 1013.910 3498.500 1014.230 3498.560 ;
        RECT 969.290 3498.360 1014.230 3498.500 ;
        RECT 969.290 3498.300 969.610 3498.360 ;
        RECT 1013.910 3498.300 1014.230 3498.360 ;
        RECT 634.870 1017.180 635.190 1017.240 ;
        RECT 969.290 1017.180 969.610 1017.240 ;
        RECT 634.870 1017.040 969.610 1017.180 ;
        RECT 634.870 1016.980 635.190 1017.040 ;
        RECT 969.290 1016.980 969.610 1017.040 ;
      LAYER via ;
        RECT 969.320 3498.300 969.580 3498.560 ;
        RECT 1013.940 3498.300 1014.200 3498.560 ;
        RECT 634.900 1016.980 635.160 1017.240 ;
        RECT 969.320 1016.980 969.580 1017.240 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3498.590 1014.140 3517.600 ;
        RECT 969.320 3498.270 969.580 3498.590 ;
        RECT 1013.940 3498.270 1014.200 3498.590 ;
        RECT 969.380 1017.270 969.520 3498.270 ;
        RECT 634.900 1016.950 635.160 1017.270 ;
        RECT 969.320 1016.950 969.580 1017.270 ;
        RECT 634.960 999.330 635.100 1016.950 ;
        RECT 635.250 999.330 635.530 1000.000 ;
        RECT 634.960 999.190 635.530 999.330 ;
        RECT 635.250 996.000 635.530 999.190 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 658.330 1011.060 658.650 1011.120 ;
        RECT 683.170 1011.060 683.490 1011.120 ;
        RECT 658.330 1010.920 683.490 1011.060 ;
        RECT 658.330 1010.860 658.650 1010.920 ;
        RECT 683.170 1010.860 683.490 1010.920 ;
      LAYER via ;
        RECT 658.360 1010.860 658.620 1011.120 ;
        RECT 683.200 1010.860 683.460 1011.120 ;
      LAYER met2 ;
        RECT 683.260 3517.910 688.460 3518.050 ;
        RECT 683.260 1011.150 683.400 3517.910 ;
        RECT 688.320 3517.370 688.460 3517.910 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.320 3517.230 689.380 3517.370 ;
        RECT 658.360 1010.830 658.620 1011.150 ;
        RECT 683.200 1010.830 683.460 1011.150 ;
        RECT 656.870 999.330 657.150 1000.000 ;
        RECT 658.420 999.330 658.560 1010.830 ;
        RECT 656.870 999.190 658.560 999.330 ;
        RECT 656.870 996.000 657.150 999.190 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 3515.160 359.190 3515.220 ;
        RECT 364.850 3515.160 365.170 3515.220 ;
        RECT 358.870 3515.020 365.170 3515.160 ;
        RECT 358.870 3514.960 359.190 3515.020 ;
        RECT 364.850 3514.960 365.170 3515.020 ;
        RECT 358.870 1010.720 359.190 1010.780 ;
        RECT 677.190 1010.720 677.510 1010.780 ;
        RECT 358.870 1010.580 677.510 1010.720 ;
        RECT 358.870 1010.520 359.190 1010.580 ;
        RECT 677.190 1010.520 677.510 1010.580 ;
      LAYER via ;
        RECT 358.900 3514.960 359.160 3515.220 ;
        RECT 364.880 3514.960 365.140 3515.220 ;
        RECT 358.900 1010.520 359.160 1010.780 ;
        RECT 677.220 1010.520 677.480 1010.780 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3515.250 365.080 3517.600 ;
        RECT 358.900 3514.930 359.160 3515.250 ;
        RECT 364.880 3514.930 365.140 3515.250 ;
        RECT 358.960 1010.810 359.100 3514.930 ;
        RECT 358.900 1010.490 359.160 1010.810 ;
        RECT 677.220 1010.490 677.480 1010.810 ;
        RECT 677.280 999.330 677.420 1010.490 ;
        RECT 678.030 999.330 678.310 1000.000 ;
        RECT 677.280 999.190 678.310 999.330 ;
        RECT 678.030 996.000 678.310 999.190 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 210.290 3501.560 210.610 3501.620 ;
        RECT 40.550 3501.420 210.610 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 210.290 3501.360 210.610 3501.420 ;
        RECT 210.290 1019.900 210.610 1019.960 ;
        RECT 696.970 1019.900 697.290 1019.960 ;
        RECT 210.290 1019.760 697.290 1019.900 ;
        RECT 210.290 1019.700 210.610 1019.760 ;
        RECT 696.970 1019.700 697.290 1019.760 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 210.320 3501.360 210.580 3501.620 ;
        RECT 210.320 1019.700 210.580 1019.960 ;
        RECT 697.000 1019.700 697.260 1019.960 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.650 40.780 3517.600 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 210.320 3501.330 210.580 3501.650 ;
        RECT 210.380 1019.990 210.520 3501.330 ;
        RECT 210.320 1019.670 210.580 1019.990 ;
        RECT 697.000 1019.670 697.260 1019.990 ;
        RECT 697.060 999.330 697.200 1019.670 ;
        RECT 699.190 999.330 699.470 1000.000 ;
        RECT 697.060 999.190 699.470 999.330 ;
        RECT 699.190 996.000 699.470 999.190 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3284.640 17.410 3284.700 ;
        RECT 717.670 3284.640 717.990 3284.700 ;
        RECT 17.090 3284.500 717.990 3284.640 ;
        RECT 17.090 3284.440 17.410 3284.500 ;
        RECT 717.670 3284.440 717.990 3284.500 ;
      LAYER via ;
        RECT 17.120 3284.440 17.380 3284.700 ;
        RECT 717.700 3284.440 717.960 3284.700 ;
      LAYER met2 ;
        RECT 17.110 3290.675 17.390 3291.045 ;
        RECT 17.180 3284.730 17.320 3290.675 ;
        RECT 17.120 3284.410 17.380 3284.730 ;
        RECT 717.700 3284.410 717.960 3284.730 ;
        RECT 717.760 1048.870 717.900 3284.410 ;
        RECT 717.760 1048.730 718.360 1048.870 ;
        RECT 718.220 999.330 718.360 1048.730 ;
        RECT 720.350 999.330 720.630 1000.000 ;
        RECT 718.220 999.190 720.630 999.330 ;
        RECT 720.350 996.000 720.630 999.190 ;
      LAYER via2 ;
        RECT 17.110 3290.720 17.390 3291.000 ;
      LAYER met3 ;
        RECT -4.800 3291.010 2.400 3291.460 ;
        RECT 17.085 3291.010 17.415 3291.025 ;
        RECT -4.800 3290.710 17.415 3291.010 ;
        RECT -4.800 3290.260 2.400 3290.710 ;
        RECT 17.085 3290.695 17.415 3290.710 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 3029.300 16.490 3029.360 ;
        RECT 738.370 3029.300 738.690 3029.360 ;
        RECT 16.170 3029.160 738.690 3029.300 ;
        RECT 16.170 3029.100 16.490 3029.160 ;
        RECT 738.370 3029.100 738.690 3029.160 ;
      LAYER via ;
        RECT 16.200 3029.100 16.460 3029.360 ;
        RECT 738.400 3029.100 738.660 3029.360 ;
      LAYER met2 ;
        RECT 16.190 3030.235 16.470 3030.605 ;
        RECT 16.260 3029.390 16.400 3030.235 ;
        RECT 16.200 3029.070 16.460 3029.390 ;
        RECT 738.400 3029.070 738.660 3029.390 ;
        RECT 738.460 1048.870 738.600 3029.070 ;
        RECT 738.460 1048.730 740.440 1048.870 ;
        RECT 740.300 999.330 740.440 1048.730 ;
        RECT 741.970 999.330 742.250 1000.000 ;
        RECT 740.300 999.190 742.250 999.330 ;
        RECT 741.970 996.000 742.250 999.190 ;
      LAYER via2 ;
        RECT 16.190 3030.280 16.470 3030.560 ;
      LAYER met3 ;
        RECT -4.800 3030.570 2.400 3031.020 ;
        RECT 16.165 3030.570 16.495 3030.585 ;
        RECT -4.800 3030.270 16.495 3030.570 ;
        RECT -4.800 3029.820 2.400 3030.270 ;
        RECT 16.165 3030.255 16.495 3030.270 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2767.160 17.410 2767.220 ;
        RECT 759.070 2767.160 759.390 2767.220 ;
        RECT 17.090 2767.020 759.390 2767.160 ;
        RECT 17.090 2766.960 17.410 2767.020 ;
        RECT 759.070 2766.960 759.390 2767.020 ;
      LAYER via ;
        RECT 17.120 2766.960 17.380 2767.220 ;
        RECT 759.100 2766.960 759.360 2767.220 ;
      LAYER met2 ;
        RECT 17.110 2769.115 17.390 2769.485 ;
        RECT 17.180 2767.250 17.320 2769.115 ;
        RECT 17.120 2766.930 17.380 2767.250 ;
        RECT 759.100 2766.930 759.360 2767.250 ;
        RECT 759.160 1048.870 759.300 2766.930 ;
        RECT 759.160 1048.730 761.600 1048.870 ;
        RECT 761.460 999.330 761.600 1048.730 ;
        RECT 763.130 999.330 763.410 1000.000 ;
        RECT 761.460 999.190 763.410 999.330 ;
        RECT 763.130 996.000 763.410 999.190 ;
      LAYER via2 ;
        RECT 17.110 2769.160 17.390 2769.440 ;
      LAYER met3 ;
        RECT -4.800 2769.450 2.400 2769.900 ;
        RECT 17.085 2769.450 17.415 2769.465 ;
        RECT -4.800 2769.150 17.415 2769.450 ;
        RECT -4.800 2768.700 2.400 2769.150 ;
        RECT 17.085 2769.135 17.415 2769.150 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2505.020 15.570 2505.080 ;
        RECT 779.770 2505.020 780.090 2505.080 ;
        RECT 15.250 2504.880 780.090 2505.020 ;
        RECT 15.250 2504.820 15.570 2504.880 ;
        RECT 779.770 2504.820 780.090 2504.880 ;
      LAYER via ;
        RECT 15.280 2504.820 15.540 2505.080 ;
        RECT 779.800 2504.820 780.060 2505.080 ;
      LAYER met2 ;
        RECT 15.270 2508.675 15.550 2509.045 ;
        RECT 15.340 2505.110 15.480 2508.675 ;
        RECT 15.280 2504.790 15.540 2505.110 ;
        RECT 779.800 2504.790 780.060 2505.110 ;
        RECT 779.860 1048.870 780.000 2504.790 ;
        RECT 779.860 1048.730 782.760 1048.870 ;
        RECT 782.620 999.330 782.760 1048.730 ;
        RECT 784.290 999.330 784.570 1000.000 ;
        RECT 782.620 999.190 784.570 999.330 ;
        RECT 784.290 996.000 784.570 999.190 ;
      LAYER via2 ;
        RECT 15.270 2508.720 15.550 2509.000 ;
      LAYER met3 ;
        RECT -4.800 2509.010 2.400 2509.460 ;
        RECT 15.245 2509.010 15.575 2509.025 ;
        RECT -4.800 2508.710 15.575 2509.010 ;
        RECT -4.800 2508.260 2.400 2508.710 ;
        RECT 15.245 2508.695 15.575 2508.710 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2242.880 16.030 2242.940 ;
        RECT 800.470 2242.880 800.790 2242.940 ;
        RECT 15.710 2242.740 800.790 2242.880 ;
        RECT 15.710 2242.680 16.030 2242.740 ;
        RECT 800.470 2242.680 800.790 2242.740 ;
      LAYER via ;
        RECT 15.740 2242.680 16.000 2242.940 ;
        RECT 800.500 2242.680 800.760 2242.940 ;
      LAYER met2 ;
        RECT 15.730 2247.555 16.010 2247.925 ;
        RECT 15.800 2242.970 15.940 2247.555 ;
        RECT 15.740 2242.650 16.000 2242.970 ;
        RECT 800.500 2242.650 800.760 2242.970 ;
        RECT 800.560 1048.870 800.700 2242.650 ;
        RECT 800.560 1048.730 803.920 1048.870 ;
        RECT 803.780 999.330 803.920 1048.730 ;
        RECT 805.450 999.330 805.730 1000.000 ;
        RECT 803.780 999.190 805.730 999.330 ;
        RECT 805.450 996.000 805.730 999.190 ;
      LAYER via2 ;
        RECT 15.730 2247.600 16.010 2247.880 ;
      LAYER met3 ;
        RECT -4.800 2247.890 2.400 2248.340 ;
        RECT 15.705 2247.890 16.035 2247.905 ;
        RECT -4.800 2247.590 16.035 2247.890 ;
        RECT -4.800 2247.140 2.400 2247.590 ;
        RECT 15.705 2247.575 16.035 2247.590 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1987.540 17.410 1987.600 ;
        RECT 821.170 1987.540 821.490 1987.600 ;
        RECT 17.090 1987.400 821.490 1987.540 ;
        RECT 17.090 1987.340 17.410 1987.400 ;
        RECT 821.170 1987.340 821.490 1987.400 ;
      LAYER via ;
        RECT 17.120 1987.340 17.380 1987.600 ;
        RECT 821.200 1987.340 821.460 1987.600 ;
      LAYER met2 ;
        RECT 17.120 1987.485 17.380 1987.630 ;
        RECT 17.110 1987.115 17.390 1987.485 ;
        RECT 821.200 1987.310 821.460 1987.630 ;
        RECT 821.260 1048.870 821.400 1987.310 ;
        RECT 821.260 1048.730 825.080 1048.870 ;
        RECT 824.940 999.330 825.080 1048.730 ;
        RECT 827.070 999.330 827.350 1000.000 ;
        RECT 824.940 999.190 827.350 999.330 ;
        RECT 827.070 996.000 827.350 999.190 ;
      LAYER via2 ;
        RECT 17.110 1987.160 17.390 1987.440 ;
      LAYER met3 ;
        RECT -4.800 1987.450 2.400 1987.900 ;
        RECT 17.085 1987.450 17.415 1987.465 ;
        RECT -4.800 1987.150 17.415 1987.450 ;
        RECT -4.800 1986.700 2.400 1987.150 ;
        RECT 17.085 1987.135 17.415 1987.150 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 253.990 1002.220 254.310 1002.280 ;
        RECT 2900.370 1002.220 2900.690 1002.280 ;
        RECT 253.990 1002.080 2900.690 1002.220 ;
        RECT 253.990 1002.020 254.310 1002.080 ;
        RECT 2900.370 1002.020 2900.690 1002.080 ;
      LAYER via ;
        RECT 254.020 1002.020 254.280 1002.280 ;
        RECT 2900.400 1002.020 2900.660 1002.280 ;
      LAYER met2 ;
        RECT 254.020 1001.990 254.280 1002.310 ;
        RECT 2900.400 1001.990 2900.660 1002.310 ;
        RECT 252.530 999.330 252.810 1000.000 ;
        RECT 254.080 999.330 254.220 1001.990 ;
        RECT 252.530 999.190 254.220 999.330 ;
        RECT 252.530 996.000 252.810 999.190 ;
        RECT 2900.460 564.245 2900.600 1001.990 ;
        RECT 2900.390 563.875 2900.670 564.245 ;
      LAYER via2 ;
        RECT 2900.390 563.920 2900.670 564.200 ;
      LAYER met3 ;
        RECT 2900.365 564.210 2900.695 564.225 ;
        RECT 2917.600 564.210 2924.800 564.660 ;
        RECT 2900.365 563.910 2924.800 564.210 ;
        RECT 2900.365 563.895 2900.695 563.910 ;
        RECT 2917.600 563.460 2924.800 563.910 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1725.400 16.950 1725.460 ;
        RECT 841.870 1725.400 842.190 1725.460 ;
        RECT 16.630 1725.260 842.190 1725.400 ;
        RECT 16.630 1725.200 16.950 1725.260 ;
        RECT 841.870 1725.200 842.190 1725.260 ;
      LAYER via ;
        RECT 16.660 1725.200 16.920 1725.460 ;
        RECT 841.900 1725.200 842.160 1725.460 ;
      LAYER met2 ;
        RECT 16.650 1726.675 16.930 1727.045 ;
        RECT 16.720 1725.490 16.860 1726.675 ;
        RECT 16.660 1725.170 16.920 1725.490 ;
        RECT 841.900 1725.170 842.160 1725.490 ;
        RECT 841.960 1048.870 842.100 1725.170 ;
        RECT 841.960 1048.730 846.240 1048.870 ;
        RECT 846.100 999.330 846.240 1048.730 ;
        RECT 848.230 999.330 848.510 1000.000 ;
        RECT 846.100 999.190 848.510 999.330 ;
        RECT 848.230 996.000 848.510 999.190 ;
      LAYER via2 ;
        RECT 16.650 1726.720 16.930 1727.000 ;
      LAYER met3 ;
        RECT -4.800 1727.010 2.400 1727.460 ;
        RECT 16.625 1727.010 16.955 1727.025 ;
        RECT -4.800 1726.710 16.955 1727.010 ;
        RECT -4.800 1726.260 2.400 1726.710 ;
        RECT 16.625 1726.695 16.955 1726.710 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1462.920 17.870 1462.980 ;
        RECT 686.390 1462.920 686.710 1462.980 ;
        RECT 17.550 1462.780 686.710 1462.920 ;
        RECT 17.550 1462.720 17.870 1462.780 ;
        RECT 686.390 1462.720 686.710 1462.780 ;
        RECT 686.390 1011.060 686.710 1011.120 ;
        RECT 869.930 1011.060 870.250 1011.120 ;
        RECT 686.390 1010.920 870.250 1011.060 ;
        RECT 686.390 1010.860 686.710 1010.920 ;
        RECT 869.930 1010.860 870.250 1010.920 ;
      LAYER via ;
        RECT 17.580 1462.720 17.840 1462.980 ;
        RECT 686.420 1462.720 686.680 1462.980 ;
        RECT 686.420 1010.860 686.680 1011.120 ;
        RECT 869.960 1010.860 870.220 1011.120 ;
      LAYER met2 ;
        RECT 17.570 1465.555 17.850 1465.925 ;
        RECT 17.640 1463.010 17.780 1465.555 ;
        RECT 17.580 1462.690 17.840 1463.010 ;
        RECT 686.420 1462.690 686.680 1463.010 ;
        RECT 686.480 1011.150 686.620 1462.690 ;
        RECT 686.420 1010.830 686.680 1011.150 ;
        RECT 869.960 1010.830 870.220 1011.150 ;
        RECT 869.390 999.330 869.670 1000.000 ;
        RECT 870.020 999.330 870.160 1010.830 ;
        RECT 869.390 999.190 870.160 999.330 ;
        RECT 869.390 996.000 869.670 999.190 ;
      LAYER via2 ;
        RECT 17.570 1465.600 17.850 1465.880 ;
      LAYER met3 ;
        RECT -4.800 1465.890 2.400 1466.340 ;
        RECT 17.545 1465.890 17.875 1465.905 ;
        RECT -4.800 1465.590 17.875 1465.890 ;
        RECT -4.800 1465.140 2.400 1465.590 ;
        RECT 17.545 1465.575 17.875 1465.590 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1200.780 15.570 1200.840 ;
        RECT 686.850 1200.780 687.170 1200.840 ;
        RECT 15.250 1200.640 687.170 1200.780 ;
        RECT 15.250 1200.580 15.570 1200.640 ;
        RECT 686.850 1200.580 687.170 1200.640 ;
        RECT 686.850 1010.720 687.170 1010.780 ;
        RECT 890.170 1010.720 890.490 1010.780 ;
        RECT 686.850 1010.580 890.490 1010.720 ;
        RECT 686.850 1010.520 687.170 1010.580 ;
        RECT 890.170 1010.520 890.490 1010.580 ;
      LAYER via ;
        RECT 15.280 1200.580 15.540 1200.840 ;
        RECT 686.880 1200.580 687.140 1200.840 ;
        RECT 686.880 1010.520 687.140 1010.780 ;
        RECT 890.200 1010.520 890.460 1010.780 ;
      LAYER met2 ;
        RECT 15.270 1205.115 15.550 1205.485 ;
        RECT 15.340 1200.870 15.480 1205.115 ;
        RECT 15.280 1200.550 15.540 1200.870 ;
        RECT 686.880 1200.550 687.140 1200.870 ;
        RECT 686.940 1010.810 687.080 1200.550 ;
        RECT 686.880 1010.490 687.140 1010.810 ;
        RECT 890.200 1010.490 890.460 1010.810 ;
        RECT 890.260 999.330 890.400 1010.490 ;
        RECT 890.550 999.330 890.830 1000.000 ;
        RECT 890.260 999.190 890.830 999.330 ;
        RECT 890.550 996.000 890.830 999.190 ;
      LAYER via2 ;
        RECT 15.270 1205.160 15.550 1205.440 ;
      LAYER met3 ;
        RECT -4.800 1205.450 2.400 1205.900 ;
        RECT 15.245 1205.450 15.575 1205.465 ;
        RECT -4.800 1205.150 15.575 1205.450 ;
        RECT -4.800 1204.700 2.400 1205.150 ;
        RECT 15.245 1205.135 15.575 1205.150 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1004.600 15.570 1004.660 ;
        RECT 910.870 1004.600 911.190 1004.660 ;
        RECT 15.250 1004.460 911.190 1004.600 ;
        RECT 15.250 1004.400 15.570 1004.460 ;
        RECT 910.870 1004.400 911.190 1004.460 ;
      LAYER via ;
        RECT 15.280 1004.400 15.540 1004.660 ;
        RECT 910.900 1004.400 911.160 1004.660 ;
      LAYER met2 ;
        RECT 15.280 1004.370 15.540 1004.690 ;
        RECT 910.900 1004.370 911.160 1004.690 ;
        RECT 15.340 944.365 15.480 1004.370 ;
        RECT 910.960 999.330 911.100 1004.370 ;
        RECT 911.710 999.330 911.990 1000.000 ;
        RECT 910.960 999.190 911.990 999.330 ;
        RECT 911.710 996.000 911.990 999.190 ;
        RECT 15.270 943.995 15.550 944.365 ;
      LAYER via2 ;
        RECT 15.270 944.040 15.550 944.320 ;
      LAYER met3 ;
        RECT -4.800 944.330 2.400 944.780 ;
        RECT 15.245 944.330 15.575 944.345 ;
        RECT -4.800 944.030 15.575 944.330 ;
        RECT -4.800 943.580 2.400 944.030 ;
        RECT 15.245 944.015 15.575 944.030 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1003.920 16.950 1003.980 ;
        RECT 932.030 1003.920 932.350 1003.980 ;
        RECT 16.630 1003.780 932.350 1003.920 ;
        RECT 16.630 1003.720 16.950 1003.780 ;
        RECT 932.030 1003.720 932.350 1003.780 ;
      LAYER via ;
        RECT 16.660 1003.720 16.920 1003.980 ;
        RECT 932.060 1003.720 932.320 1003.980 ;
      LAYER met2 ;
        RECT 16.660 1003.690 16.920 1004.010 ;
        RECT 932.060 1003.690 932.320 1004.010 ;
        RECT 16.720 683.925 16.860 1003.690 ;
        RECT 932.120 999.330 932.260 1003.690 ;
        RECT 933.330 999.330 933.610 1000.000 ;
        RECT 932.120 999.190 933.610 999.330 ;
        RECT 933.330 996.000 933.610 999.190 ;
        RECT 16.650 683.555 16.930 683.925 ;
      LAYER via2 ;
        RECT 16.650 683.600 16.930 683.880 ;
      LAYER met3 ;
        RECT -4.800 683.890 2.400 684.340 ;
        RECT 16.625 683.890 16.955 683.905 ;
        RECT -4.800 683.590 16.955 683.890 ;
        RECT -4.800 683.140 2.400 683.590 ;
        RECT 16.625 683.575 16.955 683.590 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 1003.580 19.250 1003.640 ;
        RECT 953.190 1003.580 953.510 1003.640 ;
        RECT 18.930 1003.440 953.510 1003.580 ;
        RECT 18.930 1003.380 19.250 1003.440 ;
        RECT 953.190 1003.380 953.510 1003.440 ;
      LAYER via ;
        RECT 18.960 1003.380 19.220 1003.640 ;
        RECT 953.220 1003.380 953.480 1003.640 ;
      LAYER met2 ;
        RECT 18.960 1003.350 19.220 1003.670 ;
        RECT 953.220 1003.350 953.480 1003.670 ;
        RECT 19.020 423.485 19.160 1003.350 ;
        RECT 953.280 999.330 953.420 1003.350 ;
        RECT 954.490 999.330 954.770 1000.000 ;
        RECT 953.280 999.190 954.770 999.330 ;
        RECT 954.490 996.000 954.770 999.190 ;
        RECT 18.950 423.115 19.230 423.485 ;
      LAYER via2 ;
        RECT 18.950 423.160 19.230 423.440 ;
      LAYER met3 ;
        RECT -4.800 423.450 2.400 423.900 ;
        RECT 18.925 423.450 19.255 423.465 ;
        RECT -4.800 423.150 19.255 423.450 ;
        RECT -4.800 422.700 2.400 423.150 ;
        RECT 18.925 423.135 19.255 423.150 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1002.900 17.870 1002.960 ;
        RECT 974.350 1002.900 974.670 1002.960 ;
        RECT 17.550 1002.760 974.670 1002.900 ;
        RECT 17.550 1002.700 17.870 1002.760 ;
        RECT 974.350 1002.700 974.670 1002.760 ;
      LAYER via ;
        RECT 17.580 1002.700 17.840 1002.960 ;
        RECT 974.380 1002.700 974.640 1002.960 ;
      LAYER met2 ;
        RECT 17.580 1002.670 17.840 1002.990 ;
        RECT 974.380 1002.670 974.640 1002.990 ;
        RECT 17.640 227.645 17.780 1002.670 ;
        RECT 974.440 999.330 974.580 1002.670 ;
        RECT 975.650 999.330 975.930 1000.000 ;
        RECT 974.440 999.190 975.930 999.330 ;
        RECT 975.650 996.000 975.930 999.190 ;
        RECT 17.570 227.275 17.850 227.645 ;
      LAYER via2 ;
        RECT 17.570 227.320 17.850 227.600 ;
      LAYER met3 ;
        RECT -4.800 227.610 2.400 228.060 ;
        RECT 17.545 227.610 17.875 227.625 ;
        RECT -4.800 227.310 17.875 227.610 ;
        RECT -4.800 226.860 2.400 227.310 ;
        RECT 17.545 227.295 17.875 227.310 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23.990 1002.560 24.310 1002.620 ;
        RECT 995.510 1002.560 995.830 1002.620 ;
        RECT 23.990 1002.420 995.830 1002.560 ;
        RECT 23.990 1002.360 24.310 1002.420 ;
        RECT 995.510 1002.360 995.830 1002.420 ;
        RECT 13.870 32.540 14.190 32.600 ;
        RECT 23.990 32.540 24.310 32.600 ;
        RECT 13.870 32.400 24.310 32.540 ;
        RECT 13.870 32.340 14.190 32.400 ;
        RECT 23.990 32.340 24.310 32.400 ;
      LAYER via ;
        RECT 24.020 1002.360 24.280 1002.620 ;
        RECT 995.540 1002.360 995.800 1002.620 ;
        RECT 13.900 32.340 14.160 32.600 ;
        RECT 24.020 32.340 24.280 32.600 ;
      LAYER met2 ;
        RECT 24.020 1002.330 24.280 1002.650 ;
        RECT 995.540 1002.330 995.800 1002.650 ;
        RECT 24.080 32.630 24.220 1002.330 ;
        RECT 995.600 999.330 995.740 1002.330 ;
        RECT 996.810 999.330 997.090 1000.000 ;
        RECT 995.600 999.190 997.090 999.330 ;
        RECT 996.810 996.000 997.090 999.190 ;
        RECT 13.900 32.485 14.160 32.630 ;
        RECT 13.890 32.115 14.170 32.485 ;
        RECT 24.020 32.310 24.280 32.630 ;
      LAYER via2 ;
        RECT 13.890 32.160 14.170 32.440 ;
      LAYER met3 ;
        RECT -4.800 32.450 2.400 32.900 ;
        RECT 13.865 32.450 14.195 32.465 ;
        RECT -4.800 32.150 14.195 32.450 ;
        RECT -4.800 31.700 2.400 32.150 ;
        RECT 13.865 32.135 14.195 32.150 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 275.610 1009.700 275.930 1009.760 ;
        RECT 1101.770 1009.700 1102.090 1009.760 ;
        RECT 275.610 1009.560 1102.090 1009.700 ;
        RECT 275.610 1009.500 275.930 1009.560 ;
        RECT 1101.770 1009.500 1102.090 1009.560 ;
        RECT 1101.770 765.920 1102.090 765.980 ;
        RECT 2899.910 765.920 2900.230 765.980 ;
        RECT 1101.770 765.780 2900.230 765.920 ;
        RECT 1101.770 765.720 1102.090 765.780 ;
        RECT 2899.910 765.720 2900.230 765.780 ;
      LAYER via ;
        RECT 275.640 1009.500 275.900 1009.760 ;
        RECT 1101.800 1009.500 1102.060 1009.760 ;
        RECT 1101.800 765.720 1102.060 765.980 ;
        RECT 2899.940 765.720 2900.200 765.980 ;
      LAYER met2 ;
        RECT 275.640 1009.470 275.900 1009.790 ;
        RECT 1101.800 1009.470 1102.060 1009.790 ;
        RECT 274.150 999.330 274.430 1000.000 ;
        RECT 275.700 999.330 275.840 1009.470 ;
        RECT 274.150 999.190 275.840 999.330 ;
        RECT 274.150 996.000 274.430 999.190 ;
        RECT 1101.860 766.010 1102.000 1009.470 ;
        RECT 1101.800 765.690 1102.060 766.010 ;
        RECT 2899.940 765.690 2900.200 766.010 ;
        RECT 2900.000 763.485 2900.140 765.690 ;
        RECT 2899.930 763.115 2900.210 763.485 ;
      LAYER via2 ;
        RECT 2899.930 763.160 2900.210 763.440 ;
      LAYER met3 ;
        RECT 2899.905 763.450 2900.235 763.465 ;
        RECT 2917.600 763.450 2924.800 763.900 ;
        RECT 2899.905 763.150 2924.800 763.450 ;
        RECT 2899.905 763.135 2900.235 763.150 ;
        RECT 2917.600 762.700 2924.800 763.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.310 1011.400 296.630 1011.460 ;
        RECT 1103.150 1011.400 1103.470 1011.460 ;
        RECT 296.310 1011.260 1103.470 1011.400 ;
        RECT 296.310 1011.200 296.630 1011.260 ;
        RECT 1103.150 1011.200 1103.470 1011.260 ;
        RECT 1103.150 965.840 1103.470 965.900 ;
        RECT 2899.910 965.840 2900.230 965.900 ;
        RECT 1103.150 965.700 2900.230 965.840 ;
        RECT 1103.150 965.640 1103.470 965.700 ;
        RECT 2899.910 965.640 2900.230 965.700 ;
      LAYER via ;
        RECT 296.340 1011.200 296.600 1011.460 ;
        RECT 1103.180 1011.200 1103.440 1011.460 ;
        RECT 1103.180 965.640 1103.440 965.900 ;
        RECT 2899.940 965.640 2900.200 965.900 ;
      LAYER met2 ;
        RECT 296.340 1011.170 296.600 1011.490 ;
        RECT 1103.180 1011.170 1103.440 1011.490 ;
        RECT 295.310 999.330 295.590 1000.000 ;
        RECT 296.400 999.330 296.540 1011.170 ;
        RECT 295.310 999.190 296.540 999.330 ;
        RECT 295.310 996.000 295.590 999.190 ;
        RECT 1103.240 965.930 1103.380 1011.170 ;
        RECT 1103.180 965.610 1103.440 965.930 ;
        RECT 2899.940 965.610 2900.200 965.930 ;
        RECT 2900.000 962.725 2900.140 965.610 ;
        RECT 2899.930 962.355 2900.210 962.725 ;
      LAYER via2 ;
        RECT 2899.930 962.400 2900.210 962.680 ;
      LAYER met3 ;
        RECT 2899.905 962.690 2900.235 962.705 ;
        RECT 2917.600 962.690 2924.800 963.140 ;
        RECT 2899.905 962.390 2924.800 962.690 ;
        RECT 2899.905 962.375 2900.235 962.390 ;
        RECT 2917.600 961.940 2924.800 962.390 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.570 1159.300 310.890 1159.360 ;
        RECT 2900.830 1159.300 2901.150 1159.360 ;
        RECT 310.570 1159.160 2901.150 1159.300 ;
        RECT 310.570 1159.100 310.890 1159.160 ;
        RECT 2900.830 1159.100 2901.150 1159.160 ;
      LAYER via ;
        RECT 310.600 1159.100 310.860 1159.360 ;
        RECT 2900.860 1159.100 2901.120 1159.360 ;
      LAYER met2 ;
        RECT 2900.850 1161.595 2901.130 1161.965 ;
        RECT 2900.920 1159.390 2901.060 1161.595 ;
        RECT 310.600 1159.070 310.860 1159.390 ;
        RECT 2900.860 1159.070 2901.120 1159.390 ;
        RECT 310.660 1048.870 310.800 1159.070 ;
        RECT 310.660 1048.730 314.480 1048.870 ;
        RECT 314.340 999.330 314.480 1048.730 ;
        RECT 316.470 999.330 316.750 1000.000 ;
        RECT 314.340 999.190 316.750 999.330 ;
        RECT 316.470 996.000 316.750 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1161.640 2901.130 1161.920 ;
      LAYER met3 ;
        RECT 2900.825 1161.930 2901.155 1161.945 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2900.825 1161.630 2924.800 1161.930 ;
        RECT 2900.825 1161.615 2901.155 1161.630 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 1359.560 331.590 1359.620 ;
        RECT 2900.830 1359.560 2901.150 1359.620 ;
        RECT 331.270 1359.420 2901.150 1359.560 ;
        RECT 331.270 1359.360 331.590 1359.420 ;
        RECT 2900.830 1359.360 2901.150 1359.420 ;
      LAYER via ;
        RECT 331.300 1359.360 331.560 1359.620 ;
        RECT 2900.860 1359.360 2901.120 1359.620 ;
      LAYER met2 ;
        RECT 2900.850 1360.835 2901.130 1361.205 ;
        RECT 2900.920 1359.650 2901.060 1360.835 ;
        RECT 331.300 1359.330 331.560 1359.650 ;
        RECT 2900.860 1359.330 2901.120 1359.650 ;
        RECT 331.360 1048.870 331.500 1359.330 ;
        RECT 331.360 1048.730 335.640 1048.870 ;
        RECT 335.500 999.330 335.640 1048.730 ;
        RECT 337.630 999.330 337.910 1000.000 ;
        RECT 335.500 999.190 337.910 999.330 ;
        RECT 337.630 996.000 337.910 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1360.880 2901.130 1361.160 ;
      LAYER met3 ;
        RECT 2900.825 1361.170 2901.155 1361.185 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2900.825 1360.870 2924.800 1361.170 ;
        RECT 2900.825 1360.855 2901.155 1360.870 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.330 1621.700 359.650 1621.760 ;
        RECT 2898.070 1621.700 2898.390 1621.760 ;
        RECT 359.330 1621.560 2898.390 1621.700 ;
        RECT 359.330 1621.500 359.650 1621.560 ;
        RECT 2898.070 1621.500 2898.390 1621.560 ;
      LAYER via ;
        RECT 359.360 1621.500 359.620 1621.760 ;
        RECT 2898.100 1621.500 2898.360 1621.760 ;
      LAYER met2 ;
        RECT 2898.090 1626.035 2898.370 1626.405 ;
        RECT 2898.160 1621.790 2898.300 1626.035 ;
        RECT 359.360 1621.470 359.620 1621.790 ;
        RECT 2898.100 1621.470 2898.360 1621.790 ;
        RECT 359.420 1048.870 359.560 1621.470 ;
        RECT 359.420 1048.730 360.020 1048.870 ;
        RECT 359.250 999.330 359.530 1000.000 ;
        RECT 359.880 999.330 360.020 1048.730 ;
        RECT 359.250 999.190 360.020 999.330 ;
        RECT 359.250 996.000 359.530 999.190 ;
      LAYER via2 ;
        RECT 2898.090 1626.080 2898.370 1626.360 ;
      LAYER met3 ;
        RECT 2898.065 1626.370 2898.395 1626.385 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2898.065 1626.070 2924.800 1626.370 ;
        RECT 2898.065 1626.055 2898.395 1626.070 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.570 1890.980 379.890 1891.040 ;
        RECT 2900.830 1890.980 2901.150 1891.040 ;
        RECT 379.570 1890.840 2901.150 1890.980 ;
        RECT 379.570 1890.780 379.890 1890.840 ;
        RECT 2900.830 1890.780 2901.150 1890.840 ;
      LAYER via ;
        RECT 379.600 1890.780 379.860 1891.040 ;
        RECT 2900.860 1890.780 2901.120 1891.040 ;
      LAYER met2 ;
        RECT 2900.850 1891.915 2901.130 1892.285 ;
        RECT 2900.920 1891.070 2901.060 1891.915 ;
        RECT 379.600 1890.750 379.860 1891.070 ;
        RECT 2900.860 1890.750 2901.120 1891.070 ;
        RECT 379.660 999.330 379.800 1890.750 ;
        RECT 380.410 999.330 380.690 1000.000 ;
        RECT 379.660 999.190 380.690 999.330 ;
        RECT 380.410 996.000 380.690 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1891.960 2901.130 1892.240 ;
      LAYER met3 ;
        RECT 2900.825 1892.250 2901.155 1892.265 ;
        RECT 2917.600 1892.250 2924.800 1892.700 ;
        RECT 2900.825 1891.950 2924.800 1892.250 ;
        RECT 2900.825 1891.935 2901.155 1891.950 ;
        RECT 2917.600 1891.500 2924.800 1891.950 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 2153.120 400.590 2153.180 ;
        RECT 2900.830 2153.120 2901.150 2153.180 ;
        RECT 400.270 2152.980 2901.150 2153.120 ;
        RECT 400.270 2152.920 400.590 2152.980 ;
        RECT 2900.830 2152.920 2901.150 2152.980 ;
      LAYER via ;
        RECT 400.300 2152.920 400.560 2153.180 ;
        RECT 2900.860 2152.920 2901.120 2153.180 ;
      LAYER met2 ;
        RECT 2900.850 2157.795 2901.130 2158.165 ;
        RECT 2900.920 2153.210 2901.060 2157.795 ;
        RECT 400.300 2152.890 400.560 2153.210 ;
        RECT 2900.860 2152.890 2901.120 2153.210 ;
        RECT 400.360 999.330 400.500 2152.890 ;
        RECT 401.570 999.330 401.850 1000.000 ;
        RECT 400.360 999.190 401.850 999.330 ;
        RECT 401.570 996.000 401.850 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2157.840 2901.130 2158.120 ;
      LAYER met3 ;
        RECT 2900.825 2158.130 2901.155 2158.145 ;
        RECT 2917.600 2158.130 2924.800 2158.580 ;
        RECT 2900.825 2157.830 2924.800 2158.130 ;
        RECT 2900.825 2157.815 2901.155 2157.830 ;
        RECT 2917.600 2157.380 2924.800 2157.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 218.570 997.260 218.890 997.520 ;
        RECT 218.660 994.060 218.800 997.260 ;
        RECT 2902.670 994.060 2902.990 994.120 ;
        RECT 218.660 993.920 2902.990 994.060 ;
        RECT 2902.670 993.860 2902.990 993.920 ;
      LAYER via ;
        RECT 218.600 997.260 218.860 997.520 ;
        RECT 2902.700 993.860 2902.960 994.120 ;
      LAYER met2 ;
        RECT 217.110 997.290 217.390 1000.000 ;
        RECT 218.600 997.290 218.860 997.550 ;
        RECT 217.110 997.230 218.860 997.290 ;
        RECT 217.110 997.150 218.800 997.230 ;
        RECT 217.110 996.000 217.390 997.150 ;
        RECT 2902.700 993.830 2902.960 994.150 ;
        RECT 2902.760 99.125 2902.900 993.830 ;
        RECT 2902.690 98.755 2902.970 99.125 ;
      LAYER via2 ;
        RECT 2902.690 98.800 2902.970 99.080 ;
      LAYER met3 ;
        RECT 2902.665 99.090 2902.995 99.105 ;
        RECT 2917.600 99.090 2924.800 99.540 ;
        RECT 2902.665 98.790 2924.800 99.090 ;
        RECT 2902.665 98.775 2902.995 98.790 ;
        RECT 2917.600 98.340 2924.800 98.790 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 2353.040 428.190 2353.100 ;
        RECT 2900.830 2353.040 2901.150 2353.100 ;
        RECT 427.870 2352.900 2901.150 2353.040 ;
        RECT 427.870 2352.840 428.190 2352.900 ;
        RECT 2900.830 2352.840 2901.150 2352.900 ;
      LAYER via ;
        RECT 427.900 2352.840 428.160 2353.100 ;
        RECT 2900.860 2352.840 2901.120 2353.100 ;
      LAYER met2 ;
        RECT 2900.850 2357.035 2901.130 2357.405 ;
        RECT 2900.920 2353.130 2901.060 2357.035 ;
        RECT 427.900 2352.810 428.160 2353.130 ;
        RECT 2900.860 2352.810 2901.120 2353.130 ;
        RECT 427.960 1048.870 428.100 2352.810 ;
        RECT 427.960 1048.730 428.560 1048.870 ;
        RECT 428.420 999.330 428.560 1048.730 ;
        RECT 430.090 999.330 430.370 1000.000 ;
        RECT 428.420 999.190 430.370 999.330 ;
        RECT 430.090 996.000 430.370 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2357.080 2901.130 2357.360 ;
      LAYER met3 ;
        RECT 2900.825 2357.370 2901.155 2357.385 ;
        RECT 2917.600 2357.370 2924.800 2357.820 ;
        RECT 2900.825 2357.070 2924.800 2357.370 ;
        RECT 2900.825 2357.055 2901.155 2357.070 ;
        RECT 2917.600 2356.620 2924.800 2357.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 2622.320 448.890 2622.380 ;
        RECT 2900.830 2622.320 2901.150 2622.380 ;
        RECT 448.570 2622.180 2901.150 2622.320 ;
        RECT 448.570 2622.120 448.890 2622.180 ;
        RECT 2900.830 2622.120 2901.150 2622.180 ;
      LAYER via ;
        RECT 448.600 2622.120 448.860 2622.380 ;
        RECT 2900.860 2622.120 2901.120 2622.380 ;
      LAYER met2 ;
        RECT 448.600 2622.090 448.860 2622.410 ;
        RECT 2900.850 2622.235 2901.130 2622.605 ;
        RECT 2900.860 2622.090 2901.120 2622.235 ;
        RECT 448.660 1048.870 448.800 2622.090 ;
        RECT 448.660 1048.730 449.720 1048.870 ;
        RECT 449.580 999.330 449.720 1048.730 ;
        RECT 451.250 999.330 451.530 1000.000 ;
        RECT 449.580 999.190 451.530 999.330 ;
        RECT 451.250 996.000 451.530 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2622.280 2901.130 2622.560 ;
      LAYER met3 ;
        RECT 2900.825 2622.570 2901.155 2622.585 ;
        RECT 2917.600 2622.570 2924.800 2623.020 ;
        RECT 2900.825 2622.270 2924.800 2622.570 ;
        RECT 2900.825 2622.255 2901.155 2622.270 ;
        RECT 2917.600 2621.820 2924.800 2622.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 2884.460 469.590 2884.520 ;
        RECT 2900.830 2884.460 2901.150 2884.520 ;
        RECT 469.270 2884.320 2901.150 2884.460 ;
        RECT 469.270 2884.260 469.590 2884.320 ;
        RECT 2900.830 2884.260 2901.150 2884.320 ;
      LAYER via ;
        RECT 469.300 2884.260 469.560 2884.520 ;
        RECT 2900.860 2884.260 2901.120 2884.520 ;
      LAYER met2 ;
        RECT 2900.850 2888.115 2901.130 2888.485 ;
        RECT 2900.920 2884.550 2901.060 2888.115 ;
        RECT 469.300 2884.230 469.560 2884.550 ;
        RECT 2900.860 2884.230 2901.120 2884.550 ;
        RECT 469.360 1048.870 469.500 2884.230 ;
        RECT 469.360 1048.730 470.880 1048.870 ;
        RECT 470.740 999.330 470.880 1048.730 ;
        RECT 472.410 999.330 472.690 1000.000 ;
        RECT 470.740 999.190 472.690 999.330 ;
        RECT 472.410 996.000 472.690 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2888.160 2901.130 2888.440 ;
      LAYER met3 ;
        RECT 2900.825 2888.450 2901.155 2888.465 ;
        RECT 2917.600 2888.450 2924.800 2888.900 ;
        RECT 2900.825 2888.150 2924.800 2888.450 ;
        RECT 2900.825 2888.135 2901.155 2888.150 ;
        RECT 2917.600 2887.700 2924.800 2888.150 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 3153.400 490.290 3153.460 ;
        RECT 2899.910 3153.400 2900.230 3153.460 ;
        RECT 489.970 3153.260 2900.230 3153.400 ;
        RECT 489.970 3153.200 490.290 3153.260 ;
        RECT 2899.910 3153.200 2900.230 3153.260 ;
      LAYER via ;
        RECT 490.000 3153.200 490.260 3153.460 ;
        RECT 2899.940 3153.200 2900.200 3153.460 ;
      LAYER met2 ;
        RECT 2899.930 3153.995 2900.210 3154.365 ;
        RECT 2900.000 3153.490 2900.140 3153.995 ;
        RECT 490.000 3153.170 490.260 3153.490 ;
        RECT 2899.940 3153.170 2900.200 3153.490 ;
        RECT 490.060 1048.870 490.200 3153.170 ;
        RECT 490.060 1048.730 492.040 1048.870 ;
        RECT 491.900 999.330 492.040 1048.730 ;
        RECT 493.570 999.330 493.850 1000.000 ;
        RECT 491.900 999.190 493.850 999.330 ;
        RECT 493.570 996.000 493.850 999.190 ;
      LAYER via2 ;
        RECT 2899.930 3154.040 2900.210 3154.320 ;
      LAYER met3 ;
        RECT 2899.905 3154.330 2900.235 3154.345 ;
        RECT 2917.600 3154.330 2924.800 3154.780 ;
        RECT 2899.905 3154.030 2924.800 3154.330 ;
        RECT 2899.905 3154.015 2900.235 3154.030 ;
        RECT 2917.600 3153.580 2924.800 3154.030 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 3415.880 510.990 3415.940 ;
        RECT 2900.830 3415.880 2901.150 3415.940 ;
        RECT 510.670 3415.740 2901.150 3415.880 ;
        RECT 510.670 3415.680 510.990 3415.740 ;
        RECT 2900.830 3415.680 2901.150 3415.740 ;
      LAYER via ;
        RECT 510.700 3415.680 510.960 3415.940 ;
        RECT 2900.860 3415.680 2901.120 3415.940 ;
      LAYER met2 ;
        RECT 2900.850 3419.195 2901.130 3419.565 ;
        RECT 2900.920 3415.970 2901.060 3419.195 ;
        RECT 510.700 3415.650 510.960 3415.970 ;
        RECT 2900.860 3415.650 2901.120 3415.970 ;
        RECT 510.760 1048.870 510.900 3415.650 ;
        RECT 510.760 1048.730 513.200 1048.870 ;
        RECT 513.060 999.330 513.200 1048.730 ;
        RECT 515.190 999.330 515.470 1000.000 ;
        RECT 513.060 999.190 515.470 999.330 ;
        RECT 515.190 996.000 515.470 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3419.240 2901.130 3419.520 ;
      LAYER met3 ;
        RECT 2900.825 3419.530 2901.155 3419.545 ;
        RECT 2917.600 3419.530 2924.800 3419.980 ;
        RECT 2900.825 3419.230 2924.800 3419.530 ;
        RECT 2900.825 3419.215 2901.155 3419.230 ;
        RECT 2917.600 3418.780 2924.800 3419.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 3501.560 531.690 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 531.370 3501.420 2717.610 3501.560 ;
        RECT 531.370 3501.360 531.690 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
      LAYER via ;
        RECT 531.400 3501.360 531.660 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 531.400 3501.330 531.660 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 531.460 1048.870 531.600 3501.330 ;
        RECT 531.460 1048.730 534.360 1048.870 ;
        RECT 534.220 999.330 534.360 1048.730 ;
        RECT 536.350 999.330 536.630 1000.000 ;
        RECT 534.220 999.190 536.630 999.330 ;
        RECT 536.350 996.000 536.630 999.190 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 3502.240 552.390 3502.300 ;
        RECT 2392.530 3502.240 2392.850 3502.300 ;
        RECT 552.070 3502.100 2392.850 3502.240 ;
        RECT 552.070 3502.040 552.390 3502.100 ;
        RECT 2392.530 3502.040 2392.850 3502.100 ;
      LAYER via ;
        RECT 552.100 3502.040 552.360 3502.300 ;
        RECT 2392.560 3502.040 2392.820 3502.300 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.330 2392.760 3517.600 ;
        RECT 552.100 3502.010 552.360 3502.330 ;
        RECT 2392.560 3502.010 2392.820 3502.330 ;
        RECT 552.160 1048.870 552.300 3502.010 ;
        RECT 552.160 1048.730 555.520 1048.870 ;
        RECT 555.380 999.330 555.520 1048.730 ;
        RECT 557.510 999.330 557.790 1000.000 ;
        RECT 555.380 999.190 557.790 999.330 ;
        RECT 557.510 996.000 557.790 999.190 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 3502.920 573.090 3502.980 ;
        RECT 2068.230 3502.920 2068.550 3502.980 ;
        RECT 572.770 3502.780 2068.550 3502.920 ;
        RECT 572.770 3502.720 573.090 3502.780 ;
        RECT 2068.230 3502.720 2068.550 3502.780 ;
      LAYER via ;
        RECT 572.800 3502.720 573.060 3502.980 ;
        RECT 2068.260 3502.720 2068.520 3502.980 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3503.010 2068.460 3517.600 ;
        RECT 572.800 3502.690 573.060 3503.010 ;
        RECT 2068.260 3502.690 2068.520 3503.010 ;
        RECT 572.860 1048.870 573.000 3502.690 ;
        RECT 572.860 1048.730 576.680 1048.870 ;
        RECT 576.540 999.330 576.680 1048.730 ;
        RECT 578.670 999.330 578.950 1000.000 ;
        RECT 576.540 999.190 578.950 999.330 ;
        RECT 578.670 996.000 578.950 999.190 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 3503.600 593.790 3503.660 ;
        RECT 1743.930 3503.600 1744.250 3503.660 ;
        RECT 593.470 3503.460 1744.250 3503.600 ;
        RECT 593.470 3503.400 593.790 3503.460 ;
        RECT 1743.930 3503.400 1744.250 3503.460 ;
      LAYER via ;
        RECT 593.500 3503.400 593.760 3503.660 ;
        RECT 1743.960 3503.400 1744.220 3503.660 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.690 1744.160 3517.600 ;
        RECT 593.500 3503.370 593.760 3503.690 ;
        RECT 1743.960 3503.370 1744.220 3503.690 ;
        RECT 593.560 1048.870 593.700 3503.370 ;
        RECT 593.560 1048.730 597.840 1048.870 ;
        RECT 597.700 999.330 597.840 1048.730 ;
        RECT 599.830 999.330 600.110 1000.000 ;
        RECT 597.700 999.190 600.110 999.330 ;
        RECT 599.830 996.000 600.110 999.190 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 3504.280 621.390 3504.340 ;
        RECT 1419.170 3504.280 1419.490 3504.340 ;
        RECT 621.070 3504.140 1419.490 3504.280 ;
        RECT 621.070 3504.080 621.390 3504.140 ;
        RECT 1419.170 3504.080 1419.490 3504.140 ;
      LAYER via ;
        RECT 621.100 3504.080 621.360 3504.340 ;
        RECT 1419.200 3504.080 1419.460 3504.340 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3504.370 1419.400 3517.600 ;
        RECT 621.100 3504.050 621.360 3504.370 ;
        RECT 1419.200 3504.050 1419.460 3504.370 ;
        RECT 621.160 999.330 621.300 3504.050 ;
        RECT 621.450 999.330 621.730 1000.000 ;
        RECT 621.160 999.190 621.730 999.330 ;
        RECT 621.450 996.000 621.730 999.190 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 240.650 997.460 240.970 997.520 ;
        RECT 240.650 997.320 253.300 997.460 ;
        RECT 240.650 997.260 240.970 997.320 ;
        RECT 253.160 994.400 253.300 997.320 ;
        RECT 2904.050 994.400 2904.370 994.460 ;
        RECT 253.160 994.260 2904.370 994.400 ;
        RECT 2904.050 994.200 2904.370 994.260 ;
      LAYER via ;
        RECT 240.680 997.260 240.940 997.520 ;
        RECT 2904.080 994.200 2904.340 994.460 ;
      LAYER met2 ;
        RECT 238.730 997.290 239.010 1000.000 ;
        RECT 240.680 997.290 240.940 997.550 ;
        RECT 238.730 997.230 240.940 997.290 ;
        RECT 238.730 997.150 240.880 997.230 ;
        RECT 238.730 996.000 239.010 997.150 ;
        RECT 2904.080 994.170 2904.340 994.490 ;
        RECT 2904.140 298.365 2904.280 994.170 ;
        RECT 2904.070 297.995 2904.350 298.365 ;
      LAYER via2 ;
        RECT 2904.070 298.040 2904.350 298.320 ;
      LAYER met3 ;
        RECT 2904.045 298.330 2904.375 298.345 ;
        RECT 2917.600 298.330 2924.800 298.780 ;
        RECT 2904.045 298.030 2924.800 298.330 ;
        RECT 2904.045 298.015 2904.375 298.030 ;
        RECT 2917.600 297.580 2924.800 298.030 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 3504.960 642.090 3505.020 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 641.770 3504.820 1095.190 3504.960 ;
        RECT 641.770 3504.760 642.090 3504.820 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
      LAYER via ;
        RECT 641.800 3504.760 642.060 3505.020 ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 641.800 3504.730 642.060 3505.050 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 641.860 999.330 642.000 3504.730 ;
        RECT 642.610 999.330 642.890 1000.000 ;
        RECT 641.860 999.190 642.890 999.330 ;
        RECT 642.610 996.000 642.890 999.190 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 3500.880 662.790 3500.940 ;
        RECT 770.570 3500.880 770.890 3500.940 ;
        RECT 662.470 3500.740 770.890 3500.880 ;
        RECT 662.470 3500.680 662.790 3500.740 ;
        RECT 770.570 3500.680 770.890 3500.740 ;
      LAYER via ;
        RECT 662.500 3500.680 662.760 3500.940 ;
        RECT 770.600 3500.680 770.860 3500.940 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3500.970 770.800 3517.600 ;
        RECT 662.500 3500.650 662.760 3500.970 ;
        RECT 770.600 3500.650 770.860 3500.970 ;
        RECT 662.560 999.330 662.700 3500.650 ;
        RECT 663.770 999.330 664.050 1000.000 ;
        RECT 662.560 999.190 664.050 999.330 ;
        RECT 663.770 996.000 664.050 999.190 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3501.220 446.130 3501.280 ;
        RECT 679.490 3501.220 679.810 3501.280 ;
        RECT 445.810 3501.080 679.810 3501.220 ;
        RECT 445.810 3501.020 446.130 3501.080 ;
        RECT 679.490 3501.020 679.810 3501.080 ;
        RECT 679.490 1014.120 679.810 1014.180 ;
        RECT 683.630 1014.120 683.950 1014.180 ;
        RECT 679.490 1013.980 683.950 1014.120 ;
        RECT 679.490 1013.920 679.810 1013.980 ;
        RECT 683.630 1013.920 683.950 1013.980 ;
      LAYER via ;
        RECT 445.840 3501.020 446.100 3501.280 ;
        RECT 679.520 3501.020 679.780 3501.280 ;
        RECT 679.520 1013.920 679.780 1014.180 ;
        RECT 683.660 1013.920 683.920 1014.180 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3501.310 446.040 3517.600 ;
        RECT 445.840 3500.990 446.100 3501.310 ;
        RECT 679.520 3500.990 679.780 3501.310 ;
        RECT 679.580 1014.210 679.720 3500.990 ;
        RECT 679.520 1013.890 679.780 1014.210 ;
        RECT 683.660 1013.890 683.920 1014.210 ;
        RECT 683.720 999.330 683.860 1013.890 ;
        RECT 684.930 999.330 685.210 1000.000 ;
        RECT 683.720 999.190 685.210 999.330 ;
        RECT 684.930 996.000 685.210 999.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3504.620 121.830 3504.680 ;
        RECT 703.870 3504.620 704.190 3504.680 ;
        RECT 121.510 3504.480 704.190 3504.620 ;
        RECT 121.510 3504.420 121.830 3504.480 ;
        RECT 703.870 3504.420 704.190 3504.480 ;
      LAYER via ;
        RECT 121.540 3504.420 121.800 3504.680 ;
        RECT 703.900 3504.420 704.160 3504.680 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3504.710 121.740 3517.600 ;
        RECT 121.540 3504.390 121.800 3504.710 ;
        RECT 703.900 3504.390 704.160 3504.710 ;
        RECT 703.960 1048.870 704.100 3504.390 ;
        RECT 703.960 1048.730 704.560 1048.870 ;
        RECT 704.420 999.330 704.560 1048.730 ;
        RECT 706.550 999.330 706.830 1000.000 ;
        RECT 704.420 999.190 706.830 999.330 ;
        RECT 706.550 996.000 706.830 999.190 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3354.000 17.410 3354.060 ;
        RECT 724.570 3354.000 724.890 3354.060 ;
        RECT 17.090 3353.860 724.890 3354.000 ;
        RECT 17.090 3353.800 17.410 3353.860 ;
        RECT 724.570 3353.800 724.890 3353.860 ;
      LAYER via ;
        RECT 17.120 3353.800 17.380 3354.060 ;
        RECT 724.600 3353.800 724.860 3354.060 ;
      LAYER met2 ;
        RECT 17.110 3355.955 17.390 3356.325 ;
        RECT 17.180 3354.090 17.320 3355.955 ;
        RECT 17.120 3353.770 17.380 3354.090 ;
        RECT 724.600 3353.770 724.860 3354.090 ;
        RECT 724.660 1048.870 724.800 3353.770 ;
        RECT 724.660 1048.730 725.720 1048.870 ;
        RECT 725.580 999.330 725.720 1048.730 ;
        RECT 727.710 999.330 727.990 1000.000 ;
        RECT 725.580 999.190 727.990 999.330 ;
        RECT 727.710 996.000 727.990 999.190 ;
      LAYER via2 ;
        RECT 17.110 3356.000 17.390 3356.280 ;
      LAYER met3 ;
        RECT -4.800 3356.290 2.400 3356.740 ;
        RECT 17.085 3356.290 17.415 3356.305 ;
        RECT -4.800 3355.990 17.415 3356.290 ;
        RECT -4.800 3355.540 2.400 3355.990 ;
        RECT 17.085 3355.975 17.415 3355.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 3091.520 16.030 3091.580 ;
        RECT 745.270 3091.520 745.590 3091.580 ;
        RECT 15.710 3091.380 745.590 3091.520 ;
        RECT 15.710 3091.320 16.030 3091.380 ;
        RECT 745.270 3091.320 745.590 3091.380 ;
      LAYER via ;
        RECT 15.740 3091.320 16.000 3091.580 ;
        RECT 745.300 3091.320 745.560 3091.580 ;
      LAYER met2 ;
        RECT 15.730 3095.515 16.010 3095.885 ;
        RECT 15.800 3091.610 15.940 3095.515 ;
        RECT 15.740 3091.290 16.000 3091.610 ;
        RECT 745.300 3091.290 745.560 3091.610 ;
        RECT 745.360 1048.870 745.500 3091.290 ;
        RECT 745.360 1048.730 746.880 1048.870 ;
        RECT 746.740 999.330 746.880 1048.730 ;
        RECT 748.870 999.330 749.150 1000.000 ;
        RECT 746.740 999.190 749.150 999.330 ;
        RECT 748.870 996.000 749.150 999.190 ;
      LAYER via2 ;
        RECT 15.730 3095.560 16.010 3095.840 ;
      LAYER met3 ;
        RECT -4.800 3095.850 2.400 3096.300 ;
        RECT 15.705 3095.850 16.035 3095.865 ;
        RECT -4.800 3095.550 16.035 3095.850 ;
        RECT -4.800 3095.100 2.400 3095.550 ;
        RECT 15.705 3095.535 16.035 3095.550 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2829.380 17.410 2829.440 ;
        RECT 765.970 2829.380 766.290 2829.440 ;
        RECT 17.090 2829.240 766.290 2829.380 ;
        RECT 17.090 2829.180 17.410 2829.240 ;
        RECT 765.970 2829.180 766.290 2829.240 ;
      LAYER via ;
        RECT 17.120 2829.180 17.380 2829.440 ;
        RECT 766.000 2829.180 766.260 2829.440 ;
      LAYER met2 ;
        RECT 17.110 2834.395 17.390 2834.765 ;
        RECT 17.180 2829.470 17.320 2834.395 ;
        RECT 17.120 2829.150 17.380 2829.470 ;
        RECT 766.000 2829.150 766.260 2829.470 ;
        RECT 766.060 1048.870 766.200 2829.150 ;
        RECT 766.060 1048.730 768.040 1048.870 ;
        RECT 767.900 999.330 768.040 1048.730 ;
        RECT 770.030 999.330 770.310 1000.000 ;
        RECT 767.900 999.190 770.310 999.330 ;
        RECT 770.030 996.000 770.310 999.190 ;
      LAYER via2 ;
        RECT 17.110 2834.440 17.390 2834.720 ;
      LAYER met3 ;
        RECT -4.800 2834.730 2.400 2835.180 ;
        RECT 17.085 2834.730 17.415 2834.745 ;
        RECT -4.800 2834.430 17.415 2834.730 ;
        RECT -4.800 2833.980 2.400 2834.430 ;
        RECT 17.085 2834.415 17.415 2834.430 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2574.040 17.410 2574.100 ;
        RECT 786.670 2574.040 786.990 2574.100 ;
        RECT 17.090 2573.900 786.990 2574.040 ;
        RECT 17.090 2573.840 17.410 2573.900 ;
        RECT 786.670 2573.840 786.990 2573.900 ;
      LAYER via ;
        RECT 17.120 2573.840 17.380 2574.100 ;
        RECT 786.700 2573.840 786.960 2574.100 ;
      LAYER met2 ;
        RECT 17.110 2573.955 17.390 2574.325 ;
        RECT 17.120 2573.810 17.380 2573.955 ;
        RECT 786.700 2573.810 786.960 2574.130 ;
        RECT 786.760 1048.870 786.900 2573.810 ;
        RECT 786.760 1048.730 789.200 1048.870 ;
        RECT 789.060 999.330 789.200 1048.730 ;
        RECT 791.190 999.330 791.470 1000.000 ;
        RECT 789.060 999.190 791.470 999.330 ;
        RECT 791.190 996.000 791.470 999.190 ;
      LAYER via2 ;
        RECT 17.110 2574.000 17.390 2574.280 ;
      LAYER met3 ;
        RECT -4.800 2574.290 2.400 2574.740 ;
        RECT 17.085 2574.290 17.415 2574.305 ;
        RECT -4.800 2573.990 17.415 2574.290 ;
        RECT -4.800 2573.540 2.400 2573.990 ;
        RECT 17.085 2573.975 17.415 2573.990 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2311.900 16.490 2311.960 ;
        RECT 807.370 2311.900 807.690 2311.960 ;
        RECT 16.170 2311.760 807.690 2311.900 ;
        RECT 16.170 2311.700 16.490 2311.760 ;
        RECT 807.370 2311.700 807.690 2311.760 ;
      LAYER via ;
        RECT 16.200 2311.700 16.460 2311.960 ;
        RECT 807.400 2311.700 807.660 2311.960 ;
      LAYER met2 ;
        RECT 16.190 2312.835 16.470 2313.205 ;
        RECT 16.260 2311.990 16.400 2312.835 ;
        RECT 16.200 2311.670 16.460 2311.990 ;
        RECT 807.400 2311.670 807.660 2311.990 ;
        RECT 807.460 1048.870 807.600 2311.670 ;
        RECT 807.460 1048.730 811.280 1048.870 ;
        RECT 811.140 999.330 811.280 1048.730 ;
        RECT 812.810 999.330 813.090 1000.000 ;
        RECT 811.140 999.190 813.090 999.330 ;
        RECT 812.810 996.000 813.090 999.190 ;
      LAYER via2 ;
        RECT 16.190 2312.880 16.470 2313.160 ;
      LAYER met3 ;
        RECT -4.800 2313.170 2.400 2313.620 ;
        RECT 16.165 2313.170 16.495 2313.185 ;
        RECT -4.800 2312.870 16.495 2313.170 ;
        RECT -4.800 2312.420 2.400 2312.870 ;
        RECT 16.165 2312.855 16.495 2312.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2049.420 16.030 2049.480 ;
        RECT 828.070 2049.420 828.390 2049.480 ;
        RECT 15.710 2049.280 828.390 2049.420 ;
        RECT 15.710 2049.220 16.030 2049.280 ;
        RECT 828.070 2049.220 828.390 2049.280 ;
      LAYER via ;
        RECT 15.740 2049.220 16.000 2049.480 ;
        RECT 828.100 2049.220 828.360 2049.480 ;
      LAYER met2 ;
        RECT 15.730 2052.395 16.010 2052.765 ;
        RECT 15.800 2049.510 15.940 2052.395 ;
        RECT 15.740 2049.190 16.000 2049.510 ;
        RECT 828.100 2049.190 828.360 2049.510 ;
        RECT 828.160 1048.870 828.300 2049.190 ;
        RECT 828.160 1048.730 832.440 1048.870 ;
        RECT 832.300 999.330 832.440 1048.730 ;
        RECT 833.970 999.330 834.250 1000.000 ;
        RECT 832.300 999.190 834.250 999.330 ;
        RECT 833.970 996.000 834.250 999.190 ;
      LAYER via2 ;
        RECT 15.730 2052.440 16.010 2052.720 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 15.705 2052.730 16.035 2052.745 ;
        RECT -4.800 2052.430 16.035 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 15.705 2052.415 16.035 2052.430 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 261.810 1009.020 262.130 1009.080 ;
        RECT 1100.390 1009.020 1100.710 1009.080 ;
        RECT 261.810 1008.880 1100.710 1009.020 ;
        RECT 261.810 1008.820 262.130 1008.880 ;
        RECT 1100.390 1008.820 1100.710 1008.880 ;
        RECT 1100.390 503.440 1100.710 503.500 ;
        RECT 2900.370 503.440 2900.690 503.500 ;
        RECT 1100.390 503.300 2900.690 503.440 ;
        RECT 1100.390 503.240 1100.710 503.300 ;
        RECT 2900.370 503.240 2900.690 503.300 ;
      LAYER via ;
        RECT 261.840 1008.820 262.100 1009.080 ;
        RECT 1100.420 1008.820 1100.680 1009.080 ;
        RECT 1100.420 503.240 1100.680 503.500 ;
        RECT 2900.400 503.240 2900.660 503.500 ;
      LAYER met2 ;
        RECT 261.840 1008.790 262.100 1009.110 ;
        RECT 1100.420 1008.790 1100.680 1009.110 ;
        RECT 259.890 999.330 260.170 1000.000 ;
        RECT 261.900 999.330 262.040 1008.790 ;
        RECT 259.890 999.190 262.040 999.330 ;
        RECT 259.890 996.000 260.170 999.190 ;
        RECT 1100.480 503.530 1100.620 1008.790 ;
        RECT 1100.420 503.210 1100.680 503.530 ;
        RECT 2900.400 503.210 2900.660 503.530 ;
        RECT 2900.460 497.605 2900.600 503.210 ;
        RECT 2900.390 497.235 2900.670 497.605 ;
      LAYER via2 ;
        RECT 2900.390 497.280 2900.670 497.560 ;
      LAYER met3 ;
        RECT 2900.365 497.570 2900.695 497.585 ;
        RECT 2917.600 497.570 2924.800 498.020 ;
        RECT 2900.365 497.270 2924.800 497.570 ;
        RECT 2900.365 497.255 2900.695 497.270 ;
        RECT 2917.600 496.820 2924.800 497.270 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1787.280 16.030 1787.340 ;
        RECT 849.230 1787.280 849.550 1787.340 ;
        RECT 15.710 1787.140 849.550 1787.280 ;
        RECT 15.710 1787.080 16.030 1787.140 ;
        RECT 849.230 1787.080 849.550 1787.140 ;
      LAYER via ;
        RECT 15.740 1787.080 16.000 1787.340 ;
        RECT 849.260 1787.080 849.520 1787.340 ;
      LAYER met2 ;
        RECT 15.730 1791.955 16.010 1792.325 ;
        RECT 15.800 1787.370 15.940 1791.955 ;
        RECT 15.740 1787.050 16.000 1787.370 ;
        RECT 849.260 1787.050 849.520 1787.370 ;
        RECT 849.320 1048.870 849.460 1787.050 ;
        RECT 849.320 1048.730 853.600 1048.870 ;
        RECT 853.460 999.330 853.600 1048.730 ;
        RECT 855.130 999.330 855.410 1000.000 ;
        RECT 853.460 999.190 855.410 999.330 ;
        RECT 855.130 996.000 855.410 999.190 ;
      LAYER via2 ;
        RECT 15.730 1792.000 16.010 1792.280 ;
      LAYER met3 ;
        RECT -4.800 1792.290 2.400 1792.740 ;
        RECT 15.705 1792.290 16.035 1792.305 ;
        RECT -4.800 1791.990 16.035 1792.290 ;
        RECT -4.800 1791.540 2.400 1791.990 ;
        RECT 15.705 1791.975 16.035 1791.990 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1525.140 17.870 1525.200 ;
        RECT 876.370 1525.140 876.690 1525.200 ;
        RECT 17.550 1525.000 876.690 1525.140 ;
        RECT 17.550 1524.940 17.870 1525.000 ;
        RECT 876.370 1524.940 876.690 1525.000 ;
      LAYER via ;
        RECT 17.580 1524.940 17.840 1525.200 ;
        RECT 876.400 1524.940 876.660 1525.200 ;
      LAYER met2 ;
        RECT 17.570 1530.835 17.850 1531.205 ;
        RECT 17.640 1525.230 17.780 1530.835 ;
        RECT 17.580 1524.910 17.840 1525.230 ;
        RECT 876.400 1524.910 876.660 1525.230 ;
        RECT 876.460 1048.870 876.600 1524.910 ;
        RECT 876.460 1048.730 877.060 1048.870 ;
        RECT 876.290 999.330 876.570 1000.000 ;
        RECT 876.920 999.330 877.060 1048.730 ;
        RECT 876.290 999.190 877.060 999.330 ;
        RECT 876.290 996.000 876.570 999.190 ;
      LAYER via2 ;
        RECT 17.570 1530.880 17.850 1531.160 ;
      LAYER met3 ;
        RECT -4.800 1531.170 2.400 1531.620 ;
        RECT 17.545 1531.170 17.875 1531.185 ;
        RECT -4.800 1530.870 17.875 1531.170 ;
        RECT -4.800 1530.420 2.400 1530.870 ;
        RECT 17.545 1530.855 17.875 1530.870 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1269.800 17.870 1269.860 ;
        RECT 872.690 1269.800 873.010 1269.860 ;
        RECT 17.550 1269.660 873.010 1269.800 ;
        RECT 17.550 1269.600 17.870 1269.660 ;
        RECT 872.690 1269.600 873.010 1269.660 ;
        RECT 872.690 1014.120 873.010 1014.180 ;
        RECT 897.070 1014.120 897.390 1014.180 ;
        RECT 872.690 1013.980 897.390 1014.120 ;
        RECT 872.690 1013.920 873.010 1013.980 ;
        RECT 897.070 1013.920 897.390 1013.980 ;
      LAYER via ;
        RECT 17.580 1269.600 17.840 1269.860 ;
        RECT 872.720 1269.600 872.980 1269.860 ;
        RECT 872.720 1013.920 872.980 1014.180 ;
        RECT 897.100 1013.920 897.360 1014.180 ;
      LAYER met2 ;
        RECT 17.570 1270.395 17.850 1270.765 ;
        RECT 17.640 1269.890 17.780 1270.395 ;
        RECT 17.580 1269.570 17.840 1269.890 ;
        RECT 872.720 1269.570 872.980 1269.890 ;
        RECT 872.780 1014.210 872.920 1269.570 ;
        RECT 872.720 1013.890 872.980 1014.210 ;
        RECT 897.100 1013.890 897.360 1014.210 ;
        RECT 897.160 999.330 897.300 1013.890 ;
        RECT 897.910 999.330 898.190 1000.000 ;
        RECT 897.160 999.190 898.190 999.330 ;
        RECT 897.910 996.000 898.190 999.190 ;
      LAYER via2 ;
        RECT 17.570 1270.440 17.850 1270.720 ;
      LAYER met3 ;
        RECT -4.800 1270.730 2.400 1271.180 ;
        RECT 17.545 1270.730 17.875 1270.745 ;
        RECT -4.800 1270.430 17.875 1270.730 ;
        RECT -4.800 1269.980 2.400 1270.430 ;
        RECT 17.545 1270.415 17.875 1270.430 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1008.680 17.870 1008.740 ;
        RECT 917.770 1008.680 918.090 1008.740 ;
        RECT 17.550 1008.540 918.090 1008.680 ;
        RECT 17.550 1008.480 17.870 1008.540 ;
        RECT 917.770 1008.480 918.090 1008.540 ;
      LAYER via ;
        RECT 17.580 1008.480 17.840 1008.740 ;
        RECT 917.800 1008.480 918.060 1008.740 ;
      LAYER met2 ;
        RECT 17.570 1009.275 17.850 1009.645 ;
        RECT 17.640 1008.770 17.780 1009.275 ;
        RECT 17.580 1008.450 17.840 1008.770 ;
        RECT 917.800 1008.450 918.060 1008.770 ;
        RECT 917.860 999.330 918.000 1008.450 ;
        RECT 919.070 999.330 919.350 1000.000 ;
        RECT 917.860 999.190 919.350 999.330 ;
        RECT 919.070 996.000 919.350 999.190 ;
      LAYER via2 ;
        RECT 17.570 1009.320 17.850 1009.600 ;
      LAYER met3 ;
        RECT -4.800 1009.610 2.400 1010.060 ;
        RECT 17.545 1009.610 17.875 1009.625 ;
        RECT -4.800 1009.310 17.875 1009.610 ;
        RECT -4.800 1008.860 2.400 1009.310 ;
        RECT 17.545 1009.295 17.875 1009.310 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 237.890 998.480 238.210 998.540 ;
        RECT 257.210 998.480 257.530 998.540 ;
        RECT 237.890 998.340 257.530 998.480 ;
        RECT 237.890 998.280 238.210 998.340 ;
        RECT 257.210 998.280 257.530 998.340 ;
        RECT 938.470 997.800 938.790 997.860 ;
        RECT 892.560 997.660 938.790 997.800 ;
        RECT 219.030 997.260 219.350 997.520 ;
        RECT 237.890 997.460 238.210 997.520 ;
        RECT 220.730 997.320 238.210 997.460 ;
        RECT 219.120 997.120 219.260 997.260 ;
        RECT 220.730 997.120 220.870 997.320 ;
        RECT 237.890 997.260 238.210 997.320 ;
        RECT 257.210 997.260 257.530 997.520 ;
        RECT 503.310 997.460 503.630 997.520 ;
        RECT 493.740 997.320 503.630 997.460 ;
        RECT 219.120 996.980 220.870 997.120 ;
        RECT 257.300 996.100 257.440 997.260 ;
        RECT 257.300 995.960 276.070 996.100 ;
        RECT 275.930 995.080 276.070 995.960 ;
        RECT 275.930 994.940 282.970 995.080 ;
        RECT 24.450 994.740 24.770 994.800 ;
        RECT 282.830 994.740 282.970 994.940 ;
        RECT 493.740 994.740 493.880 997.320 ;
        RECT 503.310 997.260 503.630 997.320 ;
        RECT 504.230 997.260 504.550 997.520 ;
        RECT 504.320 996.780 504.460 997.260 ;
        RECT 504.320 996.640 765.970 996.780 ;
        RECT 765.830 996.100 765.970 996.640 ;
        RECT 814.130 996.640 862.570 996.780 ;
        RECT 786.530 996.300 793.570 996.440 ;
        RECT 765.830 995.960 772.870 996.100 ;
        RECT 772.730 995.760 772.870 995.960 ;
        RECT 786.530 995.760 786.670 996.300 ;
        RECT 793.430 996.100 793.570 996.300 ;
        RECT 800.330 996.300 807.370 996.440 ;
        RECT 800.330 996.100 800.470 996.300 ;
        RECT 793.430 995.960 800.470 996.100 ;
        RECT 807.230 996.100 807.370 996.300 ;
        RECT 814.130 996.100 814.270 996.640 ;
        RECT 862.430 996.440 862.570 996.640 ;
        RECT 862.430 996.300 869.470 996.440 ;
        RECT 807.230 995.960 814.270 996.100 ;
        RECT 772.730 995.620 786.670 995.760 ;
        RECT 869.330 995.420 869.470 996.300 ;
        RECT 892.560 995.760 892.700 997.660 ;
        RECT 938.470 997.600 938.790 997.660 ;
        RECT 870.020 995.620 892.700 995.760 ;
        RECT 870.020 995.420 870.160 995.620 ;
        RECT 869.330 995.280 870.160 995.420 ;
        RECT 24.450 994.600 131.170 994.740 ;
        RECT 282.830 994.600 493.880 994.740 ;
        RECT 24.450 994.540 24.770 994.600 ;
        RECT 131.030 994.060 131.170 994.600 ;
        RECT 199.250 994.060 199.570 994.120 ;
        RECT 131.030 993.920 199.570 994.060 ;
        RECT 199.250 993.860 199.570 993.920 ;
        RECT 13.870 749.600 14.190 749.660 ;
        RECT 24.450 749.600 24.770 749.660 ;
        RECT 13.870 749.460 24.770 749.600 ;
        RECT 13.870 749.400 14.190 749.460 ;
        RECT 24.450 749.400 24.770 749.460 ;
      LAYER via ;
        RECT 237.920 998.280 238.180 998.540 ;
        RECT 257.240 998.280 257.500 998.540 ;
        RECT 219.060 997.260 219.320 997.520 ;
        RECT 237.920 997.260 238.180 997.520 ;
        RECT 257.240 997.260 257.500 997.520 ;
        RECT 24.480 994.540 24.740 994.800 ;
        RECT 503.340 997.260 503.600 997.520 ;
        RECT 504.260 997.260 504.520 997.520 ;
        RECT 938.500 997.600 938.760 997.860 ;
        RECT 199.280 993.860 199.540 994.120 ;
        RECT 13.900 749.400 14.160 749.660 ;
        RECT 24.480 749.400 24.740 749.660 ;
      LAYER met2 ;
        RECT 237.920 998.250 238.180 998.570 ;
        RECT 257.240 998.250 257.500 998.570 ;
        RECT 503.400 998.510 504.460 998.650 ;
        RECT 237.980 997.550 238.120 998.250 ;
        RECT 257.300 997.550 257.440 998.250 ;
        RECT 503.400 997.550 503.540 998.510 ;
        RECT 504.320 997.550 504.460 998.510 ;
        RECT 940.230 997.970 940.510 1000.000 ;
        RECT 938.560 997.890 940.510 997.970 ;
        RECT 938.500 997.830 940.510 997.890 ;
        RECT 938.500 997.570 938.760 997.830 ;
        RECT 219.060 997.405 219.320 997.550 ;
        RECT 199.270 997.035 199.550 997.405 ;
        RECT 219.050 997.035 219.330 997.405 ;
        RECT 237.920 997.230 238.180 997.550 ;
        RECT 257.240 997.230 257.500 997.550 ;
        RECT 503.340 997.230 503.600 997.550 ;
        RECT 504.260 997.230 504.520 997.550 ;
        RECT 24.480 994.510 24.740 994.830 ;
        RECT 24.540 749.690 24.680 994.510 ;
        RECT 199.340 994.150 199.480 997.035 ;
        RECT 940.230 996.000 940.510 997.830 ;
        RECT 199.280 993.830 199.540 994.150 ;
        RECT 13.900 749.370 14.160 749.690 ;
        RECT 24.480 749.370 24.740 749.690 ;
        RECT 13.960 749.205 14.100 749.370 ;
        RECT 13.890 748.835 14.170 749.205 ;
      LAYER via2 ;
        RECT 199.270 997.080 199.550 997.360 ;
        RECT 219.050 997.080 219.330 997.360 ;
        RECT 13.890 748.880 14.170 749.160 ;
      LAYER met3 ;
        RECT 199.245 997.370 199.575 997.385 ;
        RECT 219.025 997.370 219.355 997.385 ;
        RECT 199.245 997.070 219.355 997.370 ;
        RECT 199.245 997.055 199.575 997.070 ;
        RECT 219.025 997.055 219.355 997.070 ;
        RECT -4.800 749.170 2.400 749.620 ;
        RECT 13.865 749.170 14.195 749.185 ;
        RECT -4.800 748.870 14.195 749.170 ;
        RECT -4.800 748.420 2.400 748.870 ;
        RECT 13.865 748.855 14.195 748.870 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.390 1008.000 19.710 1008.060 ;
        RECT 959.630 1008.000 959.950 1008.060 ;
        RECT 19.390 1007.860 959.950 1008.000 ;
        RECT 19.390 1007.800 19.710 1007.860 ;
        RECT 959.630 1007.800 959.950 1007.860 ;
      LAYER via ;
        RECT 19.420 1007.800 19.680 1008.060 ;
        RECT 959.660 1007.800 959.920 1008.060 ;
      LAYER met2 ;
        RECT 19.420 1007.770 19.680 1008.090 ;
        RECT 959.660 1007.770 959.920 1008.090 ;
        RECT 19.480 488.085 19.620 1007.770 ;
        RECT 959.720 999.330 959.860 1007.770 ;
        RECT 961.390 999.330 961.670 1000.000 ;
        RECT 959.720 999.190 961.670 999.330 ;
        RECT 961.390 996.000 961.670 999.190 ;
        RECT 19.410 487.715 19.690 488.085 ;
      LAYER via2 ;
        RECT 19.410 487.760 19.690 488.040 ;
      LAYER met3 ;
        RECT -4.800 488.050 2.400 488.500 ;
        RECT 19.385 488.050 19.715 488.065 ;
        RECT -4.800 487.750 19.715 488.050 ;
        RECT -4.800 487.300 2.400 487.750 ;
        RECT 19.385 487.735 19.715 487.750 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 1007.660 18.330 1007.720 ;
        RECT 981.710 1007.660 982.030 1007.720 ;
        RECT 18.010 1007.520 982.030 1007.660 ;
        RECT 18.010 1007.460 18.330 1007.520 ;
        RECT 981.710 1007.460 982.030 1007.520 ;
      LAYER via ;
        RECT 18.040 1007.460 18.300 1007.720 ;
        RECT 981.740 1007.460 982.000 1007.720 ;
      LAYER met2 ;
        RECT 18.040 1007.430 18.300 1007.750 ;
        RECT 981.740 1007.430 982.000 1007.750 ;
        RECT 18.100 292.925 18.240 1007.430 ;
        RECT 981.800 999.330 981.940 1007.430 ;
        RECT 983.010 999.330 983.290 1000.000 ;
        RECT 981.800 999.190 983.290 999.330 ;
        RECT 983.010 996.000 983.290 999.190 ;
        RECT 18.030 292.555 18.310 292.925 ;
      LAYER via2 ;
        RECT 18.030 292.600 18.310 292.880 ;
      LAYER met3 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 18.005 292.890 18.335 292.905 ;
        RECT -4.800 292.590 18.335 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 18.005 292.575 18.335 292.590 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 1000.435 1003.170 1000.805 ;
        RECT 1002.960 999.330 1003.100 1000.435 ;
        RECT 1004.170 999.330 1004.450 1000.000 ;
        RECT 1002.960 999.190 1004.450 999.330 ;
        RECT 1004.170 996.000 1004.450 999.190 ;
      LAYER via2 ;
        RECT 1002.890 1000.480 1003.170 1000.760 ;
      LAYER met3 ;
        RECT 16.830 1000.770 17.210 1000.780 ;
        RECT 1002.865 1000.770 1003.195 1000.785 ;
        RECT 16.830 1000.470 1003.195 1000.770 ;
        RECT 16.830 1000.460 17.210 1000.470 ;
        RECT 1002.865 1000.455 1003.195 1000.470 ;
        RECT -4.800 97.050 2.400 97.500 ;
        RECT 16.830 97.050 17.210 97.060 ;
        RECT -4.800 96.750 17.210 97.050 ;
        RECT -4.800 96.300 2.400 96.750 ;
        RECT 16.830 96.740 17.210 96.750 ;
      LAYER via3 ;
        RECT 16.860 1000.460 17.180 1000.780 ;
        RECT 16.860 96.740 17.180 97.060 ;
      LAYER met4 ;
        RECT 16.855 1000.455 17.185 1000.785 ;
        RECT 16.870 97.065 17.170 1000.455 ;
        RECT 16.855 96.735 17.185 97.065 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.510 1010.040 282.830 1010.100 ;
        RECT 1101.310 1010.040 1101.630 1010.100 ;
        RECT 282.510 1009.900 1101.630 1010.040 ;
        RECT 282.510 1009.840 282.830 1009.900 ;
        RECT 1101.310 1009.840 1101.630 1009.900 ;
        RECT 1101.310 696.900 1101.630 696.960 ;
        RECT 2899.910 696.900 2900.230 696.960 ;
        RECT 1101.310 696.760 2900.230 696.900 ;
        RECT 1101.310 696.700 1101.630 696.760 ;
        RECT 2899.910 696.700 2900.230 696.760 ;
      LAYER via ;
        RECT 282.540 1009.840 282.800 1010.100 ;
        RECT 1101.340 1009.840 1101.600 1010.100 ;
        RECT 1101.340 696.700 1101.600 696.960 ;
        RECT 2899.940 696.700 2900.200 696.960 ;
      LAYER met2 ;
        RECT 282.540 1009.810 282.800 1010.130 ;
        RECT 1101.340 1009.810 1101.600 1010.130 ;
        RECT 281.050 999.330 281.330 1000.000 ;
        RECT 282.600 999.330 282.740 1009.810 ;
        RECT 281.050 999.190 282.740 999.330 ;
        RECT 281.050 996.000 281.330 999.190 ;
        RECT 1101.400 696.990 1101.540 1009.810 ;
        RECT 1101.340 696.670 1101.600 696.990 ;
        RECT 2899.940 696.845 2900.200 696.990 ;
        RECT 2899.930 696.475 2900.210 696.845 ;
      LAYER via2 ;
        RECT 2899.930 696.520 2900.210 696.800 ;
      LAYER met3 ;
        RECT 2899.905 696.810 2900.235 696.825 ;
        RECT 2917.600 696.810 2924.800 697.260 ;
        RECT 2899.905 696.510 2924.800 696.810 ;
        RECT 2899.905 696.495 2900.235 696.510 ;
        RECT 2917.600 696.060 2924.800 696.510 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.210 1011.740 303.530 1011.800 ;
        RECT 1102.690 1011.740 1103.010 1011.800 ;
        RECT 303.210 1011.600 1103.010 1011.740 ;
        RECT 303.210 1011.540 303.530 1011.600 ;
        RECT 1102.690 1011.540 1103.010 1011.600 ;
        RECT 1102.690 896.820 1103.010 896.880 ;
        RECT 2899.910 896.820 2900.230 896.880 ;
        RECT 1102.690 896.680 2900.230 896.820 ;
        RECT 1102.690 896.620 1103.010 896.680 ;
        RECT 2899.910 896.620 2900.230 896.680 ;
      LAYER via ;
        RECT 303.240 1011.540 303.500 1011.800 ;
        RECT 1102.720 1011.540 1102.980 1011.800 ;
        RECT 1102.720 896.620 1102.980 896.880 ;
        RECT 2899.940 896.620 2900.200 896.880 ;
      LAYER met2 ;
        RECT 303.240 1011.510 303.500 1011.830 ;
        RECT 1102.720 1011.510 1102.980 1011.830 ;
        RECT 302.210 999.330 302.490 1000.000 ;
        RECT 303.300 999.330 303.440 1011.510 ;
        RECT 302.210 999.190 303.440 999.330 ;
        RECT 302.210 996.000 302.490 999.190 ;
        RECT 1102.780 896.910 1102.920 1011.510 ;
        RECT 1102.720 896.590 1102.980 896.910 ;
        RECT 2899.940 896.590 2900.200 896.910 ;
        RECT 2900.000 896.085 2900.140 896.590 ;
        RECT 2899.930 895.715 2900.210 896.085 ;
      LAYER via2 ;
        RECT 2899.930 895.760 2900.210 896.040 ;
      LAYER met3 ;
        RECT 2899.905 896.050 2900.235 896.065 ;
        RECT 2917.600 896.050 2924.800 896.500 ;
        RECT 2899.905 895.750 2924.800 896.050 ;
        RECT 2899.905 895.735 2900.235 895.750 ;
        RECT 2917.600 895.300 2924.800 895.750 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.470 1090.280 317.790 1090.340 ;
        RECT 2900.830 1090.280 2901.150 1090.340 ;
        RECT 317.470 1090.140 2901.150 1090.280 ;
        RECT 317.470 1090.080 317.790 1090.140 ;
        RECT 2900.830 1090.080 2901.150 1090.140 ;
      LAYER via ;
        RECT 317.500 1090.080 317.760 1090.340 ;
        RECT 2900.860 1090.080 2901.120 1090.340 ;
      LAYER met2 ;
        RECT 2900.850 1094.955 2901.130 1095.325 ;
        RECT 2900.920 1090.370 2901.060 1094.955 ;
        RECT 317.500 1090.050 317.760 1090.370 ;
        RECT 2900.860 1090.050 2901.120 1090.370 ;
        RECT 317.560 1048.870 317.700 1090.050 ;
        RECT 317.560 1048.730 321.840 1048.870 ;
        RECT 321.700 999.330 321.840 1048.730 ;
        RECT 323.370 999.330 323.650 1000.000 ;
        RECT 321.700 999.190 323.650 999.330 ;
        RECT 323.370 996.000 323.650 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1095.000 2901.130 1095.280 ;
      LAYER met3 ;
        RECT 2900.825 1095.290 2901.155 1095.305 ;
        RECT 2917.600 1095.290 2924.800 1095.740 ;
        RECT 2900.825 1094.990 2924.800 1095.290 ;
        RECT 2900.825 1094.975 2901.155 1094.990 ;
        RECT 2917.600 1094.540 2924.800 1094.990 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 1290.540 345.390 1290.600 ;
        RECT 2899.910 1290.540 2900.230 1290.600 ;
        RECT 345.070 1290.400 2900.230 1290.540 ;
        RECT 345.070 1290.340 345.390 1290.400 ;
        RECT 2899.910 1290.340 2900.230 1290.400 ;
      LAYER via ;
        RECT 345.100 1290.340 345.360 1290.600 ;
        RECT 2899.940 1290.340 2900.200 1290.600 ;
      LAYER met2 ;
        RECT 2899.930 1294.195 2900.210 1294.565 ;
        RECT 2900.000 1290.630 2900.140 1294.195 ;
        RECT 345.100 1290.310 345.360 1290.630 ;
        RECT 2899.940 1290.310 2900.200 1290.630 ;
        RECT 345.160 1048.870 345.300 1290.310 ;
        RECT 345.160 1048.730 345.760 1048.870 ;
        RECT 344.990 999.330 345.270 1000.000 ;
        RECT 345.620 999.330 345.760 1048.730 ;
        RECT 344.990 999.190 345.760 999.330 ;
        RECT 344.990 996.000 345.270 999.190 ;
      LAYER via2 ;
        RECT 2899.930 1294.240 2900.210 1294.520 ;
      LAYER met3 ;
        RECT 2899.905 1294.530 2900.235 1294.545 ;
        RECT 2917.600 1294.530 2924.800 1294.980 ;
        RECT 2899.905 1294.230 2924.800 1294.530 ;
        RECT 2899.905 1294.215 2900.235 1294.230 ;
        RECT 2917.600 1293.780 2924.800 1294.230 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 1559.480 366.090 1559.540 ;
        RECT 2900.830 1559.480 2901.150 1559.540 ;
        RECT 365.770 1559.340 2901.150 1559.480 ;
        RECT 365.770 1559.280 366.090 1559.340 ;
        RECT 2900.830 1559.280 2901.150 1559.340 ;
      LAYER via ;
        RECT 365.800 1559.280 366.060 1559.540 ;
        RECT 2900.860 1559.280 2901.120 1559.540 ;
      LAYER met2 ;
        RECT 2900.850 1560.075 2901.130 1560.445 ;
        RECT 2900.920 1559.570 2901.060 1560.075 ;
        RECT 365.800 1559.250 366.060 1559.570 ;
        RECT 2900.860 1559.250 2901.120 1559.570 ;
        RECT 365.860 999.330 366.000 1559.250 ;
        RECT 366.150 999.330 366.430 1000.000 ;
        RECT 365.860 999.190 366.430 999.330 ;
        RECT 366.150 996.000 366.430 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1560.120 2901.130 1560.400 ;
      LAYER met3 ;
        RECT 2900.825 1560.410 2901.155 1560.425 ;
        RECT 2917.600 1560.410 2924.800 1560.860 ;
        RECT 2900.825 1560.110 2924.800 1560.410 ;
        RECT 2900.825 1560.095 2901.155 1560.110 ;
        RECT 2917.600 1559.660 2924.800 1560.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.470 1821.960 386.790 1822.020 ;
        RECT 2898.990 1821.960 2899.310 1822.020 ;
        RECT 386.470 1821.820 2899.310 1821.960 ;
        RECT 386.470 1821.760 386.790 1821.820 ;
        RECT 2898.990 1821.760 2899.310 1821.820 ;
      LAYER via ;
        RECT 386.500 1821.760 386.760 1822.020 ;
        RECT 2899.020 1821.760 2899.280 1822.020 ;
      LAYER met2 ;
        RECT 2899.010 1825.275 2899.290 1825.645 ;
        RECT 2899.080 1822.050 2899.220 1825.275 ;
        RECT 386.500 1821.730 386.760 1822.050 ;
        RECT 2899.020 1821.730 2899.280 1822.050 ;
        RECT 386.560 999.330 386.700 1821.730 ;
        RECT 387.310 999.330 387.590 1000.000 ;
        RECT 386.560 999.190 387.590 999.330 ;
        RECT 387.310 996.000 387.590 999.190 ;
      LAYER via2 ;
        RECT 2899.010 1825.320 2899.290 1825.600 ;
      LAYER met3 ;
        RECT 2898.985 1825.610 2899.315 1825.625 ;
        RECT 2917.600 1825.610 2924.800 1826.060 ;
        RECT 2898.985 1825.310 2924.800 1825.610 ;
        RECT 2898.985 1825.295 2899.315 1825.310 ;
        RECT 2917.600 1824.860 2924.800 1825.310 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 2090.900 407.490 2090.960 ;
        RECT 2900.830 2090.900 2901.150 2090.960 ;
        RECT 407.170 2090.760 2901.150 2090.900 ;
        RECT 407.170 2090.700 407.490 2090.760 ;
        RECT 2900.830 2090.700 2901.150 2090.760 ;
      LAYER via ;
        RECT 407.200 2090.700 407.460 2090.960 ;
        RECT 2900.860 2090.700 2901.120 2090.960 ;
      LAYER met2 ;
        RECT 2900.850 2091.155 2901.130 2091.525 ;
        RECT 2900.920 2090.990 2901.060 2091.155 ;
        RECT 407.200 2090.670 407.460 2090.990 ;
        RECT 2900.860 2090.670 2901.120 2090.990 ;
        RECT 407.260 999.330 407.400 2090.670 ;
        RECT 408.470 999.330 408.750 1000.000 ;
        RECT 407.260 999.190 408.750 999.330 ;
        RECT 408.470 996.000 408.750 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2091.200 2901.130 2091.480 ;
      LAYER met3 ;
        RECT 2900.825 2091.490 2901.155 2091.505 ;
        RECT 2917.600 2091.490 2924.800 2091.940 ;
        RECT 2900.825 2091.190 2924.800 2091.490 ;
        RECT 2900.825 2091.175 2901.155 2091.190 ;
        RECT 2917.600 2090.740 2924.800 2091.190 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.350 393.620 192.670 393.680 ;
        RECT 393.830 393.620 394.150 393.680 ;
        RECT 192.350 393.480 394.150 393.620 ;
        RECT 192.350 393.420 192.670 393.480 ;
        RECT 393.830 393.420 394.150 393.480 ;
        RECT 393.830 32.200 394.150 32.260 ;
        RECT 579.210 32.200 579.530 32.260 ;
        RECT 393.830 32.060 579.530 32.200 ;
        RECT 393.830 32.000 394.150 32.060 ;
        RECT 579.210 32.000 579.530 32.060 ;
        RECT 579.210 20.640 579.530 20.700 ;
        RECT 629.350 20.640 629.670 20.700 ;
        RECT 579.210 20.500 629.670 20.640 ;
        RECT 579.210 20.440 579.530 20.500 ;
        RECT 629.350 20.440 629.670 20.500 ;
      LAYER via ;
        RECT 192.380 393.420 192.640 393.680 ;
        RECT 393.860 393.420 394.120 393.680 ;
        RECT 393.860 32.000 394.120 32.260 ;
        RECT 579.240 32.000 579.500 32.260 ;
        RECT 579.240 20.440 579.500 20.700 ;
        RECT 629.380 20.440 629.640 20.700 ;
      LAYER met2 ;
        RECT 192.370 441.475 192.650 441.845 ;
        RECT 192.440 393.710 192.580 441.475 ;
        RECT 393.290 400.250 393.570 404.000 ;
        RECT 393.290 400.110 394.060 400.250 ;
        RECT 393.290 400.000 393.570 400.110 ;
        RECT 393.920 393.710 394.060 400.110 ;
        RECT 192.380 393.390 192.640 393.710 ;
        RECT 393.860 393.390 394.120 393.710 ;
        RECT 393.920 32.290 394.060 393.390 ;
        RECT 393.860 31.970 394.120 32.290 ;
        RECT 579.240 31.970 579.500 32.290 ;
        RECT 579.300 20.730 579.440 31.970 ;
        RECT 579.240 20.410 579.500 20.730 ;
        RECT 629.380 20.410 629.640 20.730 ;
        RECT 629.440 2.400 629.580 20.410 ;
        RECT 629.230 -4.800 629.790 2.400 ;
      LAYER via2 ;
        RECT 192.370 441.520 192.650 441.800 ;
      LAYER met3 ;
        RECT 200.000 442.880 204.000 443.480 ;
        RECT 192.345 441.810 192.675 441.825 ;
        RECT 200.870 441.810 201.170 442.880 ;
        RECT 192.345 441.510 201.170 441.810 ;
        RECT 192.345 441.495 192.675 441.510 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 939.850 108.700 940.170 108.760 ;
        RECT 2401.270 108.700 2401.590 108.760 ;
        RECT 939.850 108.560 2401.590 108.700 ;
        RECT 939.850 108.500 940.170 108.560 ;
        RECT 2401.270 108.500 2401.590 108.560 ;
      LAYER via ;
        RECT 939.880 108.500 940.140 108.760 ;
        RECT 2401.300 108.500 2401.560 108.760 ;
      LAYER met2 ;
        RECT 940.230 400.250 940.510 404.000 ;
        RECT 939.940 400.110 940.510 400.250 ;
        RECT 939.940 108.790 940.080 400.110 ;
        RECT 940.230 400.000 940.510 400.110 ;
        RECT 939.880 108.470 940.140 108.790 ;
        RECT 2401.300 108.470 2401.560 108.790 ;
        RECT 2401.360 82.870 2401.500 108.470 ;
        RECT 2401.360 82.730 2402.880 82.870 ;
        RECT 2402.740 2.400 2402.880 82.730 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.750 108.360 947.070 108.420 ;
        RECT 2415.070 108.360 2415.390 108.420 ;
        RECT 946.750 108.220 2415.390 108.360 ;
        RECT 946.750 108.160 947.070 108.220 ;
        RECT 2415.070 108.160 2415.390 108.220 ;
      LAYER via ;
        RECT 946.780 108.160 947.040 108.420 ;
        RECT 2415.100 108.160 2415.360 108.420 ;
      LAYER met2 ;
        RECT 945.750 400.250 946.030 404.000 ;
        RECT 945.750 400.110 947.440 400.250 ;
        RECT 945.750 400.000 946.030 400.110 ;
        RECT 947.300 351.970 947.440 400.110 ;
        RECT 947.300 351.830 947.900 351.970 ;
        RECT 947.760 324.370 947.900 351.830 ;
        RECT 946.840 324.230 947.900 324.370 ;
        RECT 946.840 108.450 946.980 324.230 ;
        RECT 946.780 108.130 947.040 108.450 ;
        RECT 2415.100 108.130 2415.360 108.450 ;
        RECT 2415.160 82.870 2415.300 108.130 ;
        RECT 2415.160 82.730 2420.360 82.870 ;
        RECT 2420.220 2.400 2420.360 82.730 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.290 376.280 946.610 376.340 ;
        RECT 949.970 376.280 950.290 376.340 ;
        RECT 946.290 376.140 950.290 376.280 ;
        RECT 946.290 376.080 946.610 376.140 ;
        RECT 949.970 376.080 950.290 376.140 ;
        RECT 946.290 108.020 946.610 108.080 ;
        RECT 2435.770 108.020 2436.090 108.080 ;
        RECT 946.290 107.880 2436.090 108.020 ;
        RECT 946.290 107.820 946.610 107.880 ;
        RECT 2435.770 107.820 2436.090 107.880 ;
      LAYER via ;
        RECT 946.320 376.080 946.580 376.340 ;
        RECT 950.000 376.080 950.260 376.340 ;
        RECT 946.320 107.820 946.580 108.080 ;
        RECT 2435.800 107.820 2436.060 108.080 ;
      LAYER met2 ;
        RECT 951.270 400.250 951.550 404.000 ;
        RECT 950.060 400.110 951.550 400.250 ;
        RECT 950.060 376.370 950.200 400.110 ;
        RECT 951.270 400.000 951.550 400.110 ;
        RECT 946.320 376.050 946.580 376.370 ;
        RECT 950.000 376.050 950.260 376.370 ;
        RECT 946.380 108.110 946.520 376.050 ;
        RECT 946.320 107.790 946.580 108.110 ;
        RECT 2435.800 107.790 2436.060 108.110 ;
        RECT 2435.860 1.770 2436.000 107.790 ;
        RECT 2437.950 1.770 2438.510 2.400 ;
        RECT 2435.860 1.630 2438.510 1.770 ;
        RECT 2437.950 -4.800 2438.510 1.630 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 953.650 107.680 953.970 107.740 ;
        RECT 2449.570 107.680 2449.890 107.740 ;
        RECT 953.650 107.540 2449.890 107.680 ;
        RECT 953.650 107.480 953.970 107.540 ;
        RECT 2449.570 107.480 2449.890 107.540 ;
        RECT 2449.570 17.580 2449.890 17.640 ;
        RECT 2453.710 17.580 2454.030 17.640 ;
        RECT 2449.570 17.440 2454.030 17.580 ;
        RECT 2449.570 17.380 2449.890 17.440 ;
        RECT 2453.710 17.380 2454.030 17.440 ;
      LAYER via ;
        RECT 953.680 107.480 953.940 107.740 ;
        RECT 2449.600 107.480 2449.860 107.740 ;
        RECT 2449.600 17.380 2449.860 17.640 ;
        RECT 2453.740 17.380 2454.000 17.640 ;
      LAYER met2 ;
        RECT 956.790 400.250 957.070 404.000 ;
        RECT 955.580 400.110 957.070 400.250 ;
        RECT 955.580 324.370 955.720 400.110 ;
        RECT 956.790 400.000 957.070 400.110 ;
        RECT 953.740 324.230 955.720 324.370 ;
        RECT 953.740 107.770 953.880 324.230 ;
        RECT 953.680 107.450 953.940 107.770 ;
        RECT 2449.600 107.450 2449.860 107.770 ;
        RECT 2449.660 17.670 2449.800 107.450 ;
        RECT 2449.600 17.350 2449.860 17.670 ;
        RECT 2453.740 17.350 2454.000 17.670 ;
        RECT 2453.800 1.770 2453.940 17.350 ;
        RECT 2455.430 1.770 2455.990 2.400 ;
        RECT 2453.800 1.630 2455.990 1.770 ;
        RECT 2455.430 -4.800 2455.990 1.630 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.550 107.340 960.870 107.400 ;
        RECT 2470.270 107.340 2470.590 107.400 ;
        RECT 960.550 107.200 2470.590 107.340 ;
        RECT 960.550 107.140 960.870 107.200 ;
        RECT 2470.270 107.140 2470.590 107.200 ;
      LAYER via ;
        RECT 960.580 107.140 960.840 107.400 ;
        RECT 2470.300 107.140 2470.560 107.400 ;
      LAYER met2 ;
        RECT 961.850 400.250 962.130 404.000 ;
        RECT 960.640 400.110 962.130 400.250 ;
        RECT 960.640 107.430 960.780 400.110 ;
        RECT 961.850 400.000 962.130 400.110 ;
        RECT 960.580 107.110 960.840 107.430 ;
        RECT 2470.300 107.110 2470.560 107.430 ;
        RECT 2470.360 82.870 2470.500 107.110 ;
        RECT 2470.360 82.730 2473.720 82.870 ;
        RECT 2473.580 2.400 2473.720 82.730 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.530 22.340 966.850 22.400 ;
        RECT 2490.970 22.340 2491.290 22.400 ;
        RECT 966.530 22.200 2491.290 22.340 ;
        RECT 966.530 22.140 966.850 22.200 ;
        RECT 2490.970 22.140 2491.290 22.200 ;
      LAYER via ;
        RECT 966.560 22.140 966.820 22.400 ;
        RECT 2491.000 22.140 2491.260 22.400 ;
      LAYER met2 ;
        RECT 967.370 400.250 967.650 404.000 ;
        RECT 966.160 400.110 967.650 400.250 ;
        RECT 966.160 34.570 966.300 400.110 ;
        RECT 967.370 400.000 967.650 400.110 ;
        RECT 966.160 34.430 966.760 34.570 ;
        RECT 966.620 22.430 966.760 34.430 ;
        RECT 966.560 22.110 966.820 22.430 ;
        RECT 2491.000 22.110 2491.260 22.430 ;
        RECT 2491.060 2.400 2491.200 22.110 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.430 22.680 973.750 22.740 ;
        RECT 2508.910 22.680 2509.230 22.740 ;
        RECT 973.430 22.540 2509.230 22.680 ;
        RECT 973.430 22.480 973.750 22.540 ;
        RECT 2508.910 22.480 2509.230 22.540 ;
      LAYER via ;
        RECT 973.460 22.480 973.720 22.740 ;
        RECT 2508.940 22.480 2509.200 22.740 ;
      LAYER met2 ;
        RECT 972.890 400.250 973.170 404.000 ;
        RECT 972.890 400.110 973.660 400.250 ;
        RECT 972.890 400.000 973.170 400.110 ;
        RECT 973.520 22.770 973.660 400.110 ;
        RECT 973.460 22.450 973.720 22.770 ;
        RECT 2508.940 22.450 2509.200 22.770 ;
        RECT 2509.000 2.400 2509.140 22.450 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.970 376.280 973.290 376.340 ;
        RECT 977.110 376.280 977.430 376.340 ;
        RECT 972.970 376.140 977.430 376.280 ;
        RECT 972.970 376.080 973.290 376.140 ;
        RECT 977.110 376.080 977.430 376.140 ;
        RECT 972.970 23.020 973.290 23.080 ;
        RECT 2526.850 23.020 2527.170 23.080 ;
        RECT 972.970 22.880 2527.170 23.020 ;
        RECT 972.970 22.820 973.290 22.880 ;
        RECT 2526.850 22.820 2527.170 22.880 ;
      LAYER via ;
        RECT 973.000 376.080 973.260 376.340 ;
        RECT 977.140 376.080 977.400 376.340 ;
        RECT 973.000 22.820 973.260 23.080 ;
        RECT 2526.880 22.820 2527.140 23.080 ;
      LAYER met2 ;
        RECT 978.410 400.250 978.690 404.000 ;
        RECT 977.200 400.110 978.690 400.250 ;
        RECT 977.200 376.370 977.340 400.110 ;
        RECT 978.410 400.000 978.690 400.110 ;
        RECT 973.000 376.050 973.260 376.370 ;
        RECT 977.140 376.050 977.400 376.370 ;
        RECT 973.060 23.110 973.200 376.050 ;
        RECT 973.000 22.790 973.260 23.110 ;
        RECT 2526.880 22.790 2527.140 23.110 ;
        RECT 2526.940 2.400 2527.080 22.790 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 979.870 375.940 980.190 376.000 ;
        RECT 982.630 375.940 982.950 376.000 ;
        RECT 979.870 375.800 982.950 375.940 ;
        RECT 979.870 375.740 980.190 375.800 ;
        RECT 982.630 375.740 982.950 375.800 ;
        RECT 979.870 23.360 980.190 23.420 ;
        RECT 2544.330 23.360 2544.650 23.420 ;
        RECT 979.870 23.220 2544.650 23.360 ;
        RECT 979.870 23.160 980.190 23.220 ;
        RECT 2544.330 23.160 2544.650 23.220 ;
      LAYER via ;
        RECT 979.900 375.740 980.160 376.000 ;
        RECT 982.660 375.740 982.920 376.000 ;
        RECT 979.900 23.160 980.160 23.420 ;
        RECT 2544.360 23.160 2544.620 23.420 ;
      LAYER met2 ;
        RECT 983.930 400.250 984.210 404.000 ;
        RECT 982.720 400.110 984.210 400.250 ;
        RECT 982.720 376.030 982.860 400.110 ;
        RECT 983.930 400.000 984.210 400.110 ;
        RECT 979.900 375.710 980.160 376.030 ;
        RECT 982.660 375.710 982.920 376.030 ;
        RECT 979.960 23.450 980.100 375.710 ;
        RECT 979.900 23.130 980.160 23.450 ;
        RECT 2544.360 23.130 2544.620 23.450 ;
        RECT 2544.420 2.400 2544.560 23.130 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 986.770 376.280 987.090 376.340 ;
        RECT 988.150 376.280 988.470 376.340 ;
        RECT 986.770 376.140 988.470 376.280 ;
        RECT 986.770 376.080 987.090 376.140 ;
        RECT 988.150 376.080 988.470 376.140 ;
        RECT 986.770 23.700 987.090 23.760 ;
        RECT 2562.270 23.700 2562.590 23.760 ;
        RECT 986.770 23.560 2562.590 23.700 ;
        RECT 986.770 23.500 987.090 23.560 ;
        RECT 2562.270 23.500 2562.590 23.560 ;
      LAYER via ;
        RECT 986.800 376.080 987.060 376.340 ;
        RECT 988.180 376.080 988.440 376.340 ;
        RECT 986.800 23.500 987.060 23.760 ;
        RECT 2562.300 23.500 2562.560 23.760 ;
      LAYER met2 ;
        RECT 989.450 400.250 989.730 404.000 ;
        RECT 988.240 400.110 989.730 400.250 ;
        RECT 988.240 376.370 988.380 400.110 ;
        RECT 989.450 400.000 989.730 400.110 ;
        RECT 986.800 376.050 987.060 376.370 ;
        RECT 988.180 376.050 988.440 376.370 ;
        RECT 986.860 23.790 987.000 376.050 ;
        RECT 986.800 23.470 987.060 23.790 ;
        RECT 2562.300 23.470 2562.560 23.790 ;
        RECT 2562.360 2.400 2562.500 23.470 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.130 376.280 442.450 376.340 ;
        RECT 446.730 376.280 447.050 376.340 ;
        RECT 442.130 376.140 447.050 376.280 ;
        RECT 442.130 376.080 442.450 376.140 ;
        RECT 446.730 376.080 447.050 376.140 ;
        RECT 442.130 32.880 442.450 32.940 ;
        RECT 586.110 32.880 586.430 32.940 ;
        RECT 442.130 32.740 586.430 32.880 ;
        RECT 442.130 32.680 442.450 32.740 ;
        RECT 586.110 32.680 586.430 32.740 ;
        RECT 586.110 19.280 586.430 19.340 ;
        RECT 806.450 19.280 806.770 19.340 ;
        RECT 586.110 19.140 806.770 19.280 ;
        RECT 586.110 19.080 586.430 19.140 ;
        RECT 806.450 19.080 806.770 19.140 ;
      LAYER via ;
        RECT 442.160 376.080 442.420 376.340 ;
        RECT 446.760 376.080 447.020 376.340 ;
        RECT 442.160 32.680 442.420 32.940 ;
        RECT 586.140 32.680 586.400 32.940 ;
        RECT 586.140 19.080 586.400 19.340 ;
        RECT 806.480 19.080 806.740 19.340 ;
      LAYER met2 ;
        RECT 448.030 400.250 448.310 404.000 ;
        RECT 446.820 400.110 448.310 400.250 ;
        RECT 446.820 376.370 446.960 400.110 ;
        RECT 448.030 400.000 448.310 400.110 ;
        RECT 442.160 376.050 442.420 376.370 ;
        RECT 446.760 376.050 447.020 376.370 ;
        RECT 442.220 32.970 442.360 376.050 ;
        RECT 442.160 32.650 442.420 32.970 ;
        RECT 586.140 32.650 586.400 32.970 ;
        RECT 586.200 19.370 586.340 32.650 ;
        RECT 586.140 19.050 586.400 19.370 ;
        RECT 806.480 19.050 806.740 19.370 ;
        RECT 806.540 2.400 806.680 19.050 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 993.670 27.440 993.990 27.500 ;
        RECT 2579.750 27.440 2580.070 27.500 ;
        RECT 993.670 27.300 2580.070 27.440 ;
        RECT 993.670 27.240 993.990 27.300 ;
        RECT 2579.750 27.240 2580.070 27.300 ;
      LAYER via ;
        RECT 993.700 27.240 993.960 27.500 ;
        RECT 2579.780 27.240 2580.040 27.500 ;
      LAYER met2 ;
        RECT 994.970 400.250 995.250 404.000 ;
        RECT 993.760 400.110 995.250 400.250 ;
        RECT 993.760 27.530 993.900 400.110 ;
        RECT 994.970 400.000 995.250 400.110 ;
        RECT 993.700 27.210 993.960 27.530 ;
        RECT 2579.780 27.210 2580.040 27.530 ;
        RECT 2579.840 2.400 2579.980 27.210 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.570 27.100 1000.890 27.160 ;
        RECT 2597.690 27.100 2598.010 27.160 ;
        RECT 1000.570 26.960 2598.010 27.100 ;
        RECT 1000.570 26.900 1000.890 26.960 ;
        RECT 2597.690 26.900 2598.010 26.960 ;
      LAYER via ;
        RECT 1000.600 26.900 1000.860 27.160 ;
        RECT 2597.720 26.900 2597.980 27.160 ;
      LAYER met2 ;
        RECT 1000.490 400.180 1000.770 404.000 ;
        RECT 1000.490 400.000 1000.800 400.180 ;
        RECT 1000.660 27.190 1000.800 400.000 ;
        RECT 1000.600 26.870 1000.860 27.190 ;
        RECT 2597.720 26.870 2597.980 27.190 ;
        RECT 2597.780 2.400 2597.920 26.870 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.030 376.280 1001.350 376.340 ;
        RECT 1004.710 376.280 1005.030 376.340 ;
        RECT 1001.030 376.140 1005.030 376.280 ;
        RECT 1001.030 376.080 1001.350 376.140 ;
        RECT 1004.710 376.080 1005.030 376.140 ;
        RECT 1001.030 26.760 1001.350 26.820 ;
        RECT 2615.170 26.760 2615.490 26.820 ;
        RECT 1001.030 26.620 2615.490 26.760 ;
        RECT 1001.030 26.560 1001.350 26.620 ;
        RECT 2615.170 26.560 2615.490 26.620 ;
      LAYER via ;
        RECT 1001.060 376.080 1001.320 376.340 ;
        RECT 1004.740 376.080 1005.000 376.340 ;
        RECT 1001.060 26.560 1001.320 26.820 ;
        RECT 2615.200 26.560 2615.460 26.820 ;
      LAYER met2 ;
        RECT 1006.010 400.250 1006.290 404.000 ;
        RECT 1004.800 400.110 1006.290 400.250 ;
        RECT 1004.800 376.370 1004.940 400.110 ;
        RECT 1006.010 400.000 1006.290 400.110 ;
        RECT 1001.060 376.050 1001.320 376.370 ;
        RECT 1004.740 376.050 1005.000 376.370 ;
        RECT 1001.120 26.850 1001.260 376.050 ;
        RECT 1001.060 26.530 1001.320 26.850 ;
        RECT 2615.200 26.530 2615.460 26.850 ;
        RECT 2615.260 2.400 2615.400 26.530 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.470 375.940 1007.790 376.000 ;
        RECT 1009.770 375.940 1010.090 376.000 ;
        RECT 1007.470 375.800 1010.090 375.940 ;
        RECT 1007.470 375.740 1007.790 375.800 ;
        RECT 1009.770 375.740 1010.090 375.800 ;
        RECT 1007.470 26.420 1007.790 26.480 ;
        RECT 2633.110 26.420 2633.430 26.480 ;
        RECT 1007.470 26.280 2633.430 26.420 ;
        RECT 1007.470 26.220 1007.790 26.280 ;
        RECT 2633.110 26.220 2633.430 26.280 ;
      LAYER via ;
        RECT 1007.500 375.740 1007.760 376.000 ;
        RECT 1009.800 375.740 1010.060 376.000 ;
        RECT 1007.500 26.220 1007.760 26.480 ;
        RECT 2633.140 26.220 2633.400 26.480 ;
      LAYER met2 ;
        RECT 1011.070 400.250 1011.350 404.000 ;
        RECT 1009.860 400.110 1011.350 400.250 ;
        RECT 1009.860 376.030 1010.000 400.110 ;
        RECT 1011.070 400.000 1011.350 400.110 ;
        RECT 1007.500 375.710 1007.760 376.030 ;
        RECT 1009.800 375.710 1010.060 376.030 ;
        RECT 1007.560 26.510 1007.700 375.710 ;
        RECT 1007.500 26.190 1007.760 26.510 ;
        RECT 2633.140 26.190 2633.400 26.510 ;
        RECT 2633.200 2.400 2633.340 26.190 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.370 399.740 1014.690 399.800 ;
        RECT 1015.290 399.740 1015.610 399.800 ;
        RECT 1014.370 399.600 1015.610 399.740 ;
        RECT 1014.370 399.540 1014.690 399.600 ;
        RECT 1015.290 399.540 1015.610 399.600 ;
        RECT 1014.370 26.080 1014.690 26.140 ;
        RECT 2650.590 26.080 2650.910 26.140 ;
        RECT 1014.370 25.940 2650.910 26.080 ;
        RECT 1014.370 25.880 1014.690 25.940 ;
        RECT 2650.590 25.880 2650.910 25.940 ;
      LAYER via ;
        RECT 1014.400 399.540 1014.660 399.800 ;
        RECT 1015.320 399.540 1015.580 399.800 ;
        RECT 1014.400 25.880 1014.660 26.140 ;
        RECT 2650.620 25.880 2650.880 26.140 ;
      LAYER met2 ;
        RECT 1016.590 400.250 1016.870 404.000 ;
        RECT 1015.380 400.110 1016.870 400.250 ;
        RECT 1015.380 399.830 1015.520 400.110 ;
        RECT 1016.590 400.000 1016.870 400.110 ;
        RECT 1014.400 399.510 1014.660 399.830 ;
        RECT 1015.320 399.510 1015.580 399.830 ;
        RECT 1014.460 26.170 1014.600 399.510 ;
        RECT 1014.400 25.850 1014.660 26.170 ;
        RECT 2650.620 25.850 2650.880 26.170 ;
        RECT 2650.680 2.400 2650.820 25.850 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.730 25.740 1022.050 25.800 ;
        RECT 2668.530 25.740 2668.850 25.800 ;
        RECT 1021.730 25.600 2668.850 25.740 ;
        RECT 1021.730 25.540 1022.050 25.600 ;
        RECT 2668.530 25.540 2668.850 25.600 ;
      LAYER via ;
        RECT 1021.760 25.540 1022.020 25.800 ;
        RECT 2668.560 25.540 2668.820 25.800 ;
      LAYER met2 ;
        RECT 1022.110 400.250 1022.390 404.000 ;
        RECT 1021.820 400.110 1022.390 400.250 ;
        RECT 1021.820 25.830 1021.960 400.110 ;
        RECT 1022.110 400.000 1022.390 400.110 ;
        RECT 1021.760 25.510 1022.020 25.830 ;
        RECT 2668.560 25.510 2668.820 25.830 ;
        RECT 2668.620 2.400 2668.760 25.510 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.270 376.280 1021.590 376.340 ;
        RECT 1026.330 376.280 1026.650 376.340 ;
        RECT 1021.270 376.140 1026.650 376.280 ;
        RECT 1021.270 376.080 1021.590 376.140 ;
        RECT 1026.330 376.080 1026.650 376.140 ;
        RECT 1021.270 25.400 1021.590 25.460 ;
        RECT 2686.010 25.400 2686.330 25.460 ;
        RECT 1021.270 25.260 2686.330 25.400 ;
        RECT 1021.270 25.200 1021.590 25.260 ;
        RECT 2686.010 25.200 2686.330 25.260 ;
      LAYER via ;
        RECT 1021.300 376.080 1021.560 376.340 ;
        RECT 1026.360 376.080 1026.620 376.340 ;
        RECT 1021.300 25.200 1021.560 25.460 ;
        RECT 2686.040 25.200 2686.300 25.460 ;
      LAYER met2 ;
        RECT 1027.630 400.250 1027.910 404.000 ;
        RECT 1026.420 400.110 1027.910 400.250 ;
        RECT 1026.420 376.370 1026.560 400.110 ;
        RECT 1027.630 400.000 1027.910 400.110 ;
        RECT 1021.300 376.050 1021.560 376.370 ;
        RECT 1026.360 376.050 1026.620 376.370 ;
        RECT 1021.360 25.490 1021.500 376.050 ;
        RECT 1021.300 25.170 1021.560 25.490 ;
        RECT 2686.040 25.170 2686.300 25.490 ;
        RECT 2686.100 2.400 2686.240 25.170 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.170 376.280 1028.490 376.340 ;
        RECT 1031.850 376.280 1032.170 376.340 ;
        RECT 1028.170 376.140 1032.170 376.280 ;
        RECT 1028.170 376.080 1028.490 376.140 ;
        RECT 1031.850 376.080 1032.170 376.140 ;
        RECT 1028.170 25.060 1028.490 25.120 ;
        RECT 2703.950 25.060 2704.270 25.120 ;
        RECT 1028.170 24.920 2704.270 25.060 ;
        RECT 1028.170 24.860 1028.490 24.920 ;
        RECT 2703.950 24.860 2704.270 24.920 ;
      LAYER via ;
        RECT 1028.200 376.080 1028.460 376.340 ;
        RECT 1031.880 376.080 1032.140 376.340 ;
        RECT 1028.200 24.860 1028.460 25.120 ;
        RECT 2703.980 24.860 2704.240 25.120 ;
      LAYER met2 ;
        RECT 1033.150 400.250 1033.430 404.000 ;
        RECT 1031.940 400.110 1033.430 400.250 ;
        RECT 1031.940 376.370 1032.080 400.110 ;
        RECT 1033.150 400.000 1033.430 400.110 ;
        RECT 1028.200 376.050 1028.460 376.370 ;
        RECT 1031.880 376.050 1032.140 376.370 ;
        RECT 1028.260 25.150 1028.400 376.050 ;
        RECT 1028.200 24.830 1028.460 25.150 ;
        RECT 2703.980 24.830 2704.240 25.150 ;
        RECT 2704.040 2.400 2704.180 24.830 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.070 375.940 1035.390 376.000 ;
        RECT 1037.370 375.940 1037.690 376.000 ;
        RECT 1035.070 375.800 1037.690 375.940 ;
        RECT 1035.070 375.740 1035.390 375.800 ;
        RECT 1037.370 375.740 1037.690 375.800 ;
        RECT 1035.070 24.720 1035.390 24.780 ;
        RECT 2721.890 24.720 2722.210 24.780 ;
        RECT 1035.070 24.580 2722.210 24.720 ;
        RECT 1035.070 24.520 1035.390 24.580 ;
        RECT 2721.890 24.520 2722.210 24.580 ;
      LAYER via ;
        RECT 1035.100 375.740 1035.360 376.000 ;
        RECT 1037.400 375.740 1037.660 376.000 ;
        RECT 1035.100 24.520 1035.360 24.780 ;
        RECT 2721.920 24.520 2722.180 24.780 ;
      LAYER met2 ;
        RECT 1038.670 400.250 1038.950 404.000 ;
        RECT 1037.460 400.110 1038.950 400.250 ;
        RECT 1037.460 376.030 1037.600 400.110 ;
        RECT 1038.670 400.000 1038.950 400.110 ;
        RECT 1035.100 375.710 1035.360 376.030 ;
        RECT 1037.400 375.710 1037.660 376.030 ;
        RECT 1035.160 24.810 1035.300 375.710 ;
        RECT 1035.100 24.490 1035.360 24.810 ;
        RECT 2721.920 24.490 2722.180 24.810 ;
        RECT 2721.980 2.400 2722.120 24.490 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.970 375.940 1042.290 376.000 ;
        RECT 1044.270 375.940 1044.590 376.000 ;
        RECT 1041.970 375.800 1044.590 375.940 ;
        RECT 1041.970 375.740 1042.290 375.800 ;
        RECT 1044.270 375.740 1044.590 375.800 ;
        RECT 1041.970 24.380 1042.290 24.440 ;
        RECT 2739.370 24.380 2739.690 24.440 ;
        RECT 1041.970 24.240 2739.690 24.380 ;
        RECT 1041.970 24.180 1042.290 24.240 ;
        RECT 2739.370 24.180 2739.690 24.240 ;
      LAYER via ;
        RECT 1042.000 375.740 1042.260 376.000 ;
        RECT 1044.300 375.740 1044.560 376.000 ;
        RECT 1042.000 24.180 1042.260 24.440 ;
        RECT 2739.400 24.180 2739.660 24.440 ;
      LAYER met2 ;
        RECT 1044.190 400.180 1044.470 404.000 ;
        RECT 1044.190 400.000 1044.500 400.180 ;
        RECT 1044.360 376.030 1044.500 400.000 ;
        RECT 1042.000 375.710 1042.260 376.030 ;
        RECT 1044.300 375.710 1044.560 376.030 ;
        RECT 1042.060 24.470 1042.200 375.710 ;
        RECT 1042.000 24.150 1042.260 24.470 ;
        RECT 2739.400 24.150 2739.660 24.470 ;
        RECT 2739.460 2.400 2739.600 24.150 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 453.630 393.280 453.950 393.340 ;
        RECT 596.690 393.280 597.010 393.340 ;
        RECT 453.630 393.140 597.010 393.280 ;
        RECT 453.630 393.080 453.950 393.140 ;
        RECT 596.690 393.080 597.010 393.140 ;
        RECT 596.690 18.940 597.010 19.000 ;
        RECT 824.390 18.940 824.710 19.000 ;
        RECT 596.690 18.800 824.710 18.940 ;
        RECT 596.690 18.740 597.010 18.800 ;
        RECT 824.390 18.740 824.710 18.800 ;
      LAYER via ;
        RECT 453.660 393.080 453.920 393.340 ;
        RECT 596.720 393.080 596.980 393.340 ;
        RECT 596.720 18.740 596.980 19.000 ;
        RECT 824.420 18.740 824.680 19.000 ;
      LAYER met2 ;
        RECT 453.550 400.180 453.830 404.000 ;
        RECT 453.550 400.000 453.860 400.180 ;
        RECT 453.720 393.370 453.860 400.000 ;
        RECT 453.660 393.050 453.920 393.370 ;
        RECT 596.720 393.050 596.980 393.370 ;
        RECT 596.780 19.030 596.920 393.050 ;
        RECT 596.720 18.710 596.980 19.030 ;
        RECT 824.420 18.710 824.680 19.030 ;
        RECT 824.480 2.400 824.620 18.710 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.330 24.040 1049.650 24.100 ;
        RECT 2757.310 24.040 2757.630 24.100 ;
        RECT 1049.330 23.900 2757.630 24.040 ;
        RECT 1049.330 23.840 1049.650 23.900 ;
        RECT 2757.310 23.840 2757.630 23.900 ;
      LAYER via ;
        RECT 1049.360 23.840 1049.620 24.100 ;
        RECT 2757.340 23.840 2757.600 24.100 ;
      LAYER met2 ;
        RECT 1049.710 400.250 1049.990 404.000 ;
        RECT 1049.420 400.110 1049.990 400.250 ;
        RECT 1049.420 24.130 1049.560 400.110 ;
        RECT 1049.710 400.000 1049.990 400.110 ;
        RECT 1049.360 23.810 1049.620 24.130 ;
        RECT 2757.340 23.810 2757.600 24.130 ;
        RECT 2757.400 2.400 2757.540 23.810 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.770 400.250 1055.050 404.000 ;
        RECT 1054.020 400.110 1055.050 400.250 ;
        RECT 1054.020 324.370 1054.160 400.110 ;
        RECT 1054.770 400.000 1055.050 400.110 ;
        RECT 1050.800 324.230 1054.160 324.370 ;
        RECT 1050.800 24.325 1050.940 324.230 ;
        RECT 1050.730 23.955 1051.010 24.325 ;
        RECT 2774.810 23.955 2775.090 24.325 ;
        RECT 2774.880 2.400 2775.020 23.955 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
      LAYER via2 ;
        RECT 1050.730 24.000 1051.010 24.280 ;
        RECT 2774.810 24.000 2775.090 24.280 ;
      LAYER met3 ;
        RECT 1050.705 24.290 1051.035 24.305 ;
        RECT 2774.785 24.290 2775.115 24.305 ;
        RECT 1050.705 23.990 2775.115 24.290 ;
        RECT 1050.705 23.975 1051.035 23.990 ;
        RECT 2774.785 23.975 2775.115 23.990 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1057.150 107.000 1057.470 107.060 ;
        RECT 2787.670 107.000 2787.990 107.060 ;
        RECT 1057.150 106.860 2787.990 107.000 ;
        RECT 1057.150 106.800 1057.470 106.860 ;
        RECT 2787.670 106.800 2787.990 106.860 ;
      LAYER via ;
        RECT 1057.180 106.800 1057.440 107.060 ;
        RECT 2787.700 106.800 2787.960 107.060 ;
      LAYER met2 ;
        RECT 1060.290 400.250 1060.570 404.000 ;
        RECT 1059.080 400.110 1060.570 400.250 ;
        RECT 1059.080 324.370 1059.220 400.110 ;
        RECT 1060.290 400.000 1060.570 400.110 ;
        RECT 1057.240 324.230 1059.220 324.370 ;
        RECT 1057.240 107.090 1057.380 324.230 ;
        RECT 1057.180 106.770 1057.440 107.090 ;
        RECT 2787.700 106.770 2787.960 107.090 ;
        RECT 2787.760 82.870 2787.900 106.770 ;
        RECT 2787.760 82.730 2792.960 82.870 ;
        RECT 2792.820 2.400 2792.960 82.730 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.810 400.250 1066.090 404.000 ;
        RECT 1064.600 400.110 1066.090 400.250 ;
        RECT 1064.600 324.370 1064.740 400.110 ;
        RECT 1065.810 400.000 1066.090 400.110 ;
        RECT 1063.680 324.230 1064.740 324.370 ;
        RECT 1063.680 107.285 1063.820 324.230 ;
        RECT 1063.610 106.915 1063.890 107.285 ;
        RECT 2808.390 106.915 2808.670 107.285 ;
        RECT 2808.460 82.870 2808.600 106.915 ;
        RECT 2808.460 82.730 2810.440 82.870 ;
        RECT 2810.300 2.400 2810.440 82.730 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
      LAYER via2 ;
        RECT 1063.610 106.960 1063.890 107.240 ;
        RECT 2808.390 106.960 2808.670 107.240 ;
      LAYER met3 ;
        RECT 1063.585 107.250 1063.915 107.265 ;
        RECT 2808.365 107.250 2808.695 107.265 ;
        RECT 1063.585 106.950 2808.695 107.250 ;
        RECT 1063.585 106.935 1063.915 106.950 ;
        RECT 2808.365 106.935 2808.695 106.950 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2822.170 17.580 2822.490 17.640 ;
        RECT 2826.310 17.580 2826.630 17.640 ;
        RECT 2822.170 17.440 2826.630 17.580 ;
        RECT 2822.170 17.380 2822.490 17.440 ;
        RECT 2826.310 17.380 2826.630 17.440 ;
      LAYER via ;
        RECT 2822.200 17.380 2822.460 17.640 ;
        RECT 2826.340 17.380 2826.600 17.640 ;
      LAYER met2 ;
        RECT 1071.330 400.250 1071.610 404.000 ;
        RECT 1071.040 400.110 1071.610 400.250 ;
        RECT 1071.040 106.605 1071.180 400.110 ;
        RECT 1071.330 400.000 1071.610 400.110 ;
        RECT 1070.970 106.235 1071.250 106.605 ;
        RECT 2822.190 106.235 2822.470 106.605 ;
        RECT 2822.260 17.670 2822.400 106.235 ;
        RECT 2822.200 17.350 2822.460 17.670 ;
        RECT 2826.340 17.350 2826.600 17.670 ;
        RECT 2826.400 1.770 2826.540 17.350 ;
        RECT 2828.030 1.770 2828.590 2.400 ;
        RECT 2826.400 1.630 2828.590 1.770 ;
        RECT 2828.030 -4.800 2828.590 1.630 ;
      LAYER via2 ;
        RECT 1070.970 106.280 1071.250 106.560 ;
        RECT 2822.190 106.280 2822.470 106.560 ;
      LAYER met3 ;
        RECT 1070.945 106.570 1071.275 106.585 ;
        RECT 2822.165 106.570 2822.495 106.585 ;
        RECT 1070.945 106.270 2822.495 106.570 ;
        RECT 1070.945 106.255 1071.275 106.270 ;
        RECT 2822.165 106.255 2822.495 106.270 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.930 31.860 1077.250 31.920 ;
        RECT 2845.630 31.860 2845.950 31.920 ;
        RECT 1076.930 31.720 2845.950 31.860 ;
        RECT 1076.930 31.660 1077.250 31.720 ;
        RECT 2845.630 31.660 2845.950 31.720 ;
      LAYER via ;
        RECT 1076.960 31.660 1077.220 31.920 ;
        RECT 2845.660 31.660 2845.920 31.920 ;
      LAYER met2 ;
        RECT 1076.850 400.180 1077.130 404.000 ;
        RECT 1076.850 400.000 1077.160 400.180 ;
        RECT 1077.020 31.950 1077.160 400.000 ;
        RECT 1076.960 31.630 1077.220 31.950 ;
        RECT 2845.660 31.630 2845.920 31.950 ;
        RECT 2845.720 2.400 2845.860 31.630 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.470 386.480 1076.790 386.540 ;
        RECT 1081.070 386.480 1081.390 386.540 ;
        RECT 1076.470 386.340 1081.390 386.480 ;
        RECT 1076.470 386.280 1076.790 386.340 ;
        RECT 1081.070 386.280 1081.390 386.340 ;
        RECT 1076.470 31.520 1076.790 31.580 ;
        RECT 2863.570 31.520 2863.890 31.580 ;
        RECT 1076.470 31.380 2863.890 31.520 ;
        RECT 1076.470 31.320 1076.790 31.380 ;
        RECT 2863.570 31.320 2863.890 31.380 ;
      LAYER via ;
        RECT 1076.500 386.280 1076.760 386.540 ;
        RECT 1081.100 386.280 1081.360 386.540 ;
        RECT 1076.500 31.320 1076.760 31.580 ;
        RECT 2863.600 31.320 2863.860 31.580 ;
      LAYER met2 ;
        RECT 1082.370 400.250 1082.650 404.000 ;
        RECT 1081.160 400.110 1082.650 400.250 ;
        RECT 1081.160 386.570 1081.300 400.110 ;
        RECT 1082.370 400.000 1082.650 400.110 ;
        RECT 1076.500 386.250 1076.760 386.570 ;
        RECT 1081.100 386.250 1081.360 386.570 ;
        RECT 1076.560 31.610 1076.700 386.250 ;
        RECT 1076.500 31.290 1076.760 31.610 ;
        RECT 2863.600 31.290 2863.860 31.610 ;
        RECT 2863.660 2.400 2863.800 31.290 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1083.370 386.140 1083.690 386.200 ;
        RECT 1086.590 386.140 1086.910 386.200 ;
        RECT 1083.370 386.000 1086.910 386.140 ;
        RECT 1083.370 385.940 1083.690 386.000 ;
        RECT 1086.590 385.940 1086.910 386.000 ;
        RECT 1083.370 31.180 1083.690 31.240 ;
        RECT 2881.510 31.180 2881.830 31.240 ;
        RECT 1083.370 31.040 2881.830 31.180 ;
        RECT 1083.370 30.980 1083.690 31.040 ;
        RECT 2881.510 30.980 2881.830 31.040 ;
      LAYER via ;
        RECT 1083.400 385.940 1083.660 386.200 ;
        RECT 1086.620 385.940 1086.880 386.200 ;
        RECT 1083.400 30.980 1083.660 31.240 ;
        RECT 2881.540 30.980 2881.800 31.240 ;
      LAYER met2 ;
        RECT 1087.890 400.250 1088.170 404.000 ;
        RECT 1086.680 400.110 1088.170 400.250 ;
        RECT 1086.680 386.230 1086.820 400.110 ;
        RECT 1087.890 400.000 1088.170 400.110 ;
        RECT 1083.400 385.910 1083.660 386.230 ;
        RECT 1086.620 385.910 1086.880 386.230 ;
        RECT 1083.460 31.270 1083.600 385.910 ;
        RECT 1083.400 30.950 1083.660 31.270 ;
        RECT 2881.540 30.950 2881.800 31.270 ;
        RECT 2881.600 2.400 2881.740 30.950 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 459.150 389.200 459.470 389.260 ;
        RECT 598.530 389.200 598.850 389.260 ;
        RECT 459.150 389.060 598.850 389.200 ;
        RECT 459.150 389.000 459.470 389.060 ;
        RECT 598.530 389.000 598.850 389.060 ;
        RECT 597.610 18.600 597.930 18.660 ;
        RECT 841.870 18.600 842.190 18.660 ;
        RECT 597.610 18.460 842.190 18.600 ;
        RECT 597.610 18.400 597.930 18.460 ;
        RECT 841.870 18.400 842.190 18.460 ;
      LAYER via ;
        RECT 459.180 389.000 459.440 389.260 ;
        RECT 598.560 389.000 598.820 389.260 ;
        RECT 597.640 18.400 597.900 18.660 ;
        RECT 841.900 18.400 842.160 18.660 ;
      LAYER met2 ;
        RECT 459.070 400.180 459.350 404.000 ;
        RECT 459.070 400.000 459.380 400.180 ;
        RECT 459.240 389.290 459.380 400.000 ;
        RECT 459.180 388.970 459.440 389.290 ;
        RECT 598.560 388.970 598.820 389.290 ;
        RECT 598.620 324.370 598.760 388.970 ;
        RECT 597.700 324.230 598.760 324.370 ;
        RECT 597.700 18.690 597.840 324.230 ;
        RECT 597.640 18.370 597.900 18.690 ;
        RECT 841.900 18.370 842.160 18.690 ;
        RECT 841.960 2.400 842.100 18.370 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.670 387.840 464.990 387.900 ;
        RECT 597.150 387.840 597.470 387.900 ;
        RECT 464.670 387.700 597.470 387.840 ;
        RECT 464.670 387.640 464.990 387.700 ;
        RECT 597.150 387.640 597.470 387.700 ;
        RECT 597.150 18.260 597.470 18.320 ;
        RECT 859.810 18.260 860.130 18.320 ;
        RECT 597.150 18.120 860.130 18.260 ;
        RECT 597.150 18.060 597.470 18.120 ;
        RECT 859.810 18.060 860.130 18.120 ;
      LAYER via ;
        RECT 464.700 387.640 464.960 387.900 ;
        RECT 597.180 387.640 597.440 387.900 ;
        RECT 597.180 18.060 597.440 18.320 ;
        RECT 859.840 18.060 860.100 18.320 ;
      LAYER met2 ;
        RECT 464.590 400.180 464.870 404.000 ;
        RECT 464.590 400.000 464.900 400.180 ;
        RECT 464.760 387.930 464.900 400.000 ;
        RECT 464.700 387.610 464.960 387.930 ;
        RECT 597.180 387.610 597.440 387.930 ;
        RECT 597.240 18.350 597.380 387.610 ;
        RECT 597.180 18.030 597.440 18.350 ;
        RECT 859.840 18.030 860.100 18.350 ;
        RECT 859.900 2.400 860.040 18.030 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.190 392.940 470.510 393.000 ;
        RECT 568.630 392.940 568.950 393.000 ;
        RECT 470.190 392.800 568.950 392.940 ;
        RECT 470.190 392.740 470.510 392.800 ;
        RECT 568.630 392.740 568.950 392.800 ;
        RECT 568.630 388.520 568.950 388.580 ;
        RECT 617.390 388.520 617.710 388.580 ;
        RECT 568.630 388.380 617.710 388.520 ;
        RECT 568.630 388.320 568.950 388.380 ;
        RECT 617.390 388.320 617.710 388.380 ;
        RECT 616.930 17.920 617.250 17.980 ;
        RECT 877.290 17.920 877.610 17.980 ;
        RECT 616.930 17.780 877.610 17.920 ;
        RECT 616.930 17.720 617.250 17.780 ;
        RECT 877.290 17.720 877.610 17.780 ;
      LAYER via ;
        RECT 470.220 392.740 470.480 393.000 ;
        RECT 568.660 392.740 568.920 393.000 ;
        RECT 568.660 388.320 568.920 388.580 ;
        RECT 617.420 388.320 617.680 388.580 ;
        RECT 616.960 17.720 617.220 17.980 ;
        RECT 877.320 17.720 877.580 17.980 ;
      LAYER met2 ;
        RECT 470.110 400.180 470.390 404.000 ;
        RECT 470.110 400.000 470.420 400.180 ;
        RECT 470.280 393.030 470.420 400.000 ;
        RECT 470.220 392.710 470.480 393.030 ;
        RECT 568.660 392.710 568.920 393.030 ;
        RECT 568.720 388.610 568.860 392.710 ;
        RECT 568.660 388.290 568.920 388.610 ;
        RECT 617.420 388.290 617.680 388.610 ;
        RECT 617.480 34.570 617.620 388.290 ;
        RECT 617.020 34.430 617.620 34.570 ;
        RECT 617.020 18.010 617.160 34.430 ;
        RECT 616.960 17.690 617.220 18.010 ;
        RECT 877.320 17.690 877.580 18.010 ;
        RECT 877.380 2.400 877.520 17.690 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 475.710 392.600 476.030 392.660 ;
        RECT 617.850 392.600 618.170 392.660 ;
        RECT 475.710 392.460 618.170 392.600 ;
        RECT 475.710 392.400 476.030 392.460 ;
        RECT 617.850 392.400 618.170 392.460 ;
        RECT 617.850 17.580 618.170 17.640 ;
        RECT 895.230 17.580 895.550 17.640 ;
        RECT 617.850 17.440 895.550 17.580 ;
        RECT 617.850 17.380 618.170 17.440 ;
        RECT 895.230 17.380 895.550 17.440 ;
      LAYER via ;
        RECT 475.740 392.400 476.000 392.660 ;
        RECT 617.880 392.400 618.140 392.660 ;
        RECT 617.880 17.380 618.140 17.640 ;
        RECT 895.260 17.380 895.520 17.640 ;
      LAYER met2 ;
        RECT 475.630 400.180 475.910 404.000 ;
        RECT 475.630 400.000 475.940 400.180 ;
        RECT 475.800 392.690 475.940 400.000 ;
        RECT 475.740 392.370 476.000 392.690 ;
        RECT 617.880 392.370 618.140 392.690 ;
        RECT 617.940 17.670 618.080 392.370 ;
        RECT 617.880 17.350 618.140 17.670 ;
        RECT 895.260 17.350 895.520 17.670 ;
        RECT 895.320 2.400 895.460 17.350 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 376.280 476.490 376.340 ;
        RECT 479.850 376.280 480.170 376.340 ;
        RECT 476.170 376.140 480.170 376.280 ;
        RECT 476.170 376.080 476.490 376.140 ;
        RECT 479.850 376.080 480.170 376.140 ;
        RECT 476.170 26.420 476.490 26.480 ;
        RECT 912.710 26.420 913.030 26.480 ;
        RECT 476.170 26.280 913.030 26.420 ;
        RECT 476.170 26.220 476.490 26.280 ;
        RECT 912.710 26.220 913.030 26.280 ;
      LAYER via ;
        RECT 476.200 376.080 476.460 376.340 ;
        RECT 479.880 376.080 480.140 376.340 ;
        RECT 476.200 26.220 476.460 26.480 ;
        RECT 912.740 26.220 913.000 26.480 ;
      LAYER met2 ;
        RECT 481.150 400.250 481.430 404.000 ;
        RECT 479.940 400.110 481.430 400.250 ;
        RECT 479.940 376.370 480.080 400.110 ;
        RECT 481.150 400.000 481.430 400.110 ;
        RECT 476.200 376.050 476.460 376.370 ;
        RECT 479.880 376.050 480.140 376.370 ;
        RECT 476.260 26.510 476.400 376.050 ;
        RECT 476.200 26.190 476.460 26.510 ;
        RECT 912.740 26.190 913.000 26.510 ;
        RECT 912.800 2.400 912.940 26.190 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 376.280 483.390 376.340 ;
        RECT 485.370 376.280 485.690 376.340 ;
        RECT 483.070 376.140 485.690 376.280 ;
        RECT 483.070 376.080 483.390 376.140 ;
        RECT 485.370 376.080 485.690 376.140 ;
        RECT 483.070 26.080 483.390 26.140 ;
        RECT 930.650 26.080 930.970 26.140 ;
        RECT 483.070 25.940 930.970 26.080 ;
        RECT 483.070 25.880 483.390 25.940 ;
        RECT 930.650 25.880 930.970 25.940 ;
      LAYER via ;
        RECT 483.100 376.080 483.360 376.340 ;
        RECT 485.400 376.080 485.660 376.340 ;
        RECT 483.100 25.880 483.360 26.140 ;
        RECT 930.680 25.880 930.940 26.140 ;
      LAYER met2 ;
        RECT 486.210 400.250 486.490 404.000 ;
        RECT 485.460 400.110 486.490 400.250 ;
        RECT 485.460 376.370 485.600 400.110 ;
        RECT 486.210 400.000 486.490 400.110 ;
        RECT 483.100 376.050 483.360 376.370 ;
        RECT 485.400 376.050 485.660 376.370 ;
        RECT 483.160 26.170 483.300 376.050 ;
        RECT 483.100 25.850 483.360 26.170 ;
        RECT 930.680 25.850 930.940 26.170 ;
        RECT 930.740 2.400 930.880 25.850 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 376.280 490.290 376.340 ;
        RECT 490.890 376.280 491.210 376.340 ;
        RECT 489.970 376.140 491.210 376.280 ;
        RECT 489.970 376.080 490.290 376.140 ;
        RECT 490.890 376.080 491.210 376.140 ;
        RECT 489.970 25.740 490.290 25.800 ;
        RECT 948.590 25.740 948.910 25.800 ;
        RECT 489.970 25.600 948.910 25.740 ;
        RECT 489.970 25.540 490.290 25.600 ;
        RECT 948.590 25.540 948.910 25.600 ;
      LAYER via ;
        RECT 490.000 376.080 490.260 376.340 ;
        RECT 490.920 376.080 491.180 376.340 ;
        RECT 490.000 25.540 490.260 25.800 ;
        RECT 948.620 25.540 948.880 25.800 ;
      LAYER met2 ;
        RECT 491.730 400.250 492.010 404.000 ;
        RECT 490.980 400.110 492.010 400.250 ;
        RECT 490.980 376.370 491.120 400.110 ;
        RECT 491.730 400.000 492.010 400.110 ;
        RECT 490.000 376.050 490.260 376.370 ;
        RECT 490.920 376.050 491.180 376.370 ;
        RECT 490.060 25.830 490.200 376.050 ;
        RECT 490.000 25.510 490.260 25.830 ;
        RECT 948.620 25.510 948.880 25.830 ;
        RECT 948.680 2.400 948.820 25.510 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 25.400 497.190 25.460 ;
        RECT 966.070 25.400 966.390 25.460 ;
        RECT 496.870 25.260 966.390 25.400 ;
        RECT 496.870 25.200 497.190 25.260 ;
        RECT 966.070 25.200 966.390 25.260 ;
      LAYER via ;
        RECT 496.900 25.200 497.160 25.460 ;
        RECT 966.100 25.200 966.360 25.460 ;
      LAYER met2 ;
        RECT 497.250 400.250 497.530 404.000 ;
        RECT 496.960 400.110 497.530 400.250 ;
        RECT 496.960 25.490 497.100 400.110 ;
        RECT 497.250 400.000 497.530 400.110 ;
        RECT 496.900 25.170 497.160 25.490 ;
        RECT 966.100 25.170 966.360 25.490 ;
        RECT 966.160 2.400 966.300 25.170 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.370 386.480 393.690 386.540 ;
        RECT 397.510 386.480 397.830 386.540 ;
        RECT 393.370 386.340 397.830 386.480 ;
        RECT 393.370 386.280 393.690 386.340 ;
        RECT 397.510 386.280 397.830 386.340 ;
        RECT 393.370 22.680 393.690 22.740 ;
        RECT 646.830 22.680 647.150 22.740 ;
        RECT 393.370 22.540 647.150 22.680 ;
        RECT 393.370 22.480 393.690 22.540 ;
        RECT 646.830 22.480 647.150 22.540 ;
      LAYER via ;
        RECT 393.400 386.280 393.660 386.540 ;
        RECT 397.540 386.280 397.800 386.540 ;
        RECT 393.400 22.480 393.660 22.740 ;
        RECT 646.860 22.480 647.120 22.740 ;
      LAYER met2 ;
        RECT 398.810 400.250 399.090 404.000 ;
        RECT 397.600 400.110 399.090 400.250 ;
        RECT 397.600 386.570 397.740 400.110 ;
        RECT 398.810 400.000 399.090 400.110 ;
        RECT 393.400 386.250 393.660 386.570 ;
        RECT 397.540 386.250 397.800 386.570 ;
        RECT 393.460 22.770 393.600 386.250 ;
        RECT 393.400 22.450 393.660 22.770 ;
        RECT 646.860 22.450 647.120 22.770 ;
        RECT 646.920 2.400 647.060 22.450 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 386.480 497.650 386.540 ;
        RECT 501.470 386.480 501.790 386.540 ;
        RECT 497.330 386.340 501.790 386.480 ;
        RECT 497.330 386.280 497.650 386.340 ;
        RECT 501.470 386.280 501.790 386.340 ;
        RECT 497.330 25.060 497.650 25.120 ;
        RECT 984.010 25.060 984.330 25.120 ;
        RECT 497.330 24.920 984.330 25.060 ;
        RECT 497.330 24.860 497.650 24.920 ;
        RECT 984.010 24.860 984.330 24.920 ;
      LAYER via ;
        RECT 497.360 386.280 497.620 386.540 ;
        RECT 501.500 386.280 501.760 386.540 ;
        RECT 497.360 24.860 497.620 25.120 ;
        RECT 984.040 24.860 984.300 25.120 ;
      LAYER met2 ;
        RECT 502.770 400.250 503.050 404.000 ;
        RECT 501.560 400.110 503.050 400.250 ;
        RECT 501.560 386.570 501.700 400.110 ;
        RECT 502.770 400.000 503.050 400.110 ;
        RECT 497.360 386.250 497.620 386.570 ;
        RECT 501.500 386.250 501.760 386.570 ;
        RECT 497.420 25.150 497.560 386.250 ;
        RECT 497.360 24.830 497.620 25.150 ;
        RECT 984.040 24.830 984.300 25.150 ;
        RECT 984.100 2.400 984.240 24.830 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 386.480 504.090 386.540 ;
        RECT 506.990 386.480 507.310 386.540 ;
        RECT 503.770 386.340 507.310 386.480 ;
        RECT 503.770 386.280 504.090 386.340 ;
        RECT 506.990 386.280 507.310 386.340 ;
        RECT 503.770 24.720 504.090 24.780 ;
        RECT 1001.490 24.720 1001.810 24.780 ;
        RECT 503.770 24.580 1001.810 24.720 ;
        RECT 503.770 24.520 504.090 24.580 ;
        RECT 1001.490 24.520 1001.810 24.580 ;
      LAYER via ;
        RECT 503.800 386.280 504.060 386.540 ;
        RECT 507.020 386.280 507.280 386.540 ;
        RECT 503.800 24.520 504.060 24.780 ;
        RECT 1001.520 24.520 1001.780 24.780 ;
      LAYER met2 ;
        RECT 508.290 400.250 508.570 404.000 ;
        RECT 507.080 400.110 508.570 400.250 ;
        RECT 507.080 386.570 507.220 400.110 ;
        RECT 508.290 400.000 508.570 400.110 ;
        RECT 503.800 386.250 504.060 386.570 ;
        RECT 507.020 386.250 507.280 386.570 ;
        RECT 503.860 24.810 504.000 386.250 ;
        RECT 503.800 24.490 504.060 24.810 ;
        RECT 1001.520 24.490 1001.780 24.810 ;
        RECT 1001.580 2.400 1001.720 24.490 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 386.480 510.990 386.540 ;
        RECT 512.510 386.480 512.830 386.540 ;
        RECT 510.670 386.340 512.830 386.480 ;
        RECT 510.670 386.280 510.990 386.340 ;
        RECT 512.510 386.280 512.830 386.340 ;
        RECT 510.670 24.380 510.990 24.440 ;
        RECT 1019.430 24.380 1019.750 24.440 ;
        RECT 510.670 24.240 1019.750 24.380 ;
        RECT 510.670 24.180 510.990 24.240 ;
        RECT 1019.430 24.180 1019.750 24.240 ;
      LAYER via ;
        RECT 510.700 386.280 510.960 386.540 ;
        RECT 512.540 386.280 512.800 386.540 ;
        RECT 510.700 24.180 510.960 24.440 ;
        RECT 1019.460 24.180 1019.720 24.440 ;
      LAYER met2 ;
        RECT 513.810 400.250 514.090 404.000 ;
        RECT 512.600 400.110 514.090 400.250 ;
        RECT 512.600 386.570 512.740 400.110 ;
        RECT 513.810 400.000 514.090 400.110 ;
        RECT 510.700 386.250 510.960 386.570 ;
        RECT 512.540 386.250 512.800 386.570 ;
        RECT 510.760 24.470 510.900 386.250 ;
        RECT 510.700 24.150 510.960 24.470 ;
        RECT 1019.460 24.150 1019.720 24.470 ;
        RECT 1019.520 2.400 1019.660 24.150 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 386.480 517.890 386.540 ;
        RECT 518.950 386.480 519.270 386.540 ;
        RECT 517.570 386.340 519.270 386.480 ;
        RECT 517.570 386.280 517.890 386.340 ;
        RECT 518.950 386.280 519.270 386.340 ;
        RECT 517.570 24.040 517.890 24.100 ;
        RECT 1036.910 24.040 1037.230 24.100 ;
        RECT 517.570 23.900 1037.230 24.040 ;
        RECT 517.570 23.840 517.890 23.900 ;
        RECT 1036.910 23.840 1037.230 23.900 ;
      LAYER via ;
        RECT 517.600 386.280 517.860 386.540 ;
        RECT 518.980 386.280 519.240 386.540 ;
        RECT 517.600 23.840 517.860 24.100 ;
        RECT 1036.940 23.840 1037.200 24.100 ;
      LAYER met2 ;
        RECT 519.330 400.250 519.610 404.000 ;
        RECT 519.040 400.110 519.610 400.250 ;
        RECT 519.040 386.570 519.180 400.110 ;
        RECT 519.330 400.000 519.610 400.110 ;
        RECT 517.600 386.250 517.860 386.570 ;
        RECT 518.980 386.250 519.240 386.570 ;
        RECT 517.660 24.130 517.800 386.250 ;
        RECT 517.600 23.810 517.860 24.130 ;
        RECT 1036.940 23.810 1037.200 24.130 ;
        RECT 1037.000 2.400 1037.140 23.810 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.850 400.250 525.130 404.000 ;
        RECT 524.560 400.110 525.130 400.250 ;
        RECT 524.560 25.685 524.700 400.110 ;
        RECT 524.850 400.000 525.130 400.110 ;
        RECT 524.490 25.315 524.770 25.685 ;
        RECT 1054.870 25.315 1055.150 25.685 ;
        RECT 1054.940 2.400 1055.080 25.315 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
      LAYER via2 ;
        RECT 524.490 25.360 524.770 25.640 ;
        RECT 1054.870 25.360 1055.150 25.640 ;
      LAYER met3 ;
        RECT 524.465 25.650 524.795 25.665 ;
        RECT 1054.845 25.650 1055.175 25.665 ;
        RECT 524.465 25.350 1055.175 25.650 ;
        RECT 524.465 25.335 524.795 25.350 ;
        RECT 1054.845 25.335 1055.175 25.350 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.370 400.250 530.650 404.000 ;
        RECT 529.160 400.110 530.650 400.250 ;
        RECT 529.160 386.650 529.300 400.110 ;
        RECT 530.370 400.000 530.650 400.110 ;
        RECT 525.480 386.510 529.300 386.650 ;
        RECT 525.480 25.005 525.620 386.510 ;
        RECT 525.410 24.635 525.690 25.005 ;
        RECT 1072.350 24.635 1072.630 25.005 ;
        RECT 1072.420 2.400 1072.560 24.635 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
      LAYER via2 ;
        RECT 525.410 24.680 525.690 24.960 ;
        RECT 1072.350 24.680 1072.630 24.960 ;
      LAYER met3 ;
        RECT 525.385 24.970 525.715 24.985 ;
        RECT 1072.325 24.970 1072.655 24.985 ;
        RECT 525.385 24.670 1072.655 24.970 ;
        RECT 525.385 24.655 525.715 24.670 ;
        RECT 1072.325 24.655 1072.655 24.670 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 547.930 390.560 548.250 390.620 ;
        RECT 755.390 390.560 755.710 390.620 ;
        RECT 547.930 390.420 755.710 390.560 ;
        RECT 547.930 390.360 548.250 390.420 ;
        RECT 755.390 390.360 755.710 390.420 ;
        RECT 535.510 388.520 535.830 388.580 ;
        RECT 547.930 388.520 548.250 388.580 ;
        RECT 535.510 388.380 548.250 388.520 ;
        RECT 535.510 388.320 535.830 388.380 ;
        RECT 547.930 388.320 548.250 388.380 ;
        RECT 755.390 28.800 755.710 28.860 ;
        RECT 1090.270 28.800 1090.590 28.860 ;
        RECT 755.390 28.660 1090.590 28.800 ;
        RECT 755.390 28.600 755.710 28.660 ;
        RECT 1090.270 28.600 1090.590 28.660 ;
      LAYER via ;
        RECT 547.960 390.360 548.220 390.620 ;
        RECT 755.420 390.360 755.680 390.620 ;
        RECT 535.540 388.320 535.800 388.580 ;
        RECT 547.960 388.320 548.220 388.580 ;
        RECT 755.420 28.600 755.680 28.860 ;
        RECT 1090.300 28.600 1090.560 28.860 ;
      LAYER met2 ;
        RECT 535.430 400.180 535.710 404.000 ;
        RECT 535.430 400.000 535.740 400.180 ;
        RECT 535.600 388.610 535.740 400.000 ;
        RECT 547.960 390.330 548.220 390.650 ;
        RECT 755.420 390.330 755.680 390.650 ;
        RECT 548.020 388.610 548.160 390.330 ;
        RECT 535.540 388.290 535.800 388.610 ;
        RECT 547.960 388.290 548.220 388.610 ;
        RECT 755.480 28.890 755.620 390.330 ;
        RECT 755.420 28.570 755.680 28.890 ;
        RECT 1090.300 28.570 1090.560 28.890 ;
        RECT 1090.360 2.400 1090.500 28.570 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.030 390.900 541.350 390.960 ;
        RECT 755.850 390.900 756.170 390.960 ;
        RECT 541.030 390.760 756.170 390.900 ;
        RECT 541.030 390.700 541.350 390.760 ;
        RECT 755.850 390.700 756.170 390.760 ;
        RECT 755.850 29.140 756.170 29.200 ;
        RECT 1107.750 29.140 1108.070 29.200 ;
        RECT 755.850 29.000 1108.070 29.140 ;
        RECT 755.850 28.940 756.170 29.000 ;
        RECT 1107.750 28.940 1108.070 29.000 ;
      LAYER via ;
        RECT 541.060 390.700 541.320 390.960 ;
        RECT 755.880 390.700 756.140 390.960 ;
        RECT 755.880 28.940 756.140 29.200 ;
        RECT 1107.780 28.940 1108.040 29.200 ;
      LAYER met2 ;
        RECT 540.950 400.180 541.230 404.000 ;
        RECT 540.950 400.000 541.260 400.180 ;
        RECT 541.120 390.990 541.260 400.000 ;
        RECT 541.060 390.670 541.320 390.990 ;
        RECT 755.880 390.670 756.140 390.990 ;
        RECT 755.940 29.230 756.080 390.670 ;
        RECT 755.880 28.910 756.140 29.230 ;
        RECT 1107.780 28.910 1108.040 29.230 ;
        RECT 1107.840 2.400 1107.980 28.910 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.550 388.860 546.870 388.920 ;
        RECT 638.550 388.860 638.870 388.920 ;
        RECT 546.550 388.720 638.870 388.860 ;
        RECT 546.550 388.660 546.870 388.720 ;
        RECT 638.550 388.660 638.870 388.720 ;
        RECT 638.090 29.480 638.410 29.540 ;
        RECT 1125.690 29.480 1126.010 29.540 ;
        RECT 638.090 29.340 1126.010 29.480 ;
        RECT 638.090 29.280 638.410 29.340 ;
        RECT 1125.690 29.280 1126.010 29.340 ;
      LAYER via ;
        RECT 546.580 388.660 546.840 388.920 ;
        RECT 638.580 388.660 638.840 388.920 ;
        RECT 638.120 29.280 638.380 29.540 ;
        RECT 1125.720 29.280 1125.980 29.540 ;
      LAYER met2 ;
        RECT 546.470 400.180 546.750 404.000 ;
        RECT 546.470 400.000 546.780 400.180 ;
        RECT 546.640 388.950 546.780 400.000 ;
        RECT 546.580 388.630 546.840 388.950 ;
        RECT 638.580 388.630 638.840 388.950 ;
        RECT 638.640 324.370 638.780 388.630 ;
        RECT 638.180 324.230 638.780 324.370 ;
        RECT 638.180 29.570 638.320 324.230 ;
        RECT 638.120 29.250 638.380 29.570 ;
        RECT 1125.720 29.250 1125.980 29.570 ;
        RECT 1125.780 2.400 1125.920 29.250 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.530 29.820 552.850 29.880 ;
        RECT 1143.630 29.820 1143.950 29.880 ;
        RECT 552.530 29.680 1143.950 29.820 ;
        RECT 552.530 29.620 552.850 29.680 ;
        RECT 1143.630 29.620 1143.950 29.680 ;
      LAYER via ;
        RECT 552.560 29.620 552.820 29.880 ;
        RECT 1143.660 29.620 1143.920 29.880 ;
      LAYER met2 ;
        RECT 551.990 400.250 552.270 404.000 ;
        RECT 551.990 400.110 552.760 400.250 ;
        RECT 551.990 400.000 552.270 400.110 ;
        RECT 552.620 29.910 552.760 400.110 ;
        RECT 552.560 29.590 552.820 29.910 ;
        RECT 1143.660 29.590 1143.920 29.910 ;
        RECT 1143.720 2.400 1143.860 29.590 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 375.940 400.590 376.000 ;
        RECT 403.030 375.940 403.350 376.000 ;
        RECT 400.270 375.800 403.350 375.940 ;
        RECT 400.270 375.740 400.590 375.800 ;
        RECT 403.030 375.740 403.350 375.800 ;
        RECT 400.270 23.020 400.590 23.080 ;
        RECT 664.770 23.020 665.090 23.080 ;
        RECT 400.270 22.880 665.090 23.020 ;
        RECT 400.270 22.820 400.590 22.880 ;
        RECT 664.770 22.820 665.090 22.880 ;
      LAYER via ;
        RECT 400.300 375.740 400.560 376.000 ;
        RECT 403.060 375.740 403.320 376.000 ;
        RECT 400.300 22.820 400.560 23.080 ;
        RECT 664.800 22.820 665.060 23.080 ;
      LAYER met2 ;
        RECT 404.330 400.250 404.610 404.000 ;
        RECT 403.120 400.110 404.610 400.250 ;
        RECT 403.120 376.030 403.260 400.110 ;
        RECT 404.330 400.000 404.610 400.110 ;
        RECT 400.300 375.710 400.560 376.030 ;
        RECT 403.060 375.710 403.320 376.030 ;
        RECT 400.360 23.110 400.500 375.710 ;
        RECT 400.300 22.790 400.560 23.110 ;
        RECT 664.800 22.790 665.060 23.110 ;
        RECT 664.860 2.400 665.000 22.790 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 376.280 552.390 376.340 ;
        RECT 556.210 376.280 556.530 376.340 ;
        RECT 552.070 376.140 556.530 376.280 ;
        RECT 552.070 376.080 552.390 376.140 ;
        RECT 556.210 376.080 556.530 376.140 ;
        RECT 552.070 30.160 552.390 30.220 ;
        RECT 1161.110 30.160 1161.430 30.220 ;
        RECT 552.070 30.020 1161.430 30.160 ;
        RECT 552.070 29.960 552.390 30.020 ;
        RECT 1161.110 29.960 1161.430 30.020 ;
      LAYER via ;
        RECT 552.100 376.080 552.360 376.340 ;
        RECT 556.240 376.080 556.500 376.340 ;
        RECT 552.100 29.960 552.360 30.220 ;
        RECT 1161.140 29.960 1161.400 30.220 ;
      LAYER met2 ;
        RECT 557.510 400.250 557.790 404.000 ;
        RECT 556.300 400.110 557.790 400.250 ;
        RECT 556.300 376.370 556.440 400.110 ;
        RECT 557.510 400.000 557.790 400.110 ;
        RECT 552.100 376.050 552.360 376.370 ;
        RECT 556.240 376.050 556.500 376.370 ;
        RECT 552.160 30.250 552.300 376.050 ;
        RECT 552.100 29.930 552.360 30.250 ;
        RECT 1161.140 29.930 1161.400 30.250 ;
        RECT 1161.200 2.400 1161.340 29.930 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 376.280 559.290 376.340 ;
        RECT 561.730 376.280 562.050 376.340 ;
        RECT 558.970 376.140 562.050 376.280 ;
        RECT 558.970 376.080 559.290 376.140 ;
        RECT 561.730 376.080 562.050 376.140 ;
        RECT 558.970 30.500 559.290 30.560 ;
        RECT 1179.050 30.500 1179.370 30.560 ;
        RECT 558.970 30.360 1179.370 30.500 ;
        RECT 558.970 30.300 559.290 30.360 ;
        RECT 1179.050 30.300 1179.370 30.360 ;
      LAYER via ;
        RECT 559.000 376.080 559.260 376.340 ;
        RECT 561.760 376.080 562.020 376.340 ;
        RECT 559.000 30.300 559.260 30.560 ;
        RECT 1179.080 30.300 1179.340 30.560 ;
      LAYER met2 ;
        RECT 563.030 400.250 563.310 404.000 ;
        RECT 561.820 400.110 563.310 400.250 ;
        RECT 561.820 376.370 561.960 400.110 ;
        RECT 563.030 400.000 563.310 400.110 ;
        RECT 559.000 376.050 559.260 376.370 ;
        RECT 561.760 376.050 562.020 376.370 ;
        RECT 559.060 30.590 559.200 376.050 ;
        RECT 559.000 30.270 559.260 30.590 ;
        RECT 1179.080 30.270 1179.340 30.590 ;
        RECT 1179.140 2.400 1179.280 30.270 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 376.280 566.190 376.340 ;
        RECT 567.250 376.280 567.570 376.340 ;
        RECT 565.870 376.140 567.570 376.280 ;
        RECT 565.870 376.080 566.190 376.140 ;
        RECT 567.250 376.080 567.570 376.140 ;
        RECT 565.870 34.240 566.190 34.300 ;
        RECT 1196.530 34.240 1196.850 34.300 ;
        RECT 565.870 34.100 1196.850 34.240 ;
        RECT 565.870 34.040 566.190 34.100 ;
        RECT 1196.530 34.040 1196.850 34.100 ;
      LAYER via ;
        RECT 565.900 376.080 566.160 376.340 ;
        RECT 567.280 376.080 567.540 376.340 ;
        RECT 565.900 34.040 566.160 34.300 ;
        RECT 1196.560 34.040 1196.820 34.300 ;
      LAYER met2 ;
        RECT 568.550 400.250 568.830 404.000 ;
        RECT 567.340 400.110 568.830 400.250 ;
        RECT 567.340 376.370 567.480 400.110 ;
        RECT 568.550 400.000 568.830 400.110 ;
        RECT 565.900 376.050 566.160 376.370 ;
        RECT 567.280 376.050 567.540 376.370 ;
        RECT 565.960 34.330 566.100 376.050 ;
        RECT 565.900 34.010 566.160 34.330 ;
        RECT 1196.560 34.010 1196.820 34.330 ;
        RECT 1196.620 2.400 1196.760 34.010 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 33.900 573.090 33.960 ;
        RECT 1214.930 33.900 1215.250 33.960 ;
        RECT 572.770 33.760 1215.250 33.900 ;
        RECT 572.770 33.700 573.090 33.760 ;
        RECT 1214.930 33.700 1215.250 33.760 ;
      LAYER via ;
        RECT 572.800 33.700 573.060 33.960 ;
        RECT 1214.960 33.700 1215.220 33.960 ;
      LAYER met2 ;
        RECT 574.070 400.250 574.350 404.000 ;
        RECT 572.860 400.110 574.350 400.250 ;
        RECT 572.860 33.990 573.000 400.110 ;
        RECT 574.070 400.000 574.350 400.110 ;
        RECT 572.800 33.670 573.060 33.990 ;
        RECT 1214.960 33.670 1215.220 33.990 ;
        RECT 1215.020 14.690 1215.160 33.670 ;
        RECT 1214.560 14.550 1215.160 14.690 ;
        RECT 1214.560 2.400 1214.700 14.550 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.130 33.560 580.450 33.620 ;
        RECT 1231.950 33.560 1232.270 33.620 ;
        RECT 580.130 33.420 1232.270 33.560 ;
        RECT 580.130 33.360 580.450 33.420 ;
        RECT 1231.950 33.360 1232.270 33.420 ;
      LAYER via ;
        RECT 580.160 33.360 580.420 33.620 ;
        RECT 1231.980 33.360 1232.240 33.620 ;
      LAYER met2 ;
        RECT 579.590 400.250 579.870 404.000 ;
        RECT 579.590 400.110 580.360 400.250 ;
        RECT 579.590 400.000 579.870 400.110 ;
        RECT 580.220 33.650 580.360 400.110 ;
        RECT 580.160 33.330 580.420 33.650 ;
        RECT 1231.980 33.330 1232.240 33.650 ;
        RECT 1232.040 2.400 1232.180 33.330 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.670 376.280 579.990 376.340 ;
        RECT 583.350 376.280 583.670 376.340 ;
        RECT 579.670 376.140 583.670 376.280 ;
        RECT 579.670 376.080 579.990 376.140 ;
        RECT 583.350 376.080 583.670 376.140 ;
        RECT 579.670 33.220 579.990 33.280 ;
        RECT 1249.890 33.220 1250.210 33.280 ;
        RECT 579.670 33.080 1250.210 33.220 ;
        RECT 579.670 33.020 579.990 33.080 ;
        RECT 1249.890 33.020 1250.210 33.080 ;
      LAYER via ;
        RECT 579.700 376.080 579.960 376.340 ;
        RECT 583.380 376.080 583.640 376.340 ;
        RECT 579.700 33.020 579.960 33.280 ;
        RECT 1249.920 33.020 1250.180 33.280 ;
      LAYER met2 ;
        RECT 584.650 400.250 584.930 404.000 ;
        RECT 583.440 400.110 584.930 400.250 ;
        RECT 583.440 376.370 583.580 400.110 ;
        RECT 584.650 400.000 584.930 400.110 ;
        RECT 579.700 376.050 579.960 376.370 ;
        RECT 583.380 376.050 583.640 376.370 ;
        RECT 579.760 33.310 579.900 376.050 ;
        RECT 579.700 32.990 579.960 33.310 ;
        RECT 1249.920 32.990 1250.180 33.310 ;
        RECT 1249.980 2.400 1250.120 32.990 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 375.940 586.890 376.000 ;
        RECT 588.870 375.940 589.190 376.000 ;
        RECT 586.570 375.800 589.190 375.940 ;
        RECT 586.570 375.740 586.890 375.800 ;
        RECT 588.870 375.740 589.190 375.800 ;
        RECT 586.570 32.880 586.890 32.940 ;
        RECT 1267.370 32.880 1267.690 32.940 ;
        RECT 586.570 32.740 1267.690 32.880 ;
        RECT 586.570 32.680 586.890 32.740 ;
        RECT 1267.370 32.680 1267.690 32.740 ;
      LAYER via ;
        RECT 586.600 375.740 586.860 376.000 ;
        RECT 588.900 375.740 589.160 376.000 ;
        RECT 586.600 32.680 586.860 32.940 ;
        RECT 1267.400 32.680 1267.660 32.940 ;
      LAYER met2 ;
        RECT 590.170 400.250 590.450 404.000 ;
        RECT 588.960 400.110 590.450 400.250 ;
        RECT 588.960 376.030 589.100 400.110 ;
        RECT 590.170 400.000 590.450 400.110 ;
        RECT 586.600 375.710 586.860 376.030 ;
        RECT 588.900 375.710 589.160 376.030 ;
        RECT 586.660 32.970 586.800 375.710 ;
        RECT 586.600 32.650 586.860 32.970 ;
        RECT 1267.400 32.650 1267.660 32.970 ;
        RECT 1267.460 2.400 1267.600 32.650 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 388.180 593.790 388.240 ;
        RECT 594.390 388.180 594.710 388.240 ;
        RECT 593.470 388.040 594.710 388.180 ;
        RECT 593.470 387.980 593.790 388.040 ;
        RECT 594.390 387.980 594.710 388.040 ;
        RECT 593.470 32.540 593.790 32.600 ;
        RECT 1285.310 32.540 1285.630 32.600 ;
        RECT 593.470 32.400 1285.630 32.540 ;
        RECT 593.470 32.340 593.790 32.400 ;
        RECT 1285.310 32.340 1285.630 32.400 ;
      LAYER via ;
        RECT 593.500 387.980 593.760 388.240 ;
        RECT 594.420 387.980 594.680 388.240 ;
        RECT 593.500 32.340 593.760 32.600 ;
        RECT 1285.340 32.340 1285.600 32.600 ;
      LAYER met2 ;
        RECT 595.690 400.250 595.970 404.000 ;
        RECT 594.480 400.110 595.970 400.250 ;
        RECT 594.480 388.270 594.620 400.110 ;
        RECT 595.690 400.000 595.970 400.110 ;
        RECT 593.500 387.950 593.760 388.270 ;
        RECT 594.420 387.950 594.680 388.270 ;
        RECT 593.560 32.630 593.700 387.950 ;
        RECT 593.500 32.310 593.760 32.630 ;
        RECT 1285.340 32.310 1285.600 32.630 ;
        RECT 1285.400 2.400 1285.540 32.310 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.830 32.200 601.150 32.260 ;
        RECT 1303.250 32.200 1303.570 32.260 ;
        RECT 600.830 32.060 1303.570 32.200 ;
        RECT 600.830 32.000 601.150 32.060 ;
        RECT 1303.250 32.000 1303.570 32.060 ;
      LAYER via ;
        RECT 600.860 32.000 601.120 32.260 ;
        RECT 1303.280 32.000 1303.540 32.260 ;
      LAYER met2 ;
        RECT 601.210 400.250 601.490 404.000 ;
        RECT 600.920 400.110 601.490 400.250 ;
        RECT 600.920 32.290 601.060 400.110 ;
        RECT 601.210 400.000 601.490 400.110 ;
        RECT 600.860 31.970 601.120 32.290 ;
        RECT 1303.280 31.970 1303.540 32.290 ;
        RECT 1303.340 2.400 1303.480 31.970 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 386.480 600.690 386.540 ;
        RECT 605.430 386.480 605.750 386.540 ;
        RECT 600.370 386.340 605.750 386.480 ;
        RECT 600.370 386.280 600.690 386.340 ;
        RECT 605.430 386.280 605.750 386.340 ;
      LAYER via ;
        RECT 600.400 386.280 600.660 386.540 ;
        RECT 605.460 386.280 605.720 386.540 ;
      LAYER met2 ;
        RECT 606.730 400.250 607.010 404.000 ;
        RECT 605.520 400.110 607.010 400.250 ;
        RECT 605.520 386.570 605.660 400.110 ;
        RECT 606.730 400.000 607.010 400.110 ;
        RECT 600.400 386.250 600.660 386.570 ;
        RECT 605.460 386.250 605.720 386.570 ;
        RECT 600.460 31.805 600.600 386.250 ;
        RECT 600.390 31.435 600.670 31.805 ;
        RECT 1320.750 31.435 1321.030 31.805 ;
        RECT 1320.820 2.400 1320.960 31.435 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
      LAYER via2 ;
        RECT 600.390 31.480 600.670 31.760 ;
        RECT 1320.750 31.480 1321.030 31.760 ;
      LAYER met3 ;
        RECT 600.365 31.770 600.695 31.785 ;
        RECT 1320.725 31.770 1321.055 31.785 ;
        RECT 600.365 31.470 1321.055 31.770 ;
        RECT 600.365 31.455 600.695 31.470 ;
        RECT 1320.725 31.455 1321.055 31.470 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 376.280 407.490 376.340 ;
        RECT 408.550 376.280 408.870 376.340 ;
        RECT 407.170 376.140 408.870 376.280 ;
        RECT 407.170 376.080 407.490 376.140 ;
        RECT 408.550 376.080 408.870 376.140 ;
        RECT 407.170 22.340 407.490 22.400 ;
        RECT 682.250 22.340 682.570 22.400 ;
        RECT 407.170 22.200 682.570 22.340 ;
        RECT 407.170 22.140 407.490 22.200 ;
        RECT 682.250 22.140 682.570 22.200 ;
      LAYER via ;
        RECT 407.200 376.080 407.460 376.340 ;
        RECT 408.580 376.080 408.840 376.340 ;
        RECT 407.200 22.140 407.460 22.400 ;
        RECT 682.280 22.140 682.540 22.400 ;
      LAYER met2 ;
        RECT 409.850 400.250 410.130 404.000 ;
        RECT 408.640 400.110 410.130 400.250 ;
        RECT 408.640 376.370 408.780 400.110 ;
        RECT 409.850 400.000 410.130 400.110 ;
        RECT 407.200 376.050 407.460 376.370 ;
        RECT 408.580 376.050 408.840 376.370 ;
        RECT 407.260 22.430 407.400 376.050 ;
        RECT 407.200 22.110 407.460 22.430 ;
        RECT 682.280 22.110 682.540 22.430 ;
        RECT 682.340 2.400 682.480 22.110 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.270 386.480 607.590 386.540 ;
        RECT 610.950 386.480 611.270 386.540 ;
        RECT 607.270 386.340 611.270 386.480 ;
        RECT 607.270 386.280 607.590 386.340 ;
        RECT 610.950 386.280 611.270 386.340 ;
      LAYER via ;
        RECT 607.300 386.280 607.560 386.540 ;
        RECT 610.980 386.280 611.240 386.540 ;
      LAYER met2 ;
        RECT 612.250 400.250 612.530 404.000 ;
        RECT 611.040 400.110 612.530 400.250 ;
        RECT 611.040 386.570 611.180 400.110 ;
        RECT 612.250 400.000 612.530 400.110 ;
        RECT 607.300 386.250 607.560 386.570 ;
        RECT 610.980 386.250 611.240 386.570 ;
        RECT 607.360 31.125 607.500 386.250 ;
        RECT 607.290 30.755 607.570 31.125 ;
        RECT 1338.690 30.755 1338.970 31.125 ;
        RECT 1338.760 2.400 1338.900 30.755 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
      LAYER via2 ;
        RECT 607.290 30.800 607.570 31.080 ;
        RECT 1338.690 30.800 1338.970 31.080 ;
      LAYER met3 ;
        RECT 607.265 31.090 607.595 31.105 ;
        RECT 1338.665 31.090 1338.995 31.105 ;
        RECT 607.265 30.790 1338.995 31.090 ;
        RECT 607.265 30.775 607.595 30.790 ;
        RECT 1338.665 30.775 1338.995 30.790 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.550 105.640 615.870 105.700 ;
        RECT 1352.470 105.640 1352.790 105.700 ;
        RECT 615.550 105.500 1352.790 105.640 ;
        RECT 615.550 105.440 615.870 105.500 ;
        RECT 1352.470 105.440 1352.790 105.500 ;
      LAYER via ;
        RECT 615.580 105.440 615.840 105.700 ;
        RECT 1352.500 105.440 1352.760 105.700 ;
      LAYER met2 ;
        RECT 617.770 400.250 618.050 404.000 ;
        RECT 616.560 400.110 618.050 400.250 ;
        RECT 616.560 324.370 616.700 400.110 ;
        RECT 617.770 400.000 618.050 400.110 ;
        RECT 615.640 324.230 616.700 324.370 ;
        RECT 615.640 105.730 615.780 324.230 ;
        RECT 615.580 105.410 615.840 105.730 ;
        RECT 1352.500 105.410 1352.760 105.730 ;
        RECT 1352.560 82.870 1352.700 105.410 ;
        RECT 1352.560 82.730 1354.080 82.870 ;
        RECT 1353.940 1.770 1354.080 82.730 ;
        RECT 1356.030 1.770 1356.590 2.400 ;
        RECT 1353.940 1.630 1356.590 1.770 ;
        RECT 1356.030 -4.800 1356.590 1.630 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 105.980 622.770 106.040 ;
        RECT 1373.170 105.980 1373.490 106.040 ;
        RECT 622.450 105.840 1373.490 105.980 ;
        RECT 622.450 105.780 622.770 105.840 ;
        RECT 1373.170 105.780 1373.490 105.840 ;
      LAYER via ;
        RECT 622.480 105.780 622.740 106.040 ;
        RECT 1373.200 105.780 1373.460 106.040 ;
      LAYER met2 ;
        RECT 623.290 400.250 623.570 404.000 ;
        RECT 622.540 400.110 623.570 400.250 ;
        RECT 622.540 106.070 622.680 400.110 ;
        RECT 623.290 400.000 623.570 400.110 ;
        RECT 622.480 105.750 622.740 106.070 ;
        RECT 1373.200 105.750 1373.460 106.070 ;
        RECT 1373.260 82.870 1373.400 105.750 ;
        RECT 1373.260 82.730 1374.320 82.870 ;
        RECT 1374.180 2.400 1374.320 82.730 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.890 106.320 629.210 106.380 ;
        RECT 1386.970 106.320 1387.290 106.380 ;
        RECT 628.890 106.180 1387.290 106.320 ;
        RECT 628.890 106.120 629.210 106.180 ;
        RECT 1386.970 106.120 1387.290 106.180 ;
      LAYER via ;
        RECT 628.920 106.120 629.180 106.380 ;
        RECT 1387.000 106.120 1387.260 106.380 ;
      LAYER met2 ;
        RECT 628.350 400.250 628.630 404.000 ;
        RECT 628.350 400.110 629.120 400.250 ;
        RECT 628.350 400.000 628.630 400.110 ;
        RECT 628.980 106.410 629.120 400.110 ;
        RECT 628.920 106.090 629.180 106.410 ;
        RECT 1387.000 106.090 1387.260 106.410 ;
        RECT 1387.060 82.870 1387.200 106.090 ;
        RECT 1387.060 82.730 1391.800 82.870 ;
        RECT 1391.660 2.400 1391.800 82.730 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.350 386.480 629.670 386.540 ;
        RECT 632.570 386.480 632.890 386.540 ;
        RECT 629.350 386.340 632.890 386.480 ;
        RECT 629.350 386.280 629.670 386.340 ;
        RECT 632.570 386.280 632.890 386.340 ;
        RECT 629.350 106.660 629.670 106.720 ;
        RECT 1407.670 106.660 1407.990 106.720 ;
        RECT 629.350 106.520 1407.990 106.660 ;
        RECT 629.350 106.460 629.670 106.520 ;
        RECT 1407.670 106.460 1407.990 106.520 ;
      LAYER via ;
        RECT 629.380 386.280 629.640 386.540 ;
        RECT 632.600 386.280 632.860 386.540 ;
        RECT 629.380 106.460 629.640 106.720 ;
        RECT 1407.700 106.460 1407.960 106.720 ;
      LAYER met2 ;
        RECT 633.870 400.250 634.150 404.000 ;
        RECT 632.660 400.110 634.150 400.250 ;
        RECT 632.660 386.570 632.800 400.110 ;
        RECT 633.870 400.000 634.150 400.110 ;
        RECT 629.380 386.250 629.640 386.570 ;
        RECT 632.600 386.250 632.860 386.570 ;
        RECT 629.440 106.750 629.580 386.250 ;
        RECT 629.380 106.430 629.640 106.750 ;
        RECT 1407.700 106.430 1407.960 106.750 ;
        RECT 1407.760 1.770 1407.900 106.430 ;
        RECT 1409.390 1.770 1409.950 2.400 ;
        RECT 1407.760 1.630 1409.950 1.770 ;
        RECT 1409.390 -4.800 1409.950 1.630 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.250 110.400 636.570 110.460 ;
        RECT 1421.470 110.400 1421.790 110.460 ;
        RECT 636.250 110.260 1421.790 110.400 ;
        RECT 636.250 110.200 636.570 110.260 ;
        RECT 1421.470 110.200 1421.790 110.260 ;
        RECT 1421.470 20.980 1421.790 21.040 ;
        RECT 1425.150 20.980 1425.470 21.040 ;
        RECT 1421.470 20.840 1425.470 20.980 ;
        RECT 1421.470 20.780 1421.790 20.840 ;
        RECT 1425.150 20.780 1425.470 20.840 ;
      LAYER via ;
        RECT 636.280 110.200 636.540 110.460 ;
        RECT 1421.500 110.200 1421.760 110.460 ;
        RECT 1421.500 20.780 1421.760 21.040 ;
        RECT 1425.180 20.780 1425.440 21.040 ;
      LAYER met2 ;
        RECT 639.390 400.250 639.670 404.000 ;
        RECT 638.180 400.110 639.670 400.250 ;
        RECT 638.180 386.140 638.320 400.110 ;
        RECT 639.390 400.000 639.670 400.110 ;
        RECT 636.340 386.000 638.320 386.140 ;
        RECT 636.340 110.490 636.480 386.000 ;
        RECT 636.280 110.170 636.540 110.490 ;
        RECT 1421.500 110.170 1421.760 110.490 ;
        RECT 1421.560 21.070 1421.700 110.170 ;
        RECT 1421.500 20.750 1421.760 21.070 ;
        RECT 1425.180 20.750 1425.440 21.070 ;
        RECT 1425.240 1.770 1425.380 20.750 ;
        RECT 1426.870 1.770 1427.430 2.400 ;
        RECT 1425.240 1.630 1427.430 1.770 ;
        RECT 1426.870 -4.800 1427.430 1.630 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 386.480 642.090 386.540 ;
        RECT 643.610 386.480 643.930 386.540 ;
        RECT 641.770 386.340 643.930 386.480 ;
        RECT 641.770 386.280 642.090 386.340 ;
        RECT 643.610 386.280 643.930 386.340 ;
        RECT 641.770 36.620 642.090 36.680 ;
        RECT 1444.930 36.620 1445.250 36.680 ;
        RECT 641.770 36.480 1445.250 36.620 ;
        RECT 641.770 36.420 642.090 36.480 ;
        RECT 1444.930 36.420 1445.250 36.480 ;
      LAYER via ;
        RECT 641.800 386.280 642.060 386.540 ;
        RECT 643.640 386.280 643.900 386.540 ;
        RECT 641.800 36.420 642.060 36.680 ;
        RECT 1444.960 36.420 1445.220 36.680 ;
      LAYER met2 ;
        RECT 644.910 400.250 645.190 404.000 ;
        RECT 643.700 400.110 645.190 400.250 ;
        RECT 643.700 386.570 643.840 400.110 ;
        RECT 644.910 400.000 645.190 400.110 ;
        RECT 641.800 386.250 642.060 386.570 ;
        RECT 643.640 386.250 643.900 386.570 ;
        RECT 641.860 36.710 642.000 386.250 ;
        RECT 641.800 36.390 642.060 36.710 ;
        RECT 1444.960 36.390 1445.220 36.710 ;
        RECT 1445.020 2.400 1445.160 36.390 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 36.960 648.990 37.020 ;
        RECT 1462.870 36.960 1463.190 37.020 ;
        RECT 648.670 36.820 1463.190 36.960 ;
        RECT 648.670 36.760 648.990 36.820 ;
        RECT 1462.870 36.760 1463.190 36.820 ;
      LAYER via ;
        RECT 648.700 36.760 648.960 37.020 ;
        RECT 1462.900 36.760 1463.160 37.020 ;
      LAYER met2 ;
        RECT 650.430 400.250 650.710 404.000 ;
        RECT 650.140 400.110 650.710 400.250 ;
        RECT 650.140 387.330 650.280 400.110 ;
        RECT 650.430 400.000 650.710 400.110 ;
        RECT 648.760 387.190 650.280 387.330 ;
        RECT 648.760 37.050 648.900 387.190 ;
        RECT 648.700 36.730 648.960 37.050 ;
        RECT 1462.900 36.730 1463.160 37.050 ;
        RECT 1462.960 2.400 1463.100 36.730 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.030 37.300 656.350 37.360 ;
        RECT 1480.350 37.300 1480.670 37.360 ;
        RECT 656.030 37.160 1480.670 37.300 ;
        RECT 656.030 37.100 656.350 37.160 ;
        RECT 1480.350 37.100 1480.670 37.160 ;
      LAYER via ;
        RECT 656.060 37.100 656.320 37.360 ;
        RECT 1480.380 37.100 1480.640 37.360 ;
      LAYER met2 ;
        RECT 655.950 400.180 656.230 404.000 ;
        RECT 655.950 400.000 656.260 400.180 ;
        RECT 656.120 37.390 656.260 400.000 ;
        RECT 656.060 37.070 656.320 37.390 ;
        RECT 1480.380 37.070 1480.640 37.390 ;
        RECT 1480.440 2.400 1480.580 37.070 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 655.570 386.480 655.890 386.540 ;
        RECT 660.170 386.480 660.490 386.540 ;
        RECT 655.570 386.340 660.490 386.480 ;
        RECT 655.570 386.280 655.890 386.340 ;
        RECT 660.170 386.280 660.490 386.340 ;
        RECT 655.570 37.640 655.890 37.700 ;
        RECT 1498.290 37.640 1498.610 37.700 ;
        RECT 655.570 37.500 1498.610 37.640 ;
        RECT 655.570 37.440 655.890 37.500 ;
        RECT 1498.290 37.440 1498.610 37.500 ;
      LAYER via ;
        RECT 655.600 386.280 655.860 386.540 ;
        RECT 660.200 386.280 660.460 386.540 ;
        RECT 655.600 37.440 655.860 37.700 ;
        RECT 1498.320 37.440 1498.580 37.700 ;
      LAYER met2 ;
        RECT 661.470 400.250 661.750 404.000 ;
        RECT 660.260 400.110 661.750 400.250 ;
        RECT 660.260 386.570 660.400 400.110 ;
        RECT 661.470 400.000 661.750 400.110 ;
        RECT 655.600 386.250 655.860 386.570 ;
        RECT 660.200 386.250 660.460 386.570 ;
        RECT 655.660 37.730 655.800 386.250 ;
        RECT 655.600 37.410 655.860 37.730 ;
        RECT 1498.320 37.410 1498.580 37.730 ;
        RECT 1498.380 2.400 1498.520 37.410 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 23.360 414.390 23.420 ;
        RECT 700.190 23.360 700.510 23.420 ;
        RECT 414.070 23.220 700.510 23.360 ;
        RECT 414.070 23.160 414.390 23.220 ;
        RECT 700.190 23.160 700.510 23.220 ;
      LAYER via ;
        RECT 414.100 23.160 414.360 23.420 ;
        RECT 700.220 23.160 700.480 23.420 ;
      LAYER met2 ;
        RECT 415.370 400.250 415.650 404.000 ;
        RECT 414.160 400.110 415.650 400.250 ;
        RECT 414.160 23.450 414.300 400.110 ;
        RECT 415.370 400.000 415.650 400.110 ;
        RECT 414.100 23.130 414.360 23.450 ;
        RECT 700.220 23.130 700.480 23.450 ;
        RECT 700.280 2.400 700.420 23.130 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 386.820 662.790 386.880 ;
        RECT 665.690 386.820 666.010 386.880 ;
        RECT 662.470 386.680 666.010 386.820 ;
        RECT 662.470 386.620 662.790 386.680 ;
        RECT 665.690 386.620 666.010 386.680 ;
        RECT 662.470 41.380 662.790 41.440 ;
        RECT 1515.770 41.380 1516.090 41.440 ;
        RECT 662.470 41.240 1516.090 41.380 ;
        RECT 662.470 41.180 662.790 41.240 ;
        RECT 1515.770 41.180 1516.090 41.240 ;
      LAYER via ;
        RECT 662.500 386.620 662.760 386.880 ;
        RECT 665.720 386.620 665.980 386.880 ;
        RECT 662.500 41.180 662.760 41.440 ;
        RECT 1515.800 41.180 1516.060 41.440 ;
      LAYER met2 ;
        RECT 666.990 400.250 667.270 404.000 ;
        RECT 665.780 400.110 667.270 400.250 ;
        RECT 665.780 386.910 665.920 400.110 ;
        RECT 666.990 400.000 667.270 400.110 ;
        RECT 662.500 386.590 662.760 386.910 ;
        RECT 665.720 386.590 665.980 386.910 ;
        RECT 662.560 41.470 662.700 386.590 ;
        RECT 662.500 41.150 662.760 41.470 ;
        RECT 1515.800 41.150 1516.060 41.470 ;
        RECT 1515.860 2.400 1516.000 41.150 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.370 41.040 669.690 41.100 ;
        RECT 1533.710 41.040 1534.030 41.100 ;
        RECT 669.370 40.900 1534.030 41.040 ;
        RECT 669.370 40.840 669.690 40.900 ;
        RECT 1533.710 40.840 1534.030 40.900 ;
      LAYER via ;
        RECT 669.400 40.840 669.660 41.100 ;
        RECT 1533.740 40.840 1534.000 41.100 ;
      LAYER met2 ;
        RECT 672.510 400.250 672.790 404.000 ;
        RECT 671.300 400.110 672.790 400.250 ;
        RECT 671.300 388.010 671.440 400.110 ;
        RECT 672.510 400.000 672.790 400.110 ;
        RECT 669.460 387.870 671.440 388.010 ;
        RECT 669.460 41.130 669.600 387.870 ;
        RECT 669.400 40.810 669.660 41.130 ;
        RECT 1533.740 40.810 1534.000 41.130 ;
        RECT 1533.800 2.400 1533.940 40.810 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.270 40.700 676.590 40.760 ;
        RECT 1551.190 40.700 1551.510 40.760 ;
        RECT 676.270 40.560 1551.510 40.700 ;
        RECT 676.270 40.500 676.590 40.560 ;
        RECT 1551.190 40.500 1551.510 40.560 ;
      LAYER via ;
        RECT 676.300 40.500 676.560 40.760 ;
        RECT 1551.220 40.500 1551.480 40.760 ;
      LAYER met2 ;
        RECT 677.570 400.250 677.850 404.000 ;
        RECT 676.360 400.110 677.850 400.250 ;
        RECT 676.360 40.790 676.500 400.110 ;
        RECT 677.570 400.000 677.850 400.110 ;
        RECT 676.300 40.470 676.560 40.790 ;
        RECT 1551.220 40.470 1551.480 40.790 ;
        RECT 1551.280 2.400 1551.420 40.470 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.170 40.360 683.490 40.420 ;
        RECT 1569.130 40.360 1569.450 40.420 ;
        RECT 683.170 40.220 1569.450 40.360 ;
        RECT 683.170 40.160 683.490 40.220 ;
        RECT 1569.130 40.160 1569.450 40.220 ;
      LAYER via ;
        RECT 683.200 40.160 683.460 40.420 ;
        RECT 1569.160 40.160 1569.420 40.420 ;
      LAYER met2 ;
        RECT 683.090 400.180 683.370 404.000 ;
        RECT 683.090 400.000 683.400 400.180 ;
        RECT 683.260 40.450 683.400 400.000 ;
        RECT 683.200 40.130 683.460 40.450 ;
        RECT 1569.160 40.130 1569.420 40.450 ;
        RECT 1569.220 2.400 1569.360 40.130 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 386.480 683.950 386.540 ;
        RECT 687.310 386.480 687.630 386.540 ;
        RECT 683.630 386.340 687.630 386.480 ;
        RECT 683.630 386.280 683.950 386.340 ;
        RECT 687.310 386.280 687.630 386.340 ;
        RECT 683.630 40.020 683.950 40.080 ;
        RECT 1586.610 40.020 1586.930 40.080 ;
        RECT 683.630 39.880 1586.930 40.020 ;
        RECT 683.630 39.820 683.950 39.880 ;
        RECT 1586.610 39.820 1586.930 39.880 ;
      LAYER via ;
        RECT 683.660 386.280 683.920 386.540 ;
        RECT 687.340 386.280 687.600 386.540 ;
        RECT 683.660 39.820 683.920 40.080 ;
        RECT 1586.640 39.820 1586.900 40.080 ;
      LAYER met2 ;
        RECT 688.610 400.250 688.890 404.000 ;
        RECT 687.400 400.110 688.890 400.250 ;
        RECT 687.400 386.570 687.540 400.110 ;
        RECT 688.610 400.000 688.890 400.110 ;
        RECT 683.660 386.250 683.920 386.570 ;
        RECT 687.340 386.250 687.600 386.570 ;
        RECT 683.720 40.110 683.860 386.250 ;
        RECT 683.660 39.790 683.920 40.110 ;
        RECT 1586.640 39.790 1586.900 40.110 ;
        RECT 1586.700 2.400 1586.840 39.790 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.070 384.100 690.390 384.160 ;
        RECT 692.830 384.100 693.150 384.160 ;
        RECT 690.070 383.960 693.150 384.100 ;
        RECT 690.070 383.900 690.390 383.960 ;
        RECT 692.830 383.900 693.150 383.960 ;
        RECT 690.070 39.680 690.390 39.740 ;
        RECT 1604.550 39.680 1604.870 39.740 ;
        RECT 690.070 39.540 1604.870 39.680 ;
        RECT 690.070 39.480 690.390 39.540 ;
        RECT 1604.550 39.480 1604.870 39.540 ;
      LAYER via ;
        RECT 690.100 383.900 690.360 384.160 ;
        RECT 692.860 383.900 693.120 384.160 ;
        RECT 690.100 39.480 690.360 39.740 ;
        RECT 1604.580 39.480 1604.840 39.740 ;
      LAYER met2 ;
        RECT 694.130 400.250 694.410 404.000 ;
        RECT 692.920 400.110 694.410 400.250 ;
        RECT 692.920 384.190 693.060 400.110 ;
        RECT 694.130 400.000 694.410 400.110 ;
        RECT 690.100 383.870 690.360 384.190 ;
        RECT 692.860 383.870 693.120 384.190 ;
        RECT 690.160 39.770 690.300 383.870 ;
        RECT 690.100 39.450 690.360 39.770 ;
        RECT 1604.580 39.450 1604.840 39.770 ;
        RECT 1604.640 2.400 1604.780 39.450 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.970 376.280 697.290 376.340 ;
        RECT 699.730 376.280 700.050 376.340 ;
        RECT 696.970 376.140 700.050 376.280 ;
        RECT 696.970 376.080 697.290 376.140 ;
        RECT 699.730 376.080 700.050 376.140 ;
        RECT 696.970 39.340 697.290 39.400 ;
        RECT 1622.030 39.340 1622.350 39.400 ;
        RECT 696.970 39.200 1622.350 39.340 ;
        RECT 696.970 39.140 697.290 39.200 ;
        RECT 1622.030 39.140 1622.350 39.200 ;
      LAYER via ;
        RECT 697.000 376.080 697.260 376.340 ;
        RECT 699.760 376.080 700.020 376.340 ;
        RECT 697.000 39.140 697.260 39.400 ;
        RECT 1622.060 39.140 1622.320 39.400 ;
      LAYER met2 ;
        RECT 699.650 400.180 699.930 404.000 ;
        RECT 699.650 400.000 699.960 400.180 ;
        RECT 699.820 376.370 699.960 400.000 ;
        RECT 697.000 376.050 697.260 376.370 ;
        RECT 699.760 376.050 700.020 376.370 ;
        RECT 697.060 39.430 697.200 376.050 ;
        RECT 697.000 39.110 697.260 39.430 ;
        RECT 1622.060 39.110 1622.320 39.430 ;
        RECT 1622.120 2.400 1622.260 39.110 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.870 39.000 704.190 39.060 ;
        RECT 1639.970 39.000 1640.290 39.060 ;
        RECT 703.870 38.860 1640.290 39.000 ;
        RECT 703.870 38.800 704.190 38.860 ;
        RECT 1639.970 38.800 1640.290 38.860 ;
      LAYER via ;
        RECT 703.900 38.800 704.160 39.060 ;
        RECT 1640.000 38.800 1640.260 39.060 ;
      LAYER met2 ;
        RECT 705.170 400.250 705.450 404.000 ;
        RECT 703.960 400.110 705.450 400.250 ;
        RECT 703.960 39.090 704.100 400.110 ;
        RECT 705.170 400.000 705.450 400.110 ;
        RECT 703.900 38.770 704.160 39.090 ;
        RECT 1640.000 38.770 1640.260 39.090 ;
        RECT 1640.060 2.400 1640.200 38.770 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 710.770 38.660 711.090 38.720 ;
        RECT 1657.910 38.660 1658.230 38.720 ;
        RECT 710.770 38.520 1658.230 38.660 ;
        RECT 710.770 38.460 711.090 38.520 ;
        RECT 1657.910 38.460 1658.230 38.520 ;
      LAYER via ;
        RECT 710.800 38.460 711.060 38.720 ;
        RECT 1657.940 38.460 1658.200 38.720 ;
      LAYER met2 ;
        RECT 710.690 400.180 710.970 404.000 ;
        RECT 710.690 400.000 711.000 400.180 ;
        RECT 710.860 38.750 711.000 400.000 ;
        RECT 710.800 38.430 711.060 38.750 ;
        RECT 1657.940 38.430 1658.200 38.750 ;
        RECT 1658.000 2.400 1658.140 38.430 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.230 376.280 711.550 376.340 ;
        RECT 714.910 376.280 715.230 376.340 ;
        RECT 711.230 376.140 715.230 376.280 ;
        RECT 711.230 376.080 711.550 376.140 ;
        RECT 714.910 376.080 715.230 376.140 ;
        RECT 711.230 38.320 711.550 38.380 ;
        RECT 1675.390 38.320 1675.710 38.380 ;
        RECT 711.230 38.180 1675.710 38.320 ;
        RECT 711.230 38.120 711.550 38.180 ;
        RECT 1675.390 38.120 1675.710 38.180 ;
      LAYER via ;
        RECT 711.260 376.080 711.520 376.340 ;
        RECT 714.940 376.080 715.200 376.340 ;
        RECT 711.260 38.120 711.520 38.380 ;
        RECT 1675.420 38.120 1675.680 38.380 ;
      LAYER met2 ;
        RECT 716.210 400.250 716.490 404.000 ;
        RECT 715.000 400.110 716.490 400.250 ;
        RECT 715.000 376.370 715.140 400.110 ;
        RECT 716.210 400.000 716.490 400.110 ;
        RECT 711.260 376.050 711.520 376.370 ;
        RECT 714.940 376.050 715.200 376.370 ;
        RECT 711.320 38.410 711.460 376.050 ;
        RECT 711.260 38.090 711.520 38.410 ;
        RECT 1675.420 38.090 1675.680 38.410 ;
        RECT 1675.480 2.400 1675.620 38.090 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 27.440 421.290 27.500 ;
        RECT 717.670 27.440 717.990 27.500 ;
        RECT 420.970 27.300 717.990 27.440 ;
        RECT 420.970 27.240 421.290 27.300 ;
        RECT 717.670 27.240 717.990 27.300 ;
      LAYER via ;
        RECT 421.000 27.240 421.260 27.500 ;
        RECT 717.700 27.240 717.960 27.500 ;
      LAYER met2 ;
        RECT 420.890 400.180 421.170 404.000 ;
        RECT 420.890 400.000 421.200 400.180 ;
        RECT 421.060 27.530 421.200 400.000 ;
        RECT 421.000 27.210 421.260 27.530 ;
        RECT 717.700 27.210 717.960 27.530 ;
        RECT 717.760 2.400 717.900 27.210 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 717.670 375.940 717.990 376.000 ;
        RECT 720.430 375.940 720.750 376.000 ;
        RECT 717.670 375.800 720.750 375.940 ;
        RECT 717.670 375.740 717.990 375.800 ;
        RECT 720.430 375.740 720.750 375.800 ;
        RECT 717.670 37.980 717.990 38.040 ;
        RECT 1693.330 37.980 1693.650 38.040 ;
        RECT 717.670 37.840 1693.650 37.980 ;
        RECT 717.670 37.780 717.990 37.840 ;
        RECT 1693.330 37.780 1693.650 37.840 ;
      LAYER via ;
        RECT 717.700 375.740 717.960 376.000 ;
        RECT 720.460 375.740 720.720 376.000 ;
        RECT 717.700 37.780 717.960 38.040 ;
        RECT 1693.360 37.780 1693.620 38.040 ;
      LAYER met2 ;
        RECT 721.730 400.250 722.010 404.000 ;
        RECT 720.520 400.110 722.010 400.250 ;
        RECT 720.520 376.030 720.660 400.110 ;
        RECT 721.730 400.000 722.010 400.110 ;
        RECT 717.700 375.710 717.960 376.030 ;
        RECT 720.460 375.710 720.720 376.030 ;
        RECT 717.760 38.070 717.900 375.710 ;
        RECT 717.700 37.750 717.960 38.070 ;
        RECT 1693.360 37.750 1693.620 38.070 ;
        RECT 1693.420 2.400 1693.560 37.750 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.570 379.000 724.890 379.060 ;
        RECT 726.870 379.000 727.190 379.060 ;
        RECT 724.570 378.860 727.190 379.000 ;
        RECT 724.570 378.800 724.890 378.860 ;
        RECT 726.870 378.800 727.190 378.860 ;
      LAYER via ;
        RECT 724.600 378.800 724.860 379.060 ;
        RECT 726.900 378.800 727.160 379.060 ;
      LAYER met2 ;
        RECT 726.790 400.180 727.070 404.000 ;
        RECT 726.790 400.000 727.100 400.180 ;
        RECT 726.960 379.090 727.100 400.000 ;
        RECT 724.600 378.770 724.860 379.090 ;
        RECT 726.900 378.770 727.160 379.090 ;
        RECT 724.660 38.605 724.800 378.770 ;
        RECT 724.590 38.235 724.870 38.605 ;
        RECT 1710.830 38.235 1711.110 38.605 ;
        RECT 1710.900 2.400 1711.040 38.235 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
      LAYER via2 ;
        RECT 724.590 38.280 724.870 38.560 ;
        RECT 1710.830 38.280 1711.110 38.560 ;
      LAYER met3 ;
        RECT 724.565 38.570 724.895 38.585 ;
        RECT 1710.805 38.570 1711.135 38.585 ;
        RECT 724.565 38.270 1711.135 38.570 ;
        RECT 724.565 38.255 724.895 38.270 ;
        RECT 1710.805 38.255 1711.135 38.270 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.310 400.250 732.590 404.000 ;
        RECT 731.560 400.110 732.590 400.250 ;
        RECT 731.560 37.925 731.700 400.110 ;
        RECT 732.310 400.000 732.590 400.110 ;
        RECT 731.490 37.555 731.770 37.925 ;
        RECT 1728.770 37.555 1729.050 37.925 ;
        RECT 1728.840 2.400 1728.980 37.555 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
      LAYER via2 ;
        RECT 731.490 37.600 731.770 37.880 ;
        RECT 1728.770 37.600 1729.050 37.880 ;
      LAYER met3 ;
        RECT 731.465 37.890 731.795 37.905 ;
        RECT 1728.745 37.890 1729.075 37.905 ;
        RECT 731.465 37.590 1729.075 37.890 ;
        RECT 731.465 37.575 731.795 37.590 ;
        RECT 1728.745 37.575 1729.075 37.590 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.390 376.280 732.710 376.340 ;
        RECT 736.530 376.280 736.850 376.340 ;
        RECT 732.390 376.140 736.850 376.280 ;
        RECT 732.390 376.080 732.710 376.140 ;
        RECT 736.530 376.080 736.850 376.140 ;
        RECT 732.390 110.060 732.710 110.120 ;
        RECT 1745.770 110.060 1746.090 110.120 ;
        RECT 732.390 109.920 1746.090 110.060 ;
        RECT 732.390 109.860 732.710 109.920 ;
        RECT 1745.770 109.860 1746.090 109.920 ;
      LAYER via ;
        RECT 732.420 376.080 732.680 376.340 ;
        RECT 736.560 376.080 736.820 376.340 ;
        RECT 732.420 109.860 732.680 110.120 ;
        RECT 1745.800 109.860 1746.060 110.120 ;
      LAYER met2 ;
        RECT 737.830 400.250 738.110 404.000 ;
        RECT 736.620 400.110 738.110 400.250 ;
        RECT 736.620 376.370 736.760 400.110 ;
        RECT 737.830 400.000 738.110 400.110 ;
        RECT 732.420 376.050 732.680 376.370 ;
        RECT 736.560 376.050 736.820 376.370 ;
        RECT 732.480 110.150 732.620 376.050 ;
        RECT 732.420 109.830 732.680 110.150 ;
        RECT 1745.800 109.830 1746.060 110.150 ;
        RECT 1745.860 14.690 1746.000 109.830 ;
        RECT 1745.860 14.550 1746.460 14.690 ;
        RECT 1746.320 2.400 1746.460 14.550 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.830 376.280 739.150 376.340 ;
        RECT 742.050 376.280 742.370 376.340 ;
        RECT 738.830 376.140 742.370 376.280 ;
        RECT 738.830 376.080 739.150 376.140 ;
        RECT 742.050 376.080 742.370 376.140 ;
        RECT 738.830 109.720 739.150 109.780 ;
        RECT 1759.570 109.720 1759.890 109.780 ;
        RECT 738.830 109.580 1759.890 109.720 ;
        RECT 738.830 109.520 739.150 109.580 ;
        RECT 1759.570 109.520 1759.890 109.580 ;
      LAYER via ;
        RECT 738.860 376.080 739.120 376.340 ;
        RECT 742.080 376.080 742.340 376.340 ;
        RECT 738.860 109.520 739.120 109.780 ;
        RECT 1759.600 109.520 1759.860 109.780 ;
      LAYER met2 ;
        RECT 743.350 400.250 743.630 404.000 ;
        RECT 742.140 400.110 743.630 400.250 ;
        RECT 742.140 376.370 742.280 400.110 ;
        RECT 743.350 400.000 743.630 400.110 ;
        RECT 738.860 376.050 739.120 376.370 ;
        RECT 742.080 376.050 742.340 376.370 ;
        RECT 738.920 109.810 739.060 376.050 ;
        RECT 738.860 109.490 739.120 109.810 ;
        RECT 1759.600 109.490 1759.860 109.810 ;
        RECT 1759.660 82.870 1759.800 109.490 ;
        RECT 1759.660 82.730 1764.400 82.870 ;
        RECT 1764.260 2.400 1764.400 82.730 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 746.190 375.940 746.510 376.000 ;
        RECT 747.570 375.940 747.890 376.000 ;
        RECT 746.190 375.800 747.890 375.940 ;
        RECT 746.190 375.740 746.510 375.800 ;
        RECT 747.570 375.740 747.890 375.800 ;
        RECT 746.190 109.380 746.510 109.440 ;
        RECT 1780.270 109.380 1780.590 109.440 ;
        RECT 746.190 109.240 1780.590 109.380 ;
        RECT 746.190 109.180 746.510 109.240 ;
        RECT 1780.270 109.180 1780.590 109.240 ;
      LAYER via ;
        RECT 746.220 375.740 746.480 376.000 ;
        RECT 747.600 375.740 747.860 376.000 ;
        RECT 746.220 109.180 746.480 109.440 ;
        RECT 1780.300 109.180 1780.560 109.440 ;
      LAYER met2 ;
        RECT 748.870 400.250 749.150 404.000 ;
        RECT 747.660 400.110 749.150 400.250 ;
        RECT 747.660 376.030 747.800 400.110 ;
        RECT 748.870 400.000 749.150 400.110 ;
        RECT 746.220 375.710 746.480 376.030 ;
        RECT 747.600 375.710 747.860 376.030 ;
        RECT 746.280 109.470 746.420 375.710 ;
        RECT 746.220 109.150 746.480 109.470 ;
        RECT 1780.300 109.150 1780.560 109.470 ;
        RECT 1780.360 82.870 1780.500 109.150 ;
        RECT 1780.360 82.730 1781.880 82.870 ;
        RECT 1781.740 2.400 1781.880 82.730 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.630 386.820 752.950 386.880 ;
        RECT 754.470 386.820 754.790 386.880 ;
        RECT 752.630 386.680 754.790 386.820 ;
        RECT 752.630 386.620 752.950 386.680 ;
        RECT 754.470 386.620 754.790 386.680 ;
        RECT 752.630 109.040 752.950 109.100 ;
        RECT 1794.070 109.040 1794.390 109.100 ;
        RECT 752.630 108.900 1794.390 109.040 ;
        RECT 752.630 108.840 752.950 108.900 ;
        RECT 1794.070 108.840 1794.390 108.900 ;
      LAYER via ;
        RECT 752.660 386.620 752.920 386.880 ;
        RECT 754.500 386.620 754.760 386.880 ;
        RECT 752.660 108.840 752.920 109.100 ;
        RECT 1794.100 108.840 1794.360 109.100 ;
      LAYER met2 ;
        RECT 754.390 400.180 754.670 404.000 ;
        RECT 754.390 400.000 754.700 400.180 ;
        RECT 754.560 386.910 754.700 400.000 ;
        RECT 752.660 386.590 752.920 386.910 ;
        RECT 754.500 386.590 754.760 386.910 ;
        RECT 752.720 109.130 752.860 386.590 ;
        RECT 752.660 108.810 752.920 109.130 ;
        RECT 1794.100 108.810 1794.360 109.130 ;
        RECT 1794.160 82.870 1794.300 108.810 ;
        RECT 1794.160 82.730 1797.520 82.870 ;
        RECT 1797.380 1.770 1797.520 82.730 ;
        RECT 1799.470 1.770 1800.030 2.400 ;
        RECT 1797.380 1.630 1800.030 1.770 ;
        RECT 1799.470 -4.800 1800.030 1.630 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.990 116.520 760.310 116.580 ;
        RECT 1814.770 116.520 1815.090 116.580 ;
        RECT 759.990 116.380 1815.090 116.520 ;
        RECT 759.990 116.320 760.310 116.380 ;
        RECT 1814.770 116.320 1815.090 116.380 ;
      LAYER via ;
        RECT 760.020 116.320 760.280 116.580 ;
        RECT 1814.800 116.320 1815.060 116.580 ;
      LAYER met2 ;
        RECT 759.910 400.180 760.190 404.000 ;
        RECT 759.910 400.000 760.220 400.180 ;
        RECT 760.080 116.610 760.220 400.000 ;
        RECT 760.020 116.290 760.280 116.610 ;
        RECT 1814.800 116.290 1815.060 116.610 ;
        RECT 1814.860 82.870 1815.000 116.290 ;
        RECT 1814.860 82.730 1817.760 82.870 ;
        RECT 1817.620 2.400 1817.760 82.730 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.070 375.940 759.390 376.000 ;
        RECT 764.130 375.940 764.450 376.000 ;
        RECT 759.070 375.800 764.450 375.940 ;
        RECT 759.070 375.740 759.390 375.800 ;
        RECT 764.130 375.740 764.450 375.800 ;
        RECT 759.530 43.420 759.850 43.480 ;
        RECT 1835.010 43.420 1835.330 43.480 ;
        RECT 759.530 43.280 1835.330 43.420 ;
        RECT 759.530 43.220 759.850 43.280 ;
        RECT 1835.010 43.220 1835.330 43.280 ;
      LAYER via ;
        RECT 759.100 375.740 759.360 376.000 ;
        RECT 764.160 375.740 764.420 376.000 ;
        RECT 759.560 43.220 759.820 43.480 ;
        RECT 1835.040 43.220 1835.300 43.480 ;
      LAYER met2 ;
        RECT 765.430 400.250 765.710 404.000 ;
        RECT 764.220 400.110 765.710 400.250 ;
        RECT 764.220 376.030 764.360 400.110 ;
        RECT 765.430 400.000 765.710 400.110 ;
        RECT 759.100 375.710 759.360 376.030 ;
        RECT 764.160 375.710 764.420 376.030 ;
        RECT 759.160 62.970 759.300 375.710 ;
        RECT 759.160 62.830 759.760 62.970 ;
        RECT 759.620 43.510 759.760 62.830 ;
        RECT 759.560 43.190 759.820 43.510 ;
        RECT 1835.040 43.190 1835.300 43.510 ;
        RECT 1835.100 2.400 1835.240 43.190 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.970 376.280 766.290 376.340 ;
        RECT 769.650 376.280 769.970 376.340 ;
        RECT 765.970 376.140 769.970 376.280 ;
        RECT 765.970 376.080 766.290 376.140 ;
        RECT 769.650 376.080 769.970 376.140 ;
        RECT 765.970 43.760 766.290 43.820 ;
        RECT 1852.950 43.760 1853.270 43.820 ;
        RECT 765.970 43.620 1853.270 43.760 ;
        RECT 765.970 43.560 766.290 43.620 ;
        RECT 1852.950 43.560 1853.270 43.620 ;
      LAYER via ;
        RECT 766.000 376.080 766.260 376.340 ;
        RECT 769.680 376.080 769.940 376.340 ;
        RECT 766.000 43.560 766.260 43.820 ;
        RECT 1852.980 43.560 1853.240 43.820 ;
      LAYER met2 ;
        RECT 770.490 400.250 770.770 404.000 ;
        RECT 769.740 400.110 770.770 400.250 ;
        RECT 769.740 376.370 769.880 400.110 ;
        RECT 770.490 400.000 770.770 400.110 ;
        RECT 766.000 376.050 766.260 376.370 ;
        RECT 769.680 376.050 769.940 376.370 ;
        RECT 766.060 43.850 766.200 376.050 ;
        RECT 766.000 43.530 766.260 43.850 ;
        RECT 1852.980 43.530 1853.240 43.850 ;
        RECT 1853.040 2.400 1853.180 43.530 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.430 376.280 421.750 376.340 ;
        RECT 425.110 376.280 425.430 376.340 ;
        RECT 421.430 376.140 425.430 376.280 ;
        RECT 421.430 376.080 421.750 376.140 ;
        RECT 425.110 376.080 425.430 376.140 ;
        RECT 421.430 27.100 421.750 27.160 ;
        RECT 735.610 27.100 735.930 27.160 ;
        RECT 421.430 26.960 735.930 27.100 ;
        RECT 421.430 26.900 421.750 26.960 ;
        RECT 735.610 26.900 735.930 26.960 ;
      LAYER via ;
        RECT 421.460 376.080 421.720 376.340 ;
        RECT 425.140 376.080 425.400 376.340 ;
        RECT 421.460 26.900 421.720 27.160 ;
        RECT 735.640 26.900 735.900 27.160 ;
      LAYER met2 ;
        RECT 426.410 400.250 426.690 404.000 ;
        RECT 425.200 400.110 426.690 400.250 ;
        RECT 425.200 376.370 425.340 400.110 ;
        RECT 426.410 400.000 426.690 400.110 ;
        RECT 421.460 376.050 421.720 376.370 ;
        RECT 425.140 376.050 425.400 376.370 ;
        RECT 421.520 27.190 421.660 376.050 ;
        RECT 421.460 26.870 421.720 27.190 ;
        RECT 735.640 26.870 735.900 27.190 ;
        RECT 735.700 2.400 735.840 26.870 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 772.870 376.280 773.190 376.340 ;
        RECT 774.710 376.280 775.030 376.340 ;
        RECT 772.870 376.140 775.030 376.280 ;
        RECT 772.870 376.080 773.190 376.140 ;
        RECT 774.710 376.080 775.030 376.140 ;
        RECT 772.870 44.100 773.190 44.160 ;
        RECT 1870.430 44.100 1870.750 44.160 ;
        RECT 772.870 43.960 1870.750 44.100 ;
        RECT 772.870 43.900 773.190 43.960 ;
        RECT 1870.430 43.900 1870.750 43.960 ;
      LAYER via ;
        RECT 772.900 376.080 773.160 376.340 ;
        RECT 774.740 376.080 775.000 376.340 ;
        RECT 772.900 43.900 773.160 44.160 ;
        RECT 1870.460 43.900 1870.720 44.160 ;
      LAYER met2 ;
        RECT 776.010 400.250 776.290 404.000 ;
        RECT 774.800 400.110 776.290 400.250 ;
        RECT 774.800 376.370 774.940 400.110 ;
        RECT 776.010 400.000 776.290 400.110 ;
        RECT 772.900 376.050 773.160 376.370 ;
        RECT 774.740 376.050 775.000 376.370 ;
        RECT 772.960 44.190 773.100 376.050 ;
        RECT 772.900 43.870 773.160 44.190 ;
        RECT 1870.460 43.870 1870.720 44.190 ;
        RECT 1870.520 2.400 1870.660 43.870 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 779.770 44.440 780.090 44.500 ;
        RECT 1888.370 44.440 1888.690 44.500 ;
        RECT 779.770 44.300 1888.690 44.440 ;
        RECT 779.770 44.240 780.090 44.300 ;
        RECT 1888.370 44.240 1888.690 44.300 ;
      LAYER via ;
        RECT 779.800 44.240 780.060 44.500 ;
        RECT 1888.400 44.240 1888.660 44.500 ;
      LAYER met2 ;
        RECT 781.530 400.250 781.810 404.000 ;
        RECT 781.240 400.110 781.810 400.250 ;
        RECT 781.240 391.410 781.380 400.110 ;
        RECT 781.530 400.000 781.810 400.110 ;
        RECT 779.860 391.270 781.380 391.410 ;
        RECT 779.860 44.530 780.000 391.270 ;
        RECT 779.800 44.210 780.060 44.530 ;
        RECT 1888.400 44.210 1888.660 44.530 ;
        RECT 1888.460 2.400 1888.600 44.210 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 786.670 48.180 786.990 48.240 ;
        RECT 1905.850 48.180 1906.170 48.240 ;
        RECT 786.670 48.040 1906.170 48.180 ;
        RECT 786.670 47.980 786.990 48.040 ;
        RECT 1905.850 47.980 1906.170 48.040 ;
      LAYER via ;
        RECT 786.700 47.980 786.960 48.240 ;
        RECT 1905.880 47.980 1906.140 48.240 ;
      LAYER met2 ;
        RECT 787.050 400.250 787.330 404.000 ;
        RECT 786.760 400.110 787.330 400.250 ;
        RECT 786.760 48.270 786.900 400.110 ;
        RECT 787.050 400.000 787.330 400.110 ;
        RECT 786.700 47.950 786.960 48.270 ;
        RECT 1905.880 47.950 1906.140 48.270 ;
        RECT 1905.940 2.400 1906.080 47.950 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.130 376.280 787.450 376.340 ;
        RECT 791.270 376.280 791.590 376.340 ;
        RECT 787.130 376.140 791.590 376.280 ;
        RECT 787.130 376.080 787.450 376.140 ;
        RECT 791.270 376.080 791.590 376.140 ;
        RECT 787.130 47.840 787.450 47.900 ;
        RECT 1923.790 47.840 1924.110 47.900 ;
        RECT 787.130 47.700 1924.110 47.840 ;
        RECT 787.130 47.640 787.450 47.700 ;
        RECT 1923.790 47.640 1924.110 47.700 ;
      LAYER via ;
        RECT 787.160 376.080 787.420 376.340 ;
        RECT 791.300 376.080 791.560 376.340 ;
        RECT 787.160 47.640 787.420 47.900 ;
        RECT 1923.820 47.640 1924.080 47.900 ;
      LAYER met2 ;
        RECT 792.570 400.250 792.850 404.000 ;
        RECT 791.360 400.110 792.850 400.250 ;
        RECT 791.360 376.370 791.500 400.110 ;
        RECT 792.570 400.000 792.850 400.110 ;
        RECT 787.160 376.050 787.420 376.370 ;
        RECT 791.300 376.050 791.560 376.370 ;
        RECT 787.220 47.930 787.360 376.050 ;
        RECT 787.160 47.610 787.420 47.930 ;
        RECT 1923.820 47.610 1924.080 47.930 ;
        RECT 1923.880 2.400 1924.020 47.610 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 793.570 376.280 793.890 376.340 ;
        RECT 796.790 376.280 797.110 376.340 ;
        RECT 793.570 376.140 797.110 376.280 ;
        RECT 793.570 376.080 793.890 376.140 ;
        RECT 796.790 376.080 797.110 376.140 ;
        RECT 793.570 47.500 793.890 47.560 ;
        RECT 1941.270 47.500 1941.590 47.560 ;
        RECT 793.570 47.360 1941.590 47.500 ;
        RECT 793.570 47.300 793.890 47.360 ;
        RECT 1941.270 47.300 1941.590 47.360 ;
      LAYER via ;
        RECT 793.600 376.080 793.860 376.340 ;
        RECT 796.820 376.080 797.080 376.340 ;
        RECT 793.600 47.300 793.860 47.560 ;
        RECT 1941.300 47.300 1941.560 47.560 ;
      LAYER met2 ;
        RECT 798.090 400.250 798.370 404.000 ;
        RECT 796.880 400.110 798.370 400.250 ;
        RECT 796.880 376.370 797.020 400.110 ;
        RECT 798.090 400.000 798.370 400.110 ;
        RECT 793.600 376.050 793.860 376.370 ;
        RECT 796.820 376.050 797.080 376.370 ;
        RECT 793.660 47.590 793.800 376.050 ;
        RECT 793.600 47.270 793.860 47.590 ;
        RECT 1941.300 47.270 1941.560 47.590 ;
        RECT 1941.360 2.400 1941.500 47.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.470 47.160 800.790 47.220 ;
        RECT 1959.210 47.160 1959.530 47.220 ;
        RECT 800.470 47.020 1959.530 47.160 ;
        RECT 800.470 46.960 800.790 47.020 ;
        RECT 1959.210 46.960 1959.530 47.020 ;
      LAYER via ;
        RECT 800.500 46.960 800.760 47.220 ;
        RECT 1959.240 46.960 1959.500 47.220 ;
      LAYER met2 ;
        RECT 803.610 400.250 803.890 404.000 ;
        RECT 802.400 400.110 803.890 400.250 ;
        RECT 802.400 351.970 802.540 400.110 ;
        RECT 803.610 400.000 803.890 400.110 ;
        RECT 800.560 351.830 802.540 351.970 ;
        RECT 800.560 47.250 800.700 351.830 ;
        RECT 800.500 46.930 800.760 47.250 ;
        RECT 1959.240 46.930 1959.500 47.250 ;
        RECT 1959.300 2.400 1959.440 46.930 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.370 398.380 807.690 398.440 ;
        RECT 808.290 398.380 808.610 398.440 ;
        RECT 807.370 398.240 808.610 398.380 ;
        RECT 807.370 398.180 807.690 398.240 ;
        RECT 808.290 398.180 808.610 398.240 ;
        RECT 807.370 46.820 807.690 46.880 ;
        RECT 1976.690 46.820 1977.010 46.880 ;
        RECT 807.370 46.680 1977.010 46.820 ;
        RECT 807.370 46.620 807.690 46.680 ;
        RECT 1976.690 46.620 1977.010 46.680 ;
      LAYER via ;
        RECT 807.400 398.180 807.660 398.440 ;
        RECT 808.320 398.180 808.580 398.440 ;
        RECT 807.400 46.620 807.660 46.880 ;
        RECT 1976.720 46.620 1976.980 46.880 ;
      LAYER met2 ;
        RECT 809.130 400.250 809.410 404.000 ;
        RECT 808.380 400.110 809.410 400.250 ;
        RECT 808.380 398.470 808.520 400.110 ;
        RECT 809.130 400.000 809.410 400.110 ;
        RECT 807.400 398.150 807.660 398.470 ;
        RECT 808.320 398.150 808.580 398.470 ;
        RECT 807.460 46.910 807.600 398.150 ;
        RECT 807.400 46.590 807.660 46.910 ;
        RECT 1976.720 46.590 1976.980 46.910 ;
        RECT 1976.780 2.400 1976.920 46.590 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.270 46.480 814.590 46.540 ;
        RECT 1994.630 46.480 1994.950 46.540 ;
        RECT 814.270 46.340 1994.950 46.480 ;
        RECT 814.270 46.280 814.590 46.340 ;
        RECT 1994.630 46.280 1994.950 46.340 ;
      LAYER via ;
        RECT 814.300 46.280 814.560 46.540 ;
        RECT 1994.660 46.280 1994.920 46.540 ;
      LAYER met2 ;
        RECT 814.650 400.250 814.930 404.000 ;
        RECT 814.360 400.110 814.930 400.250 ;
        RECT 814.360 46.570 814.500 400.110 ;
        RECT 814.650 400.000 814.930 400.110 ;
        RECT 814.300 46.250 814.560 46.570 ;
        RECT 1994.660 46.250 1994.920 46.570 ;
        RECT 1994.720 2.400 1994.860 46.250 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.730 376.280 815.050 376.340 ;
        RECT 818.410 376.280 818.730 376.340 ;
        RECT 814.730 376.140 818.730 376.280 ;
        RECT 814.730 376.080 815.050 376.140 ;
        RECT 818.410 376.080 818.730 376.140 ;
        RECT 814.730 46.140 815.050 46.200 ;
        RECT 2012.570 46.140 2012.890 46.200 ;
        RECT 814.730 46.000 2012.890 46.140 ;
        RECT 814.730 45.940 815.050 46.000 ;
        RECT 2012.570 45.940 2012.890 46.000 ;
      LAYER via ;
        RECT 814.760 376.080 815.020 376.340 ;
        RECT 818.440 376.080 818.700 376.340 ;
        RECT 814.760 45.940 815.020 46.200 ;
        RECT 2012.600 45.940 2012.860 46.200 ;
      LAYER met2 ;
        RECT 819.710 400.250 819.990 404.000 ;
        RECT 818.500 400.110 819.990 400.250 ;
        RECT 818.500 376.370 818.640 400.110 ;
        RECT 819.710 400.000 819.990 400.110 ;
        RECT 814.760 376.050 815.020 376.370 ;
        RECT 818.440 376.050 818.700 376.370 ;
        RECT 814.820 46.230 814.960 376.050 ;
        RECT 814.760 45.910 815.020 46.230 ;
        RECT 2012.600 45.910 2012.860 46.230 ;
        RECT 2012.660 2.400 2012.800 45.910 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.170 376.280 821.490 376.340 ;
        RECT 823.930 376.280 824.250 376.340 ;
        RECT 821.170 376.140 824.250 376.280 ;
        RECT 821.170 376.080 821.490 376.140 ;
        RECT 823.930 376.080 824.250 376.140 ;
        RECT 821.170 45.800 821.490 45.860 ;
        RECT 2030.050 45.800 2030.370 45.860 ;
        RECT 821.170 45.660 2030.370 45.800 ;
        RECT 821.170 45.600 821.490 45.660 ;
        RECT 2030.050 45.600 2030.370 45.660 ;
      LAYER via ;
        RECT 821.200 376.080 821.460 376.340 ;
        RECT 823.960 376.080 824.220 376.340 ;
        RECT 821.200 45.600 821.460 45.860 ;
        RECT 2030.080 45.600 2030.340 45.860 ;
      LAYER met2 ;
        RECT 825.230 400.250 825.510 404.000 ;
        RECT 824.020 400.110 825.510 400.250 ;
        RECT 824.020 376.370 824.160 400.110 ;
        RECT 825.230 400.000 825.510 400.110 ;
        RECT 821.200 376.050 821.460 376.370 ;
        RECT 823.960 376.050 824.220 376.370 ;
        RECT 821.260 45.890 821.400 376.050 ;
        RECT 821.200 45.570 821.460 45.890 ;
        RECT 2030.080 45.570 2030.340 45.890 ;
        RECT 2030.140 2.400 2030.280 45.570 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 376.280 428.190 376.340 ;
        RECT 430.630 376.280 430.950 376.340 ;
        RECT 427.870 376.140 430.950 376.280 ;
        RECT 427.870 376.080 428.190 376.140 ;
        RECT 430.630 376.080 430.950 376.140 ;
        RECT 427.870 26.760 428.190 26.820 ;
        RECT 753.090 26.760 753.410 26.820 ;
        RECT 427.870 26.620 753.410 26.760 ;
        RECT 427.870 26.560 428.190 26.620 ;
        RECT 753.090 26.560 753.410 26.620 ;
      LAYER via ;
        RECT 427.900 376.080 428.160 376.340 ;
        RECT 430.660 376.080 430.920 376.340 ;
        RECT 427.900 26.560 428.160 26.820 ;
        RECT 753.120 26.560 753.380 26.820 ;
      LAYER met2 ;
        RECT 431.930 400.250 432.210 404.000 ;
        RECT 430.720 400.110 432.210 400.250 ;
        RECT 430.720 376.370 430.860 400.110 ;
        RECT 431.930 400.000 432.210 400.110 ;
        RECT 427.900 376.050 428.160 376.370 ;
        RECT 430.660 376.050 430.920 376.370 ;
        RECT 427.960 26.850 428.100 376.050 ;
        RECT 427.900 26.530 428.160 26.850 ;
        RECT 753.120 26.530 753.380 26.850 ;
        RECT 753.180 2.400 753.320 26.530 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.070 376.280 828.390 376.340 ;
        RECT 830.370 376.280 830.690 376.340 ;
        RECT 828.070 376.140 830.690 376.280 ;
        RECT 828.070 376.080 828.390 376.140 ;
        RECT 830.370 376.080 830.690 376.140 ;
        RECT 828.070 45.460 828.390 45.520 ;
        RECT 2047.990 45.460 2048.310 45.520 ;
        RECT 828.070 45.320 2048.310 45.460 ;
        RECT 828.070 45.260 828.390 45.320 ;
        RECT 2047.990 45.260 2048.310 45.320 ;
      LAYER via ;
        RECT 828.100 376.080 828.360 376.340 ;
        RECT 830.400 376.080 830.660 376.340 ;
        RECT 828.100 45.260 828.360 45.520 ;
        RECT 2048.020 45.260 2048.280 45.520 ;
      LAYER met2 ;
        RECT 830.750 400.250 831.030 404.000 ;
        RECT 830.460 400.110 831.030 400.250 ;
        RECT 830.460 376.370 830.600 400.110 ;
        RECT 830.750 400.000 831.030 400.110 ;
        RECT 828.100 376.050 828.360 376.370 ;
        RECT 830.400 376.050 830.660 376.370 ;
        RECT 828.160 45.550 828.300 376.050 ;
        RECT 828.100 45.230 828.360 45.550 ;
        RECT 2048.020 45.230 2048.280 45.550 ;
        RECT 2048.080 2.400 2048.220 45.230 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 834.970 45.120 835.290 45.180 ;
        RECT 2065.470 45.120 2065.790 45.180 ;
        RECT 834.970 44.980 2065.790 45.120 ;
        RECT 834.970 44.920 835.290 44.980 ;
        RECT 2065.470 44.920 2065.790 44.980 ;
      LAYER via ;
        RECT 835.000 44.920 835.260 45.180 ;
        RECT 2065.500 44.920 2065.760 45.180 ;
      LAYER met2 ;
        RECT 836.270 400.250 836.550 404.000 ;
        RECT 835.060 400.110 836.550 400.250 ;
        RECT 835.060 45.210 835.200 400.110 ;
        RECT 836.270 400.000 836.550 400.110 ;
        RECT 835.000 44.890 835.260 45.210 ;
        RECT 2065.500 44.890 2065.760 45.210 ;
        RECT 2065.560 2.400 2065.700 44.890 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 841.870 44.780 842.190 44.840 ;
        RECT 2083.410 44.780 2083.730 44.840 ;
        RECT 841.870 44.640 2083.730 44.780 ;
        RECT 841.870 44.580 842.190 44.640 ;
        RECT 2083.410 44.580 2083.730 44.640 ;
      LAYER via ;
        RECT 841.900 44.580 842.160 44.840 ;
        RECT 2083.440 44.580 2083.700 44.840 ;
      LAYER met2 ;
        RECT 841.790 400.180 842.070 404.000 ;
        RECT 841.790 400.000 842.100 400.180 ;
        RECT 841.960 44.870 842.100 400.000 ;
        RECT 841.900 44.550 842.160 44.870 ;
        RECT 2083.440 44.550 2083.700 44.870 ;
        RECT 2083.500 2.400 2083.640 44.550 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.330 386.480 842.650 386.540 ;
        RECT 846.010 386.480 846.330 386.540 ;
        RECT 842.330 386.340 846.330 386.480 ;
        RECT 842.330 386.280 842.650 386.340 ;
        RECT 846.010 386.280 846.330 386.340 ;
      LAYER via ;
        RECT 842.360 386.280 842.620 386.540 ;
        RECT 846.040 386.280 846.300 386.540 ;
      LAYER met2 ;
        RECT 847.310 400.250 847.590 404.000 ;
        RECT 846.100 400.110 847.590 400.250 ;
        RECT 846.100 386.570 846.240 400.110 ;
        RECT 847.310 400.000 847.590 400.110 ;
        RECT 842.360 386.250 842.620 386.570 ;
        RECT 846.040 386.250 846.300 386.570 ;
        RECT 842.420 45.405 842.560 386.250 ;
        RECT 842.350 45.035 842.630 45.405 ;
        RECT 2100.910 45.035 2101.190 45.405 ;
        RECT 2100.980 2.400 2101.120 45.035 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
      LAYER via2 ;
        RECT 842.350 45.080 842.630 45.360 ;
        RECT 2100.910 45.080 2101.190 45.360 ;
      LAYER met3 ;
        RECT 842.325 45.370 842.655 45.385 ;
        RECT 2100.885 45.370 2101.215 45.385 ;
        RECT 842.325 45.070 2101.215 45.370 ;
        RECT 842.325 45.055 842.655 45.070 ;
        RECT 2100.885 45.055 2101.215 45.070 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 848.770 386.140 849.090 386.200 ;
        RECT 851.530 386.140 851.850 386.200 ;
        RECT 848.770 386.000 851.850 386.140 ;
        RECT 848.770 385.940 849.090 386.000 ;
        RECT 851.530 385.940 851.850 386.000 ;
      LAYER via ;
        RECT 848.800 385.940 849.060 386.200 ;
        RECT 851.560 385.940 851.820 386.200 ;
      LAYER met2 ;
        RECT 852.830 400.250 853.110 404.000 ;
        RECT 851.620 400.110 853.110 400.250 ;
        RECT 851.620 386.230 851.760 400.110 ;
        RECT 852.830 400.000 853.110 400.110 ;
        RECT 848.800 385.910 849.060 386.230 ;
        RECT 851.560 385.910 851.820 386.230 ;
        RECT 848.860 44.725 849.000 385.910 ;
        RECT 848.790 44.355 849.070 44.725 ;
        RECT 2118.850 44.355 2119.130 44.725 ;
        RECT 2118.920 2.400 2119.060 44.355 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
      LAYER via2 ;
        RECT 848.790 44.400 849.070 44.680 ;
        RECT 2118.850 44.400 2119.130 44.680 ;
      LAYER met3 ;
        RECT 848.765 44.690 849.095 44.705 ;
        RECT 2118.825 44.690 2119.155 44.705 ;
        RECT 848.765 44.390 2119.155 44.690 ;
        RECT 848.765 44.375 849.095 44.390 ;
        RECT 2118.825 44.375 2119.155 44.390 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 857.050 116.180 857.370 116.240 ;
        RECT 2132.170 116.180 2132.490 116.240 ;
        RECT 857.050 116.040 2132.490 116.180 ;
        RECT 857.050 115.980 857.370 116.040 ;
        RECT 2132.170 115.980 2132.490 116.040 ;
      LAYER via ;
        RECT 857.080 115.980 857.340 116.240 ;
        RECT 2132.200 115.980 2132.460 116.240 ;
      LAYER met2 ;
        RECT 858.350 400.250 858.630 404.000 ;
        RECT 857.140 400.110 858.630 400.250 ;
        RECT 857.140 116.270 857.280 400.110 ;
        RECT 858.350 400.000 858.630 400.110 ;
        RECT 857.080 115.950 857.340 116.270 ;
        RECT 2132.200 115.950 2132.460 116.270 ;
        RECT 2132.260 82.870 2132.400 115.950 ;
        RECT 2132.260 82.730 2134.240 82.870 ;
        RECT 2134.100 1.770 2134.240 82.730 ;
        RECT 2136.190 1.770 2136.750 2.400 ;
        RECT 2134.100 1.630 2136.750 1.770 ;
        RECT 2136.190 -4.800 2136.750 1.630 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.490 115.840 863.810 115.900 ;
        RECT 2152.870 115.840 2153.190 115.900 ;
        RECT 863.490 115.700 2153.190 115.840 ;
        RECT 863.490 115.640 863.810 115.700 ;
        RECT 2152.870 115.640 2153.190 115.700 ;
      LAYER via ;
        RECT 863.520 115.640 863.780 115.900 ;
        RECT 2152.900 115.640 2153.160 115.900 ;
      LAYER met2 ;
        RECT 863.870 400.250 864.150 404.000 ;
        RECT 863.580 400.110 864.150 400.250 ;
        RECT 863.580 115.930 863.720 400.110 ;
        RECT 863.870 400.000 864.150 400.110 ;
        RECT 863.520 115.610 863.780 115.930 ;
        RECT 2152.900 115.610 2153.160 115.930 ;
        RECT 2152.960 82.870 2153.100 115.610 ;
        RECT 2152.960 82.730 2154.480 82.870 ;
        RECT 2154.340 2.400 2154.480 82.730 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.950 115.500 864.270 115.560 ;
        RECT 2166.670 115.500 2166.990 115.560 ;
        RECT 863.950 115.360 2166.990 115.500 ;
        RECT 863.950 115.300 864.270 115.360 ;
        RECT 2166.670 115.300 2166.990 115.360 ;
      LAYER via ;
        RECT 863.980 115.300 864.240 115.560 ;
        RECT 2166.700 115.300 2166.960 115.560 ;
      LAYER met2 ;
        RECT 868.930 400.250 869.210 404.000 ;
        RECT 867.720 400.110 869.210 400.250 ;
        RECT 867.720 324.370 867.860 400.110 ;
        RECT 868.930 400.000 869.210 400.110 ;
        RECT 864.040 324.230 867.860 324.370 ;
        RECT 864.040 115.590 864.180 324.230 ;
        RECT 863.980 115.270 864.240 115.590 ;
        RECT 2166.700 115.270 2166.960 115.590 ;
        RECT 2166.760 82.870 2166.900 115.270 ;
        RECT 2166.760 82.730 2170.120 82.870 ;
        RECT 2169.980 1.770 2170.120 82.730 ;
        RECT 2172.070 1.770 2172.630 2.400 ;
        RECT 2169.980 1.630 2172.630 1.770 ;
        RECT 2172.070 -4.800 2172.630 1.630 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 870.390 115.160 870.710 115.220 ;
        RECT 2187.370 115.160 2187.690 115.220 ;
        RECT 870.390 115.020 2187.690 115.160 ;
        RECT 870.390 114.960 870.710 115.020 ;
        RECT 2187.370 114.960 2187.690 115.020 ;
      LAYER via ;
        RECT 870.420 114.960 870.680 115.220 ;
        RECT 2187.400 114.960 2187.660 115.220 ;
      LAYER met2 ;
        RECT 874.450 400.250 874.730 404.000 ;
        RECT 873.240 400.110 874.730 400.250 ;
        RECT 873.240 324.370 873.380 400.110 ;
        RECT 874.450 400.000 874.730 400.110 ;
        RECT 870.480 324.230 873.380 324.370 ;
        RECT 870.480 115.250 870.620 324.230 ;
        RECT 870.420 114.930 870.680 115.250 ;
        RECT 2187.400 114.930 2187.660 115.250 ;
        RECT 2187.460 1.770 2187.600 114.930 ;
        RECT 2189.550 1.770 2190.110 2.400 ;
        RECT 2187.460 1.630 2190.110 1.770 ;
        RECT 2189.550 -4.800 2190.110 1.630 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 877.750 114.820 878.070 114.880 ;
        RECT 2201.630 114.820 2201.950 114.880 ;
        RECT 877.750 114.680 2201.950 114.820 ;
        RECT 877.750 114.620 878.070 114.680 ;
        RECT 2201.630 114.620 2201.950 114.680 ;
        RECT 2201.630 16.900 2201.950 16.960 ;
        RECT 2207.610 16.900 2207.930 16.960 ;
        RECT 2201.630 16.760 2207.930 16.900 ;
        RECT 2201.630 16.700 2201.950 16.760 ;
        RECT 2207.610 16.700 2207.930 16.760 ;
      LAYER via ;
        RECT 877.780 114.620 878.040 114.880 ;
        RECT 2201.660 114.620 2201.920 114.880 ;
        RECT 2201.660 16.700 2201.920 16.960 ;
        RECT 2207.640 16.700 2207.900 16.960 ;
      LAYER met2 ;
        RECT 879.970 400.250 880.250 404.000 ;
        RECT 878.760 400.110 880.250 400.250 ;
        RECT 878.760 324.370 878.900 400.110 ;
        RECT 879.970 400.000 880.250 400.110 ;
        RECT 877.840 324.230 878.900 324.370 ;
        RECT 877.840 114.910 877.980 324.230 ;
        RECT 877.780 114.590 878.040 114.910 ;
        RECT 2201.660 114.590 2201.920 114.910 ;
        RECT 2201.720 16.990 2201.860 114.590 ;
        RECT 2201.660 16.670 2201.920 16.990 ;
        RECT 2207.640 16.670 2207.900 16.990 ;
        RECT 2207.700 2.400 2207.840 16.670 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.230 355.540 435.550 355.600 ;
        RECT 436.150 355.540 436.470 355.600 ;
        RECT 435.230 355.400 436.470 355.540 ;
        RECT 435.230 355.340 435.550 355.400 ;
        RECT 436.150 355.340 436.470 355.400 ;
        RECT 435.230 28.800 435.550 28.860 ;
        RECT 607.270 28.800 607.590 28.860 ;
        RECT 435.230 28.660 607.590 28.800 ;
        RECT 435.230 28.600 435.550 28.660 ;
        RECT 607.270 28.600 607.590 28.660 ;
        RECT 607.270 15.880 607.590 15.940 ;
        RECT 771.030 15.880 771.350 15.940 ;
        RECT 607.270 15.740 771.350 15.880 ;
        RECT 607.270 15.680 607.590 15.740 ;
        RECT 771.030 15.680 771.350 15.740 ;
      LAYER via ;
        RECT 435.260 355.340 435.520 355.600 ;
        RECT 436.180 355.340 436.440 355.600 ;
        RECT 435.260 28.600 435.520 28.860 ;
        RECT 607.300 28.600 607.560 28.860 ;
        RECT 607.300 15.680 607.560 15.940 ;
        RECT 771.060 15.680 771.320 15.940 ;
      LAYER met2 ;
        RECT 437.450 400.250 437.730 404.000 ;
        RECT 436.240 400.110 437.730 400.250 ;
        RECT 436.240 355.630 436.380 400.110 ;
        RECT 437.450 400.000 437.730 400.110 ;
        RECT 435.260 355.310 435.520 355.630 ;
        RECT 436.180 355.310 436.440 355.630 ;
        RECT 435.320 28.890 435.460 355.310 ;
        RECT 435.260 28.570 435.520 28.890 ;
        RECT 607.300 28.570 607.560 28.890 ;
        RECT 607.360 15.970 607.500 28.570 ;
        RECT 607.300 15.650 607.560 15.970 ;
        RECT 771.060 15.650 771.320 15.970 ;
        RECT 771.120 2.400 771.260 15.650 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 884.190 50.220 884.510 50.280 ;
        RECT 2225.090 50.220 2225.410 50.280 ;
        RECT 884.190 50.080 2225.410 50.220 ;
        RECT 884.190 50.020 884.510 50.080 ;
        RECT 2225.090 50.020 2225.410 50.080 ;
      LAYER via ;
        RECT 884.220 50.020 884.480 50.280 ;
        RECT 2225.120 50.020 2225.380 50.280 ;
      LAYER met2 ;
        RECT 885.490 400.250 885.770 404.000 ;
        RECT 884.280 400.110 885.770 400.250 ;
        RECT 884.280 50.310 884.420 400.110 ;
        RECT 885.490 400.000 885.770 400.110 ;
        RECT 884.220 49.990 884.480 50.310 ;
        RECT 2225.120 49.990 2225.380 50.310 ;
        RECT 2225.180 2.400 2225.320 49.990 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.630 50.560 890.950 50.620 ;
        RECT 2243.030 50.560 2243.350 50.620 ;
        RECT 890.630 50.420 2243.350 50.560 ;
        RECT 890.630 50.360 890.950 50.420 ;
        RECT 2243.030 50.360 2243.350 50.420 ;
      LAYER via ;
        RECT 890.660 50.360 890.920 50.620 ;
        RECT 2243.060 50.360 2243.320 50.620 ;
      LAYER met2 ;
        RECT 891.010 400.250 891.290 404.000 ;
        RECT 890.720 400.110 891.290 400.250 ;
        RECT 890.720 50.650 890.860 400.110 ;
        RECT 891.010 400.000 891.290 400.110 ;
        RECT 890.660 50.330 890.920 50.650 ;
        RECT 2243.060 50.330 2243.320 50.650 ;
        RECT 2243.120 2.400 2243.260 50.330 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 891.090 386.480 891.410 386.540 ;
        RECT 895.230 386.480 895.550 386.540 ;
        RECT 891.090 386.340 895.550 386.480 ;
        RECT 891.090 386.280 891.410 386.340 ;
        RECT 895.230 386.280 895.550 386.340 ;
        RECT 891.090 50.900 891.410 50.960 ;
        RECT 2258.210 50.900 2258.530 50.960 ;
        RECT 891.090 50.760 2258.530 50.900 ;
        RECT 891.090 50.700 891.410 50.760 ;
        RECT 2258.210 50.700 2258.530 50.760 ;
      LAYER via ;
        RECT 891.120 386.280 891.380 386.540 ;
        RECT 895.260 386.280 895.520 386.540 ;
        RECT 891.120 50.700 891.380 50.960 ;
        RECT 2258.240 50.700 2258.500 50.960 ;
      LAYER met2 ;
        RECT 896.530 400.250 896.810 404.000 ;
        RECT 895.320 400.110 896.810 400.250 ;
        RECT 895.320 386.570 895.460 400.110 ;
        RECT 896.530 400.000 896.810 400.110 ;
        RECT 891.120 386.250 891.380 386.570 ;
        RECT 895.260 386.250 895.520 386.570 ;
        RECT 891.180 50.990 891.320 386.250 ;
        RECT 891.120 50.670 891.380 50.990 ;
        RECT 2258.240 50.670 2258.500 50.990 ;
        RECT 2258.300 1.770 2258.440 50.670 ;
        RECT 2260.390 1.770 2260.950 2.400 ;
        RECT 2258.300 1.630 2260.950 1.770 ;
        RECT 2260.390 -4.800 2260.950 1.630 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.530 385.800 897.850 385.860 ;
        RECT 900.750 385.800 901.070 385.860 ;
        RECT 897.530 385.660 901.070 385.800 ;
        RECT 897.530 385.600 897.850 385.660 ;
        RECT 900.750 385.600 901.070 385.660 ;
        RECT 897.530 51.240 897.850 51.300 ;
        RECT 2278.450 51.240 2278.770 51.300 ;
        RECT 897.530 51.100 2278.770 51.240 ;
        RECT 897.530 51.040 897.850 51.100 ;
        RECT 2278.450 51.040 2278.770 51.100 ;
      LAYER via ;
        RECT 897.560 385.600 897.820 385.860 ;
        RECT 900.780 385.600 901.040 385.860 ;
        RECT 897.560 51.040 897.820 51.300 ;
        RECT 2278.480 51.040 2278.740 51.300 ;
      LAYER met2 ;
        RECT 902.050 400.250 902.330 404.000 ;
        RECT 900.840 400.110 902.330 400.250 ;
        RECT 900.840 385.890 900.980 400.110 ;
        RECT 902.050 400.000 902.330 400.110 ;
        RECT 897.560 385.570 897.820 385.890 ;
        RECT 900.780 385.570 901.040 385.890 ;
        RECT 897.620 51.330 897.760 385.570 ;
        RECT 897.560 51.010 897.820 51.330 ;
        RECT 2278.480 51.010 2278.740 51.330 ;
        RECT 2278.540 2.400 2278.680 51.010 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.430 386.480 904.750 386.540 ;
        RECT 906.270 386.480 906.590 386.540 ;
        RECT 904.430 386.340 906.590 386.480 ;
        RECT 904.430 386.280 904.750 386.340 ;
        RECT 906.270 386.280 906.590 386.340 ;
        RECT 904.430 54.980 904.750 55.040 ;
        RECT 2295.930 54.980 2296.250 55.040 ;
        RECT 904.430 54.840 2296.250 54.980 ;
        RECT 904.430 54.780 904.750 54.840 ;
        RECT 2295.930 54.780 2296.250 54.840 ;
      LAYER via ;
        RECT 904.460 386.280 904.720 386.540 ;
        RECT 906.300 386.280 906.560 386.540 ;
        RECT 904.460 54.780 904.720 55.040 ;
        RECT 2295.960 54.780 2296.220 55.040 ;
      LAYER met2 ;
        RECT 907.570 400.250 907.850 404.000 ;
        RECT 906.360 400.110 907.850 400.250 ;
        RECT 906.360 386.570 906.500 400.110 ;
        RECT 907.570 400.000 907.850 400.110 ;
        RECT 904.460 386.250 904.720 386.570 ;
        RECT 906.300 386.250 906.560 386.570 ;
        RECT 904.520 55.070 904.660 386.250 ;
        RECT 904.460 54.750 904.720 55.070 ;
        RECT 2295.960 54.750 2296.220 55.070 ;
        RECT 2296.020 2.400 2296.160 54.750 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.790 54.640 912.110 54.700 ;
        RECT 2311.570 54.640 2311.890 54.700 ;
        RECT 911.790 54.500 2311.890 54.640 ;
        RECT 911.790 54.440 912.110 54.500 ;
        RECT 2311.570 54.440 2311.890 54.500 ;
      LAYER via ;
        RECT 911.820 54.440 912.080 54.700 ;
        RECT 2311.600 54.440 2311.860 54.700 ;
      LAYER met2 ;
        RECT 912.630 400.250 912.910 404.000 ;
        RECT 911.880 400.110 912.910 400.250 ;
        RECT 911.880 54.730 912.020 400.110 ;
        RECT 912.630 400.000 912.910 400.110 ;
        RECT 911.820 54.410 912.080 54.730 ;
        RECT 2311.600 54.410 2311.860 54.730 ;
        RECT 2311.660 1.770 2311.800 54.410 ;
        RECT 2313.750 1.770 2314.310 2.400 ;
        RECT 2311.660 1.630 2314.310 1.770 ;
        RECT 2313.750 -4.800 2314.310 1.630 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.230 54.300 918.550 54.360 ;
        RECT 2329.050 54.300 2329.370 54.360 ;
        RECT 918.230 54.160 2329.370 54.300 ;
        RECT 918.230 54.100 918.550 54.160 ;
        RECT 2329.050 54.100 2329.370 54.160 ;
      LAYER via ;
        RECT 918.260 54.100 918.520 54.360 ;
        RECT 2329.080 54.100 2329.340 54.360 ;
      LAYER met2 ;
        RECT 918.150 400.180 918.430 404.000 ;
        RECT 918.150 400.000 918.460 400.180 ;
        RECT 918.320 54.390 918.460 400.000 ;
        RECT 918.260 54.070 918.520 54.390 ;
        RECT 2329.080 54.070 2329.340 54.390 ;
        RECT 2329.140 1.770 2329.280 54.070 ;
        RECT 2331.230 1.770 2331.790 2.400 ;
        RECT 2329.140 1.630 2331.790 1.770 ;
        RECT 2331.230 -4.800 2331.790 1.630 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.690 386.480 919.010 386.540 ;
        RECT 922.370 386.480 922.690 386.540 ;
        RECT 918.690 386.340 922.690 386.480 ;
        RECT 918.690 386.280 919.010 386.340 ;
        RECT 922.370 386.280 922.690 386.340 ;
        RECT 918.690 53.960 919.010 54.020 ;
        RECT 2349.290 53.960 2349.610 54.020 ;
        RECT 918.690 53.820 2349.610 53.960 ;
        RECT 918.690 53.760 919.010 53.820 ;
        RECT 2349.290 53.760 2349.610 53.820 ;
      LAYER via ;
        RECT 918.720 386.280 918.980 386.540 ;
        RECT 922.400 386.280 922.660 386.540 ;
        RECT 918.720 53.760 918.980 54.020 ;
        RECT 2349.320 53.760 2349.580 54.020 ;
      LAYER met2 ;
        RECT 923.670 400.250 923.950 404.000 ;
        RECT 922.460 400.110 923.950 400.250 ;
        RECT 922.460 386.570 922.600 400.110 ;
        RECT 923.670 400.000 923.950 400.110 ;
        RECT 918.720 386.250 918.980 386.570 ;
        RECT 922.400 386.250 922.660 386.570 ;
        RECT 918.780 54.050 918.920 386.250 ;
        RECT 918.720 53.730 918.980 54.050 ;
        RECT 2349.320 53.730 2349.580 54.050 ;
        RECT 2349.380 2.400 2349.520 53.730 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.130 386.140 925.450 386.200 ;
        RECT 927.890 386.140 928.210 386.200 ;
        RECT 925.130 386.000 928.210 386.140 ;
        RECT 925.130 385.940 925.450 386.000 ;
        RECT 927.890 385.940 928.210 386.000 ;
        RECT 925.130 53.620 925.450 53.680 ;
        RECT 2367.230 53.620 2367.550 53.680 ;
        RECT 925.130 53.480 2367.550 53.620 ;
        RECT 925.130 53.420 925.450 53.480 ;
        RECT 2367.230 53.420 2367.550 53.480 ;
      LAYER via ;
        RECT 925.160 385.940 925.420 386.200 ;
        RECT 927.920 385.940 928.180 386.200 ;
        RECT 925.160 53.420 925.420 53.680 ;
        RECT 2367.260 53.420 2367.520 53.680 ;
      LAYER met2 ;
        RECT 929.190 400.250 929.470 404.000 ;
        RECT 927.980 400.110 929.470 400.250 ;
        RECT 927.980 386.230 928.120 400.110 ;
        RECT 929.190 400.000 929.470 400.110 ;
        RECT 925.160 385.910 925.420 386.230 ;
        RECT 927.920 385.910 928.180 386.230 ;
        RECT 925.220 53.710 925.360 385.910 ;
        RECT 925.160 53.390 925.420 53.710 ;
        RECT 2367.260 53.390 2367.520 53.710 ;
        RECT 2367.320 2.400 2367.460 53.390 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.030 53.280 932.350 53.340 ;
        RECT 2382.410 53.280 2382.730 53.340 ;
        RECT 932.030 53.140 2382.730 53.280 ;
        RECT 932.030 53.080 932.350 53.140 ;
        RECT 2382.410 53.080 2382.730 53.140 ;
      LAYER via ;
        RECT 932.060 53.080 932.320 53.340 ;
        RECT 2382.440 53.080 2382.700 53.340 ;
      LAYER met2 ;
        RECT 934.710 400.250 934.990 404.000 ;
        RECT 933.500 400.110 934.990 400.250 ;
        RECT 933.500 351.970 933.640 400.110 ;
        RECT 934.710 400.000 934.990 400.110 ;
        RECT 932.120 351.830 933.640 351.970 ;
        RECT 932.120 53.370 932.260 351.830 ;
        RECT 932.060 53.050 932.320 53.370 ;
        RECT 2382.440 53.050 2382.700 53.370 ;
        RECT 2382.500 1.770 2382.640 53.050 ;
        RECT 2384.590 1.770 2385.150 2.400 ;
        RECT 2382.500 1.630 2385.150 1.770 ;
        RECT 2384.590 -4.800 2385.150 1.630 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 31.180 441.990 31.240 ;
        RECT 788.970 31.180 789.290 31.240 ;
        RECT 441.670 31.040 789.290 31.180 ;
        RECT 441.670 30.980 441.990 31.040 ;
        RECT 788.970 30.980 789.290 31.040 ;
      LAYER via ;
        RECT 441.700 30.980 441.960 31.240 ;
        RECT 789.000 30.980 789.260 31.240 ;
      LAYER met2 ;
        RECT 442.510 400.250 442.790 404.000 ;
        RECT 441.760 400.110 442.790 400.250 ;
        RECT 441.760 31.270 441.900 400.110 ;
        RECT 442.510 400.000 442.790 400.110 ;
        RECT 441.700 30.950 441.960 31.270 ;
        RECT 789.000 30.950 789.260 31.270 ;
        RECT 789.060 2.400 789.200 30.950 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.290 31.520 394.610 31.580 ;
        RECT 634.870 31.520 635.190 31.580 ;
        RECT 394.290 31.380 635.190 31.520 ;
        RECT 394.290 31.320 394.610 31.380 ;
        RECT 634.870 31.320 635.190 31.380 ;
      LAYER via ;
        RECT 394.320 31.320 394.580 31.580 ;
        RECT 634.900 31.320 635.160 31.580 ;
      LAYER met2 ;
        RECT 395.130 400.250 395.410 404.000 ;
        RECT 394.380 400.110 395.410 400.250 ;
        RECT 394.380 31.610 394.520 400.110 ;
        RECT 395.130 400.000 395.410 400.110 ;
        RECT 394.320 31.290 394.580 31.610 ;
        RECT 634.900 31.290 635.160 31.610 ;
        RECT 634.960 2.400 635.100 31.290 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.930 375.940 939.250 376.000 ;
        RECT 940.770 375.940 941.090 376.000 ;
        RECT 938.930 375.800 941.090 375.940 ;
        RECT 938.930 375.740 939.250 375.800 ;
        RECT 940.770 375.740 941.090 375.800 ;
        RECT 938.930 52.940 939.250 53.000 ;
        RECT 2408.630 52.940 2408.950 53.000 ;
        RECT 938.930 52.800 2408.950 52.940 ;
        RECT 938.930 52.740 939.250 52.800 ;
        RECT 2408.630 52.740 2408.950 52.800 ;
      LAYER via ;
        RECT 938.960 375.740 939.220 376.000 ;
        RECT 940.800 375.740 941.060 376.000 ;
        RECT 938.960 52.740 939.220 53.000 ;
        RECT 2408.660 52.740 2408.920 53.000 ;
      LAYER met2 ;
        RECT 942.070 400.250 942.350 404.000 ;
        RECT 940.860 400.110 942.350 400.250 ;
        RECT 940.860 376.030 941.000 400.110 ;
        RECT 942.070 400.000 942.350 400.110 ;
        RECT 938.960 375.710 939.220 376.030 ;
        RECT 940.800 375.710 941.060 376.030 ;
        RECT 939.020 53.030 939.160 375.710 ;
        RECT 938.960 52.710 939.220 53.030 ;
        RECT 2408.660 52.710 2408.920 53.030 ;
        RECT 2408.720 2.400 2408.860 52.710 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.370 375.940 945.690 376.000 ;
        RECT 947.670 375.940 947.990 376.000 ;
        RECT 945.370 375.800 947.990 375.940 ;
        RECT 945.370 375.740 945.690 375.800 ;
        RECT 947.670 375.740 947.990 375.800 ;
        RECT 945.370 52.600 945.690 52.660 ;
        RECT 2423.810 52.600 2424.130 52.660 ;
        RECT 945.370 52.460 2424.130 52.600 ;
        RECT 945.370 52.400 945.690 52.460 ;
        RECT 2423.810 52.400 2424.130 52.460 ;
      LAYER via ;
        RECT 945.400 375.740 945.660 376.000 ;
        RECT 947.700 375.740 947.960 376.000 ;
        RECT 945.400 52.400 945.660 52.660 ;
        RECT 2423.840 52.400 2424.100 52.660 ;
      LAYER met2 ;
        RECT 947.590 400.180 947.870 404.000 ;
        RECT 947.590 400.000 947.900 400.180 ;
        RECT 947.760 376.030 947.900 400.000 ;
        RECT 945.400 375.710 945.660 376.030 ;
        RECT 947.700 375.710 947.960 376.030 ;
        RECT 945.460 52.690 945.600 375.710 ;
        RECT 945.400 52.370 945.660 52.690 ;
        RECT 2423.840 52.370 2424.100 52.690 ;
        RECT 2423.900 1.770 2424.040 52.370 ;
        RECT 2425.990 1.770 2426.550 2.400 ;
        RECT 2423.900 1.630 2426.550 1.770 ;
        RECT 2425.990 -4.800 2426.550 1.630 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.270 52.260 952.590 52.320 ;
        RECT 2444.050 52.260 2444.370 52.320 ;
        RECT 952.270 52.120 2444.370 52.260 ;
        RECT 952.270 52.060 952.590 52.120 ;
        RECT 2444.050 52.060 2444.370 52.120 ;
      LAYER via ;
        RECT 952.300 52.060 952.560 52.320 ;
        RECT 2444.080 52.060 2444.340 52.320 ;
      LAYER met2 ;
        RECT 953.110 400.250 953.390 404.000 ;
        RECT 952.360 400.110 953.390 400.250 ;
        RECT 952.360 52.350 952.500 400.110 ;
        RECT 953.110 400.000 953.390 400.110 ;
        RECT 952.300 52.030 952.560 52.350 ;
        RECT 2444.080 52.030 2444.340 52.350 ;
        RECT 2444.140 2.400 2444.280 52.030 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.730 376.280 953.050 376.340 ;
        RECT 957.330 376.280 957.650 376.340 ;
        RECT 952.730 376.140 957.650 376.280 ;
        RECT 952.730 376.080 953.050 376.140 ;
        RECT 957.330 376.080 957.650 376.140 ;
        RECT 952.730 51.920 953.050 51.980 ;
        RECT 2461.530 51.920 2461.850 51.980 ;
        RECT 952.730 51.780 2461.850 51.920 ;
        RECT 952.730 51.720 953.050 51.780 ;
        RECT 2461.530 51.720 2461.850 51.780 ;
      LAYER via ;
        RECT 952.760 376.080 953.020 376.340 ;
        RECT 957.360 376.080 957.620 376.340 ;
        RECT 952.760 51.720 953.020 51.980 ;
        RECT 2461.560 51.720 2461.820 51.980 ;
      LAYER met2 ;
        RECT 958.630 400.250 958.910 404.000 ;
        RECT 957.420 400.110 958.910 400.250 ;
        RECT 957.420 376.370 957.560 400.110 ;
        RECT 958.630 400.000 958.910 400.110 ;
        RECT 952.760 376.050 953.020 376.370 ;
        RECT 957.360 376.050 957.620 376.370 ;
        RECT 952.820 52.010 952.960 376.050 ;
        RECT 952.760 51.690 953.020 52.010 ;
        RECT 2461.560 51.690 2461.820 52.010 ;
        RECT 2461.620 2.400 2461.760 51.690 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.170 375.940 959.490 376.000 ;
        RECT 962.390 375.940 962.710 376.000 ;
        RECT 959.170 375.800 962.710 375.940 ;
        RECT 959.170 375.740 959.490 375.800 ;
        RECT 962.390 375.740 962.710 375.800 ;
        RECT 959.170 51.580 959.490 51.640 ;
        RECT 2477.170 51.580 2477.490 51.640 ;
        RECT 959.170 51.440 2477.490 51.580 ;
        RECT 959.170 51.380 959.490 51.440 ;
        RECT 2477.170 51.380 2477.490 51.440 ;
      LAYER via ;
        RECT 959.200 375.740 959.460 376.000 ;
        RECT 962.420 375.740 962.680 376.000 ;
        RECT 959.200 51.380 959.460 51.640 ;
        RECT 2477.200 51.380 2477.460 51.640 ;
      LAYER met2 ;
        RECT 963.690 400.250 963.970 404.000 ;
        RECT 962.480 400.110 963.970 400.250 ;
        RECT 962.480 376.030 962.620 400.110 ;
        RECT 963.690 400.000 963.970 400.110 ;
        RECT 959.200 375.710 959.460 376.030 ;
        RECT 962.420 375.710 962.680 376.030 ;
        RECT 959.260 51.670 959.400 375.710 ;
        RECT 959.200 51.350 959.460 51.670 ;
        RECT 2477.200 51.350 2477.460 51.670 ;
        RECT 2477.260 1.770 2477.400 51.350 ;
        RECT 2479.350 1.770 2479.910 2.400 ;
        RECT 2477.260 1.630 2479.910 1.770 ;
        RECT 2479.350 -4.800 2479.910 1.630 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.210 400.250 969.490 404.000 ;
        RECT 968.000 400.110 969.490 400.250 ;
        RECT 968.000 351.970 968.140 400.110 ;
        RECT 969.210 400.000 969.490 400.110 ;
        RECT 966.620 351.830 968.140 351.970 ;
        RECT 966.620 52.205 966.760 351.830 ;
        RECT 966.550 51.835 966.830 52.205 ;
        RECT 2494.670 51.835 2494.950 52.205 ;
        RECT 2494.740 1.770 2494.880 51.835 ;
        RECT 2496.830 1.770 2497.390 2.400 ;
        RECT 2494.740 1.630 2497.390 1.770 ;
        RECT 2496.830 -4.800 2497.390 1.630 ;
      LAYER via2 ;
        RECT 966.550 51.880 966.830 52.160 ;
        RECT 2494.670 51.880 2494.950 52.160 ;
      LAYER met3 ;
        RECT 966.525 52.170 966.855 52.185 ;
        RECT 2494.645 52.170 2494.975 52.185 ;
        RECT 966.525 51.870 2494.975 52.170 ;
        RECT 966.525 51.855 966.855 51.870 ;
        RECT 2494.645 51.855 2494.975 51.870 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.730 400.250 975.010 404.000 ;
        RECT 973.980 400.110 975.010 400.250 ;
        RECT 973.980 51.525 974.120 400.110 ;
        RECT 974.730 400.000 975.010 400.110 ;
        RECT 973.910 51.155 974.190 51.525 ;
        RECT 2514.910 51.155 2515.190 51.525 ;
        RECT 2514.980 2.400 2515.120 51.155 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
      LAYER via2 ;
        RECT 973.910 51.200 974.190 51.480 ;
        RECT 2514.910 51.200 2515.190 51.480 ;
      LAYER met3 ;
        RECT 973.885 51.490 974.215 51.505 ;
        RECT 2514.885 51.490 2515.215 51.505 ;
        RECT 973.885 51.190 2515.215 51.490 ;
        RECT 973.885 51.175 974.215 51.190 ;
        RECT 2514.885 51.175 2515.215 51.190 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.790 114.480 981.110 114.540 ;
        RECT 2532.370 114.480 2532.690 114.540 ;
        RECT 980.790 114.340 2532.690 114.480 ;
        RECT 980.790 114.280 981.110 114.340 ;
        RECT 2532.370 114.280 2532.690 114.340 ;
      LAYER via ;
        RECT 980.820 114.280 981.080 114.540 ;
        RECT 2532.400 114.280 2532.660 114.540 ;
      LAYER met2 ;
        RECT 980.250 400.250 980.530 404.000 ;
        RECT 980.250 400.110 981.020 400.250 ;
        RECT 980.250 400.000 980.530 400.110 ;
        RECT 980.880 114.570 981.020 400.110 ;
        RECT 980.820 114.250 981.080 114.570 ;
        RECT 2532.400 114.250 2532.660 114.570 ;
        RECT 2532.460 2.400 2532.600 114.250 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 981.250 114.140 981.570 114.200 ;
        RECT 2546.170 114.140 2546.490 114.200 ;
        RECT 981.250 114.000 2546.490 114.140 ;
        RECT 981.250 113.940 981.570 114.000 ;
        RECT 2546.170 113.940 2546.490 114.000 ;
      LAYER via ;
        RECT 981.280 113.940 981.540 114.200 ;
        RECT 2546.200 113.940 2546.460 114.200 ;
      LAYER met2 ;
        RECT 985.770 400.250 986.050 404.000 ;
        RECT 984.560 400.110 986.050 400.250 ;
        RECT 984.560 324.370 984.700 400.110 ;
        RECT 985.770 400.000 986.050 400.110 ;
        RECT 981.340 324.230 984.700 324.370 ;
        RECT 981.340 114.230 981.480 324.230 ;
        RECT 981.280 113.910 981.540 114.230 ;
        RECT 2546.200 113.910 2546.460 114.230 ;
        RECT 2546.260 82.870 2546.400 113.910 ;
        RECT 2546.260 82.730 2548.240 82.870 ;
        RECT 2548.100 1.770 2548.240 82.730 ;
        RECT 2550.190 1.770 2550.750 2.400 ;
        RECT 2548.100 1.630 2550.750 1.770 ;
        RECT 2550.190 -4.800 2550.750 1.630 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 988.150 113.800 988.470 113.860 ;
        RECT 2566.870 113.800 2567.190 113.860 ;
        RECT 988.150 113.660 2567.190 113.800 ;
        RECT 988.150 113.600 988.470 113.660 ;
        RECT 2566.870 113.600 2567.190 113.660 ;
      LAYER via ;
        RECT 988.180 113.600 988.440 113.860 ;
        RECT 2566.900 113.600 2567.160 113.860 ;
      LAYER met2 ;
        RECT 991.290 400.250 991.570 404.000 ;
        RECT 990.080 400.110 991.570 400.250 ;
        RECT 990.080 324.370 990.220 400.110 ;
        RECT 991.290 400.000 991.570 400.110 ;
        RECT 988.240 324.230 990.220 324.370 ;
        RECT 988.240 113.890 988.380 324.230 ;
        RECT 988.180 113.570 988.440 113.890 ;
        RECT 2566.900 113.570 2567.160 113.890 ;
        RECT 2566.960 1.770 2567.100 113.570 ;
        RECT 2567.670 1.770 2568.230 2.400 ;
        RECT 2566.960 1.630 2568.230 1.770 ;
        RECT 2567.670 -4.800 2568.230 1.630 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 30.840 448.890 30.900 ;
        RECT 812.430 30.840 812.750 30.900 ;
        RECT 448.570 30.700 812.750 30.840 ;
        RECT 448.570 30.640 448.890 30.700 ;
        RECT 812.430 30.640 812.750 30.700 ;
      LAYER via ;
        RECT 448.600 30.640 448.860 30.900 ;
        RECT 812.460 30.640 812.720 30.900 ;
      LAYER met2 ;
        RECT 449.870 400.250 450.150 404.000 ;
        RECT 448.660 400.110 450.150 400.250 ;
        RECT 448.660 30.930 448.800 400.110 ;
        RECT 449.870 400.000 450.150 400.110 ;
        RECT 448.600 30.610 448.860 30.930 ;
        RECT 812.460 30.610 812.720 30.930 ;
        RECT 812.520 2.400 812.660 30.610 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.810 400.250 997.090 404.000 ;
        RECT 995.600 400.110 997.090 400.250 ;
        RECT 995.600 324.370 995.740 400.110 ;
        RECT 996.810 400.000 997.090 400.110 ;
        RECT 994.680 324.230 995.740 324.370 ;
        RECT 994.680 113.405 994.820 324.230 ;
        RECT 994.610 113.035 994.890 113.405 ;
        RECT 2580.690 113.035 2580.970 113.405 ;
        RECT 2580.760 82.870 2580.900 113.035 ;
        RECT 2580.760 82.730 2585.960 82.870 ;
        RECT 2585.820 2.400 2585.960 82.730 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
      LAYER via2 ;
        RECT 994.610 113.080 994.890 113.360 ;
        RECT 2580.690 113.080 2580.970 113.360 ;
      LAYER met3 ;
        RECT 994.585 113.370 994.915 113.385 ;
        RECT 2580.665 113.370 2580.995 113.385 ;
        RECT 994.585 113.070 2580.995 113.370 ;
        RECT 994.585 113.055 994.915 113.070 ;
        RECT 2580.665 113.055 2580.995 113.070 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.490 57.360 1001.810 57.420 ;
        RECT 2601.370 57.360 2601.690 57.420 ;
        RECT 1001.490 57.220 2601.690 57.360 ;
        RECT 1001.490 57.160 1001.810 57.220 ;
        RECT 2601.370 57.160 2601.690 57.220 ;
      LAYER via ;
        RECT 1001.520 57.160 1001.780 57.420 ;
        RECT 2601.400 57.160 2601.660 57.420 ;
      LAYER met2 ;
        RECT 1002.330 400.250 1002.610 404.000 ;
        RECT 1001.580 400.110 1002.610 400.250 ;
        RECT 1001.580 57.450 1001.720 400.110 ;
        RECT 1002.330 400.000 1002.610 400.110 ;
        RECT 1001.520 57.130 1001.780 57.450 ;
        RECT 2601.400 57.130 2601.660 57.450 ;
        RECT 2601.460 1.770 2601.600 57.130 ;
        RECT 2603.550 1.770 2604.110 2.400 ;
        RECT 2601.460 1.630 2604.110 1.770 ;
        RECT 2603.550 -4.800 2604.110 1.630 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1008.390 57.700 1008.710 57.760 ;
        RECT 2618.850 57.700 2619.170 57.760 ;
        RECT 1008.390 57.560 2619.170 57.700 ;
        RECT 1008.390 57.500 1008.710 57.560 ;
        RECT 2618.850 57.500 2619.170 57.560 ;
      LAYER via ;
        RECT 1008.420 57.500 1008.680 57.760 ;
        RECT 2618.880 57.500 2619.140 57.760 ;
      LAYER met2 ;
        RECT 1007.390 400.250 1007.670 404.000 ;
        RECT 1007.390 400.110 1008.620 400.250 ;
        RECT 1007.390 400.000 1007.670 400.110 ;
        RECT 1008.480 57.790 1008.620 400.110 ;
        RECT 1008.420 57.470 1008.680 57.790 ;
        RECT 2618.880 57.470 2619.140 57.790 ;
        RECT 2618.940 1.770 2619.080 57.470 ;
        RECT 2621.030 1.770 2621.590 2.400 ;
        RECT 2618.940 1.630 2621.590 1.770 ;
        RECT 2621.030 -4.800 2621.590 1.630 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.930 376.280 1008.250 376.340 ;
        RECT 1011.610 376.280 1011.930 376.340 ;
        RECT 1007.930 376.140 1011.930 376.280 ;
        RECT 1007.930 376.080 1008.250 376.140 ;
        RECT 1011.610 376.080 1011.930 376.140 ;
        RECT 1007.930 58.040 1008.250 58.100 ;
        RECT 2639.090 58.040 2639.410 58.100 ;
        RECT 1007.930 57.900 2639.410 58.040 ;
        RECT 1007.930 57.840 1008.250 57.900 ;
        RECT 2639.090 57.840 2639.410 57.900 ;
      LAYER via ;
        RECT 1007.960 376.080 1008.220 376.340 ;
        RECT 1011.640 376.080 1011.900 376.340 ;
        RECT 1007.960 57.840 1008.220 58.100 ;
        RECT 2639.120 57.840 2639.380 58.100 ;
      LAYER met2 ;
        RECT 1012.910 400.250 1013.190 404.000 ;
        RECT 1011.700 400.110 1013.190 400.250 ;
        RECT 1011.700 376.370 1011.840 400.110 ;
        RECT 1012.910 400.000 1013.190 400.110 ;
        RECT 1007.960 376.050 1008.220 376.370 ;
        RECT 1011.640 376.050 1011.900 376.370 ;
        RECT 1008.020 58.130 1008.160 376.050 ;
        RECT 1007.960 57.810 1008.220 58.130 ;
        RECT 2639.120 57.810 2639.380 58.130 ;
        RECT 2639.180 2.400 2639.320 57.810 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.830 376.280 1015.150 376.340 ;
        RECT 1017.130 376.280 1017.450 376.340 ;
        RECT 1014.830 376.140 1017.450 376.280 ;
        RECT 1014.830 376.080 1015.150 376.140 ;
        RECT 1017.130 376.080 1017.450 376.140 ;
        RECT 1014.830 58.380 1015.150 58.440 ;
        RECT 2657.030 58.380 2657.350 58.440 ;
        RECT 1014.830 58.240 2657.350 58.380 ;
        RECT 1014.830 58.180 1015.150 58.240 ;
        RECT 2657.030 58.180 2657.350 58.240 ;
      LAYER via ;
        RECT 1014.860 376.080 1015.120 376.340 ;
        RECT 1017.160 376.080 1017.420 376.340 ;
        RECT 1014.860 58.180 1015.120 58.440 ;
        RECT 2657.060 58.180 2657.320 58.440 ;
      LAYER met2 ;
        RECT 1018.430 400.250 1018.710 404.000 ;
        RECT 1017.220 400.110 1018.710 400.250 ;
        RECT 1017.220 376.370 1017.360 400.110 ;
        RECT 1018.430 400.000 1018.710 400.110 ;
        RECT 1014.860 376.050 1015.120 376.370 ;
        RECT 1017.160 376.050 1017.420 376.370 ;
        RECT 1014.920 58.470 1015.060 376.050 ;
        RECT 1014.860 58.150 1015.120 58.470 ;
        RECT 2657.060 58.150 2657.320 58.470 ;
        RECT 2657.120 16.730 2657.260 58.150 ;
        RECT 2656.660 16.590 2657.260 16.730 ;
        RECT 2656.660 2.400 2656.800 16.590 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.190 62.120 1022.510 62.180 ;
        RECT 2672.210 62.120 2672.530 62.180 ;
        RECT 1022.190 61.980 2672.530 62.120 ;
        RECT 1022.190 61.920 1022.510 61.980 ;
        RECT 2672.210 61.920 2672.530 61.980 ;
      LAYER via ;
        RECT 1022.220 61.920 1022.480 62.180 ;
        RECT 2672.240 61.920 2672.500 62.180 ;
      LAYER met2 ;
        RECT 1023.950 400.250 1024.230 404.000 ;
        RECT 1022.740 400.110 1024.230 400.250 ;
        RECT 1022.740 351.970 1022.880 400.110 ;
        RECT 1023.950 400.000 1024.230 400.110 ;
        RECT 1022.280 351.830 1022.880 351.970 ;
        RECT 1022.280 62.210 1022.420 351.830 ;
        RECT 1022.220 61.890 1022.480 62.210 ;
        RECT 2672.240 61.890 2672.500 62.210 ;
        RECT 2672.300 1.770 2672.440 61.890 ;
        RECT 2674.390 1.770 2674.950 2.400 ;
        RECT 2672.300 1.630 2674.950 1.770 ;
        RECT 2674.390 -4.800 2674.950 1.630 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.630 61.780 1028.950 61.840 ;
        RECT 2691.070 61.780 2691.390 61.840 ;
        RECT 1028.630 61.640 2691.390 61.780 ;
        RECT 1028.630 61.580 1028.950 61.640 ;
        RECT 2691.070 61.580 2691.390 61.640 ;
      LAYER via ;
        RECT 1028.660 61.580 1028.920 61.840 ;
        RECT 2691.100 61.580 2691.360 61.840 ;
      LAYER met2 ;
        RECT 1029.470 400.250 1029.750 404.000 ;
        RECT 1028.720 400.110 1029.750 400.250 ;
        RECT 1028.720 61.870 1028.860 400.110 ;
        RECT 1029.470 400.000 1029.750 400.110 ;
        RECT 1028.660 61.550 1028.920 61.870 ;
        RECT 2691.100 61.550 2691.360 61.870 ;
        RECT 2691.160 1.770 2691.300 61.550 ;
        RECT 2691.870 1.770 2692.430 2.400 ;
        RECT 2691.160 1.630 2692.430 1.770 ;
        RECT 2691.870 -4.800 2692.430 1.630 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.530 61.440 1035.850 61.500 ;
        RECT 2709.930 61.440 2710.250 61.500 ;
        RECT 1035.530 61.300 2710.250 61.440 ;
        RECT 1035.530 61.240 1035.850 61.300 ;
        RECT 2709.930 61.240 2710.250 61.300 ;
      LAYER via ;
        RECT 1035.560 61.240 1035.820 61.500 ;
        RECT 2709.960 61.240 2710.220 61.500 ;
      LAYER met2 ;
        RECT 1034.990 400.250 1035.270 404.000 ;
        RECT 1034.990 400.110 1035.760 400.250 ;
        RECT 1034.990 400.000 1035.270 400.110 ;
        RECT 1035.620 61.530 1035.760 400.110 ;
        RECT 1035.560 61.210 1035.820 61.530 ;
        RECT 2709.960 61.210 2710.220 61.530 ;
        RECT 2710.020 2.400 2710.160 61.210 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.990 376.280 1036.310 376.340 ;
        RECT 1039.210 376.280 1039.530 376.340 ;
        RECT 1035.990 376.140 1039.530 376.280 ;
        RECT 1035.990 376.080 1036.310 376.140 ;
        RECT 1039.210 376.080 1039.530 376.140 ;
        RECT 1035.990 61.100 1036.310 61.160 ;
        RECT 2727.410 61.100 2727.730 61.160 ;
        RECT 1035.990 60.960 2727.730 61.100 ;
        RECT 1035.990 60.900 1036.310 60.960 ;
        RECT 2727.410 60.900 2727.730 60.960 ;
      LAYER via ;
        RECT 1036.020 376.080 1036.280 376.340 ;
        RECT 1039.240 376.080 1039.500 376.340 ;
        RECT 1036.020 60.900 1036.280 61.160 ;
        RECT 2727.440 60.900 2727.700 61.160 ;
      LAYER met2 ;
        RECT 1040.510 400.250 1040.790 404.000 ;
        RECT 1039.300 400.110 1040.790 400.250 ;
        RECT 1039.300 376.370 1039.440 400.110 ;
        RECT 1040.510 400.000 1040.790 400.110 ;
        RECT 1036.020 376.050 1036.280 376.370 ;
        RECT 1039.240 376.050 1039.500 376.370 ;
        RECT 1036.080 61.190 1036.220 376.050 ;
        RECT 1036.020 60.870 1036.280 61.190 ;
        RECT 2727.440 60.870 2727.700 61.190 ;
        RECT 2727.500 2.400 2727.640 60.870 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.430 376.620 1042.750 376.680 ;
        RECT 1044.730 376.620 1045.050 376.680 ;
        RECT 1042.430 376.480 1045.050 376.620 ;
        RECT 1042.430 376.420 1042.750 376.480 ;
        RECT 1044.730 376.420 1045.050 376.480 ;
        RECT 1042.430 60.760 1042.750 60.820 ;
        RECT 2743.050 60.760 2743.370 60.820 ;
        RECT 1042.430 60.620 2743.370 60.760 ;
        RECT 1042.430 60.560 1042.750 60.620 ;
        RECT 2743.050 60.560 2743.370 60.620 ;
      LAYER via ;
        RECT 1042.460 376.420 1042.720 376.680 ;
        RECT 1044.760 376.420 1045.020 376.680 ;
        RECT 1042.460 60.560 1042.720 60.820 ;
        RECT 2743.080 60.560 2743.340 60.820 ;
      LAYER met2 ;
        RECT 1046.030 400.250 1046.310 404.000 ;
        RECT 1044.820 400.110 1046.310 400.250 ;
        RECT 1044.820 376.710 1044.960 400.110 ;
        RECT 1046.030 400.000 1046.310 400.110 ;
        RECT 1042.460 376.390 1042.720 376.710 ;
        RECT 1044.760 376.390 1045.020 376.710 ;
        RECT 1042.520 60.850 1042.660 376.390 ;
        RECT 1042.460 60.530 1042.720 60.850 ;
        RECT 2743.080 60.530 2743.340 60.850 ;
        RECT 2743.140 1.770 2743.280 60.530 ;
        RECT 2745.230 1.770 2745.790 2.400 ;
        RECT 2743.140 1.630 2745.790 1.770 ;
        RECT 2745.230 -4.800 2745.790 1.630 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.930 29.140 456.250 29.200 ;
        RECT 630.270 29.140 630.590 29.200 ;
        RECT 455.930 29.000 630.590 29.140 ;
        RECT 455.930 28.940 456.250 29.000 ;
        RECT 630.270 28.940 630.590 29.000 ;
        RECT 630.270 20.640 630.590 20.700 ;
        RECT 830.370 20.640 830.690 20.700 ;
        RECT 630.270 20.500 830.690 20.640 ;
        RECT 630.270 20.440 630.590 20.500 ;
        RECT 830.370 20.440 830.690 20.500 ;
      LAYER via ;
        RECT 455.960 28.940 456.220 29.200 ;
        RECT 630.300 28.940 630.560 29.200 ;
        RECT 630.300 20.440 630.560 20.700 ;
        RECT 830.400 20.440 830.660 20.700 ;
      LAYER met2 ;
        RECT 455.390 400.250 455.670 404.000 ;
        RECT 455.390 400.110 456.160 400.250 ;
        RECT 455.390 400.000 455.670 400.110 ;
        RECT 456.020 29.230 456.160 400.110 ;
        RECT 455.960 28.910 456.220 29.230 ;
        RECT 630.300 28.910 630.560 29.230 ;
        RECT 630.360 20.730 630.500 28.910 ;
        RECT 630.300 20.410 630.560 20.730 ;
        RECT 830.400 20.410 830.660 20.730 ;
        RECT 830.460 2.400 830.600 20.410 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.790 60.420 1050.110 60.480 ;
        RECT 2763.290 60.420 2763.610 60.480 ;
        RECT 1049.790 60.280 2763.610 60.420 ;
        RECT 1049.790 60.220 1050.110 60.280 ;
        RECT 2763.290 60.220 2763.610 60.280 ;
      LAYER via ;
        RECT 1049.820 60.220 1050.080 60.480 ;
        RECT 2763.320 60.220 2763.580 60.480 ;
      LAYER met2 ;
        RECT 1051.550 400.250 1051.830 404.000 ;
        RECT 1050.340 400.110 1051.830 400.250 ;
        RECT 1050.340 398.210 1050.480 400.110 ;
        RECT 1051.550 400.000 1051.830 400.110 ;
        RECT 1049.880 398.070 1050.480 398.210 ;
        RECT 1049.880 60.510 1050.020 398.070 ;
        RECT 1049.820 60.190 1050.080 60.510 ;
        RECT 2763.320 60.190 2763.580 60.510 ;
        RECT 2763.380 2.400 2763.520 60.190 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1056.230 60.080 1056.550 60.140 ;
        RECT 2781.230 60.080 2781.550 60.140 ;
        RECT 1056.230 59.940 2781.550 60.080 ;
        RECT 1056.230 59.880 1056.550 59.940 ;
        RECT 2781.230 59.880 2781.550 59.940 ;
      LAYER via ;
        RECT 1056.260 59.880 1056.520 60.140 ;
        RECT 2781.260 59.880 2781.520 60.140 ;
      LAYER met2 ;
        RECT 1056.610 400.250 1056.890 404.000 ;
        RECT 1056.320 400.110 1056.890 400.250 ;
        RECT 1056.320 60.170 1056.460 400.110 ;
        RECT 1056.610 400.000 1056.890 400.110 ;
        RECT 1056.260 59.850 1056.520 60.170 ;
        RECT 2781.260 59.850 2781.520 60.170 ;
        RECT 2781.320 16.730 2781.460 59.850 ;
        RECT 2780.860 16.590 2781.460 16.730 ;
        RECT 2780.860 2.400 2781.000 16.590 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.770 376.280 1056.090 376.340 ;
        RECT 1060.830 376.280 1061.150 376.340 ;
        RECT 1055.770 376.140 1061.150 376.280 ;
        RECT 1055.770 376.080 1056.090 376.140 ;
        RECT 1060.830 376.080 1061.150 376.140 ;
        RECT 1055.770 59.740 1056.090 59.800 ;
        RECT 2796.410 59.740 2796.730 59.800 ;
        RECT 1055.770 59.600 2796.730 59.740 ;
        RECT 1055.770 59.540 1056.090 59.600 ;
        RECT 2796.410 59.540 2796.730 59.600 ;
      LAYER via ;
        RECT 1055.800 376.080 1056.060 376.340 ;
        RECT 1060.860 376.080 1061.120 376.340 ;
        RECT 1055.800 59.540 1056.060 59.800 ;
        RECT 2796.440 59.540 2796.700 59.800 ;
      LAYER met2 ;
        RECT 1062.130 400.250 1062.410 404.000 ;
        RECT 1060.920 400.110 1062.410 400.250 ;
        RECT 1060.920 376.370 1061.060 400.110 ;
        RECT 1062.130 400.000 1062.410 400.110 ;
        RECT 1055.800 376.050 1056.060 376.370 ;
        RECT 1060.860 376.050 1061.120 376.370 ;
        RECT 1055.860 59.830 1056.000 376.050 ;
        RECT 1055.800 59.510 1056.060 59.830 ;
        RECT 2796.440 59.510 2796.700 59.830 ;
        RECT 2796.500 1.770 2796.640 59.510 ;
        RECT 2798.590 1.770 2799.150 2.400 ;
        RECT 2796.500 1.630 2799.150 1.770 ;
        RECT 2798.590 -4.800 2799.150 1.630 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1062.670 376.280 1062.990 376.340 ;
        RECT 1066.350 376.280 1066.670 376.340 ;
        RECT 1062.670 376.140 1066.670 376.280 ;
        RECT 1062.670 376.080 1062.990 376.140 ;
        RECT 1066.350 376.080 1066.670 376.140 ;
        RECT 1062.670 59.400 1062.990 59.460 ;
        RECT 2815.270 59.400 2815.590 59.460 ;
        RECT 1062.670 59.260 2815.590 59.400 ;
        RECT 1062.670 59.200 1062.990 59.260 ;
        RECT 2815.270 59.200 2815.590 59.260 ;
      LAYER via ;
        RECT 1062.700 376.080 1062.960 376.340 ;
        RECT 1066.380 376.080 1066.640 376.340 ;
        RECT 1062.700 59.200 1062.960 59.460 ;
        RECT 2815.300 59.200 2815.560 59.460 ;
      LAYER met2 ;
        RECT 1067.650 400.250 1067.930 404.000 ;
        RECT 1066.440 400.110 1067.930 400.250 ;
        RECT 1066.440 376.370 1066.580 400.110 ;
        RECT 1067.650 400.000 1067.930 400.110 ;
        RECT 1062.700 376.050 1062.960 376.370 ;
        RECT 1066.380 376.050 1066.640 376.370 ;
        RECT 1062.760 59.490 1062.900 376.050 ;
        RECT 1062.700 59.170 1062.960 59.490 ;
        RECT 2815.300 59.170 2815.560 59.490 ;
        RECT 2815.360 1.770 2815.500 59.170 ;
        RECT 2816.070 1.770 2816.630 2.400 ;
        RECT 2815.360 1.630 2816.630 1.770 ;
        RECT 2816.070 -4.800 2816.630 1.630 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.570 375.940 1069.890 376.000 ;
        RECT 1071.870 375.940 1072.190 376.000 ;
        RECT 1069.570 375.800 1072.190 375.940 ;
        RECT 1069.570 375.740 1069.890 375.800 ;
        RECT 1071.870 375.740 1072.190 375.800 ;
        RECT 1069.570 59.060 1069.890 59.120 ;
        RECT 2834.130 59.060 2834.450 59.120 ;
        RECT 1069.570 58.920 2834.450 59.060 ;
        RECT 1069.570 58.860 1069.890 58.920 ;
        RECT 2834.130 58.860 2834.450 58.920 ;
      LAYER via ;
        RECT 1069.600 375.740 1069.860 376.000 ;
        RECT 1071.900 375.740 1072.160 376.000 ;
        RECT 1069.600 58.860 1069.860 59.120 ;
        RECT 2834.160 58.860 2834.420 59.120 ;
      LAYER met2 ;
        RECT 1073.170 400.250 1073.450 404.000 ;
        RECT 1071.960 400.110 1073.450 400.250 ;
        RECT 1071.960 376.030 1072.100 400.110 ;
        RECT 1073.170 400.000 1073.450 400.110 ;
        RECT 1069.600 375.710 1069.860 376.030 ;
        RECT 1071.900 375.710 1072.160 376.030 ;
        RECT 1069.660 59.150 1069.800 375.710 ;
        RECT 1069.600 58.830 1069.860 59.150 ;
        RECT 2834.160 58.830 2834.420 59.150 ;
        RECT 2834.220 2.400 2834.360 58.830 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.690 400.250 1078.970 404.000 ;
        RECT 1077.480 400.110 1078.970 400.250 ;
        RECT 1077.480 59.005 1077.620 400.110 ;
        RECT 1078.690 400.000 1078.970 400.110 ;
        RECT 1077.410 58.635 1077.690 59.005 ;
        RECT 2851.630 58.635 2851.910 59.005 ;
        RECT 2851.700 2.400 2851.840 58.635 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
      LAYER via2 ;
        RECT 1077.410 58.680 1077.690 58.960 ;
        RECT 2851.630 58.680 2851.910 58.960 ;
      LAYER met3 ;
        RECT 1077.385 58.970 1077.715 58.985 ;
        RECT 2851.605 58.970 2851.935 58.985 ;
        RECT 1077.385 58.670 2851.935 58.970 ;
        RECT 1077.385 58.655 1077.715 58.670 ;
        RECT 2851.605 58.655 2851.935 58.670 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1083.830 58.720 1084.150 58.780 ;
        RECT 2867.250 58.720 2867.570 58.780 ;
        RECT 1083.830 58.580 2867.570 58.720 ;
        RECT 1083.830 58.520 1084.150 58.580 ;
        RECT 2867.250 58.520 2867.570 58.580 ;
      LAYER via ;
        RECT 1083.860 58.520 1084.120 58.780 ;
        RECT 2867.280 58.520 2867.540 58.780 ;
      LAYER met2 ;
        RECT 1084.210 400.250 1084.490 404.000 ;
        RECT 1083.920 400.110 1084.490 400.250 ;
        RECT 1083.920 58.810 1084.060 400.110 ;
        RECT 1084.210 400.000 1084.490 400.110 ;
        RECT 1083.860 58.490 1084.120 58.810 ;
        RECT 2867.280 58.490 2867.540 58.810 ;
        RECT 2867.340 1.770 2867.480 58.490 ;
        RECT 2869.430 1.770 2869.990 2.400 ;
        RECT 2867.340 1.630 2869.990 1.770 ;
        RECT 2869.430 -4.800 2869.990 1.630 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.290 386.480 1084.610 386.540 ;
        RECT 1088.430 386.480 1088.750 386.540 ;
        RECT 1084.290 386.340 1088.750 386.480 ;
        RECT 1084.290 386.280 1084.610 386.340 ;
        RECT 1088.430 386.280 1088.750 386.340 ;
      LAYER via ;
        RECT 1084.320 386.280 1084.580 386.540 ;
        RECT 1088.460 386.280 1088.720 386.540 ;
      LAYER met2 ;
        RECT 1089.730 400.250 1090.010 404.000 ;
        RECT 1088.520 400.110 1090.010 400.250 ;
        RECT 1088.520 386.570 1088.660 400.110 ;
        RECT 1089.730 400.000 1090.010 400.110 ;
        RECT 1084.320 386.250 1084.580 386.570 ;
        RECT 1088.460 386.250 1088.720 386.570 ;
        RECT 1084.380 58.325 1084.520 386.250 ;
        RECT 1084.310 57.955 1084.590 58.325 ;
        RECT 2884.750 57.955 2885.030 58.325 ;
        RECT 2884.820 1.770 2884.960 57.955 ;
        RECT 2886.910 1.770 2887.470 2.400 ;
        RECT 2884.820 1.630 2887.470 1.770 ;
        RECT 2886.910 -4.800 2887.470 1.630 ;
      LAYER via2 ;
        RECT 1084.310 58.000 1084.590 58.280 ;
        RECT 2884.750 58.000 2885.030 58.280 ;
      LAYER met3 ;
        RECT 1084.285 58.290 1084.615 58.305 ;
        RECT 2884.725 58.290 2885.055 58.305 ;
        RECT 1084.285 57.990 2885.055 58.290 ;
        RECT 1084.285 57.975 1084.615 57.990 ;
        RECT 2884.725 57.975 2885.055 57.990 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 376.280 455.790 376.340 ;
        RECT 459.610 376.280 459.930 376.340 ;
        RECT 455.470 376.140 459.930 376.280 ;
        RECT 455.470 376.080 455.790 376.140 ;
        RECT 459.610 376.080 459.930 376.140 ;
        RECT 455.470 31.860 455.790 31.920 ;
        RECT 655.570 31.860 655.890 31.920 ;
        RECT 455.470 31.720 655.890 31.860 ;
        RECT 455.470 31.660 455.790 31.720 ;
        RECT 655.570 31.660 655.890 31.720 ;
        RECT 655.570 16.900 655.890 16.960 ;
        RECT 847.850 16.900 848.170 16.960 ;
        RECT 655.570 16.760 848.170 16.900 ;
        RECT 655.570 16.700 655.890 16.760 ;
        RECT 847.850 16.700 848.170 16.760 ;
      LAYER via ;
        RECT 455.500 376.080 455.760 376.340 ;
        RECT 459.640 376.080 459.900 376.340 ;
        RECT 455.500 31.660 455.760 31.920 ;
        RECT 655.600 31.660 655.860 31.920 ;
        RECT 655.600 16.700 655.860 16.960 ;
        RECT 847.880 16.700 848.140 16.960 ;
      LAYER met2 ;
        RECT 460.910 400.250 461.190 404.000 ;
        RECT 459.700 400.110 461.190 400.250 ;
        RECT 459.700 376.370 459.840 400.110 ;
        RECT 460.910 400.000 461.190 400.110 ;
        RECT 455.500 376.050 455.760 376.370 ;
        RECT 459.640 376.050 459.900 376.370 ;
        RECT 455.560 31.950 455.700 376.050 ;
        RECT 455.500 31.630 455.760 31.950 ;
        RECT 655.600 31.630 655.860 31.950 ;
        RECT 655.660 16.990 655.800 31.630 ;
        RECT 655.600 16.670 655.860 16.990 ;
        RECT 847.880 16.670 848.140 16.990 ;
        RECT 847.940 2.400 848.080 16.670 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 400.080 463.610 400.140 ;
        RECT 465.130 400.080 465.450 400.140 ;
        RECT 463.290 399.940 465.450 400.080 ;
        RECT 463.290 399.880 463.610 399.940 ;
        RECT 465.130 399.880 465.450 399.940 ;
        RECT 462.830 40.700 463.150 40.760 ;
        RECT 662.470 40.700 662.790 40.760 ;
        RECT 462.830 40.560 662.790 40.700 ;
        RECT 462.830 40.500 463.150 40.560 ;
        RECT 662.470 40.500 662.790 40.560 ;
        RECT 662.470 20.300 662.790 20.360 ;
        RECT 865.790 20.300 866.110 20.360 ;
        RECT 662.470 20.160 866.110 20.300 ;
        RECT 662.470 20.100 662.790 20.160 ;
        RECT 865.790 20.100 866.110 20.160 ;
      LAYER via ;
        RECT 463.320 399.880 463.580 400.140 ;
        RECT 465.160 399.880 465.420 400.140 ;
        RECT 462.860 40.500 463.120 40.760 ;
        RECT 662.500 40.500 662.760 40.760 ;
        RECT 662.500 20.100 662.760 20.360 ;
        RECT 865.820 20.100 866.080 20.360 ;
      LAYER met2 ;
        RECT 466.430 400.250 466.710 404.000 ;
        RECT 465.220 400.170 466.710 400.250 ;
        RECT 463.320 399.850 463.580 400.170 ;
        RECT 465.160 400.110 466.710 400.170 ;
        RECT 465.160 399.850 465.420 400.110 ;
        RECT 466.430 400.000 466.710 400.110 ;
        RECT 463.380 398.210 463.520 399.850 ;
        RECT 462.920 398.070 463.520 398.210 ;
        RECT 462.920 40.790 463.060 398.070 ;
        RECT 462.860 40.470 463.120 40.790 ;
        RECT 662.500 40.470 662.760 40.790 ;
        RECT 662.560 20.390 662.700 40.470 ;
        RECT 662.500 20.070 662.760 20.390 ;
        RECT 865.820 20.070 866.080 20.390 ;
        RECT 865.880 2.400 866.020 20.070 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 40.360 469.590 40.420 ;
        RECT 679.030 40.360 679.350 40.420 ;
        RECT 469.270 40.220 679.350 40.360 ;
        RECT 469.270 40.160 469.590 40.220 ;
        RECT 679.030 40.160 679.350 40.220 ;
        RECT 679.030 19.620 679.350 19.680 ;
        RECT 883.270 19.620 883.590 19.680 ;
        RECT 679.030 19.480 883.590 19.620 ;
        RECT 679.030 19.420 679.350 19.480 ;
        RECT 883.270 19.420 883.590 19.480 ;
      LAYER via ;
        RECT 469.300 40.160 469.560 40.420 ;
        RECT 679.060 40.160 679.320 40.420 ;
        RECT 679.060 19.420 679.320 19.680 ;
        RECT 883.300 19.420 883.560 19.680 ;
      LAYER met2 ;
        RECT 471.950 400.250 472.230 404.000 ;
        RECT 470.740 400.110 472.230 400.250 ;
        RECT 470.740 351.970 470.880 400.110 ;
        RECT 471.950 400.000 472.230 400.110 ;
        RECT 469.360 351.830 470.880 351.970 ;
        RECT 469.360 40.450 469.500 351.830 ;
        RECT 469.300 40.130 469.560 40.450 ;
        RECT 679.060 40.130 679.320 40.450 ;
        RECT 679.120 19.710 679.260 40.130 ;
        RECT 679.060 19.390 679.320 19.710 ;
        RECT 883.300 19.390 883.560 19.710 ;
        RECT 883.360 2.400 883.500 19.390 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.630 52.260 476.950 52.320 ;
        RECT 901.210 52.260 901.530 52.320 ;
        RECT 476.630 52.120 901.530 52.260 ;
        RECT 476.630 52.060 476.950 52.120 ;
        RECT 901.210 52.060 901.530 52.120 ;
      LAYER via ;
        RECT 476.660 52.060 476.920 52.320 ;
        RECT 901.240 52.060 901.500 52.320 ;
      LAYER met2 ;
        RECT 477.470 400.250 477.750 404.000 ;
        RECT 476.720 400.110 477.750 400.250 ;
        RECT 476.720 52.350 476.860 400.110 ;
        RECT 477.470 400.000 477.750 400.110 ;
        RECT 476.660 52.030 476.920 52.350 ;
        RECT 901.240 52.030 901.500 52.350 ;
        RECT 901.300 2.400 901.440 52.030 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 390.900 483.390 390.960 ;
        RECT 483.070 390.760 500.320 390.900 ;
        RECT 483.070 390.700 483.390 390.760 ;
        RECT 500.180 390.560 500.320 390.760 ;
        RECT 500.180 390.420 517.570 390.560 ;
        RECT 517.430 389.880 517.570 390.420 ;
        RECT 517.430 389.740 518.260 389.880 ;
        RECT 518.120 389.540 518.260 389.740 ;
        RECT 631.190 389.540 631.510 389.600 ;
        RECT 518.120 389.400 631.510 389.540 ;
        RECT 631.190 389.340 631.510 389.400 ;
        RECT 631.190 23.700 631.510 23.760 ;
        RECT 918.690 23.700 919.010 23.760 ;
        RECT 631.190 23.560 919.010 23.700 ;
        RECT 631.190 23.500 631.510 23.560 ;
        RECT 918.690 23.500 919.010 23.560 ;
      LAYER via ;
        RECT 483.100 390.700 483.360 390.960 ;
        RECT 631.220 389.340 631.480 389.600 ;
        RECT 631.220 23.500 631.480 23.760 ;
        RECT 918.720 23.500 918.980 23.760 ;
      LAYER met2 ;
        RECT 482.990 400.180 483.270 404.000 ;
        RECT 482.990 400.000 483.300 400.180 ;
        RECT 483.160 390.990 483.300 400.000 ;
        RECT 483.100 390.670 483.360 390.990 ;
        RECT 631.220 389.310 631.480 389.630 ;
        RECT 631.280 23.790 631.420 389.310 ;
        RECT 631.220 23.470 631.480 23.790 ;
        RECT 918.720 23.470 918.980 23.790 ;
        RECT 918.780 2.400 918.920 23.470 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 488.130 392.260 488.450 392.320 ;
        RECT 658.790 392.260 659.110 392.320 ;
        RECT 488.130 392.120 659.110 392.260 ;
        RECT 488.130 392.060 488.450 392.120 ;
        RECT 658.790 392.060 659.110 392.120 ;
        RECT 658.790 22.680 659.110 22.740 ;
        RECT 936.630 22.680 936.950 22.740 ;
        RECT 658.790 22.540 936.950 22.680 ;
        RECT 658.790 22.480 659.110 22.540 ;
        RECT 936.630 22.480 936.950 22.540 ;
      LAYER via ;
        RECT 488.160 392.060 488.420 392.320 ;
        RECT 658.820 392.060 659.080 392.320 ;
        RECT 658.820 22.480 659.080 22.740 ;
        RECT 936.660 22.480 936.920 22.740 ;
      LAYER met2 ;
        RECT 488.050 400.180 488.330 404.000 ;
        RECT 488.050 400.000 488.360 400.180 ;
        RECT 488.220 392.350 488.360 400.000 ;
        RECT 488.160 392.030 488.420 392.350 ;
        RECT 658.820 392.030 659.080 392.350 ;
        RECT 658.880 22.770 659.020 392.030 ;
        RECT 658.820 22.450 659.080 22.770 ;
        RECT 936.660 22.450 936.920 22.770 ;
        RECT 936.720 2.400 936.860 22.450 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.270 391.920 492.590 391.980 ;
        RECT 673.510 391.920 673.830 391.980 ;
        RECT 492.270 391.780 673.830 391.920 ;
        RECT 492.270 391.720 492.590 391.780 ;
        RECT 673.510 391.720 673.830 391.780 ;
        RECT 672.590 23.020 672.910 23.080 ;
        RECT 954.110 23.020 954.430 23.080 ;
        RECT 672.590 22.880 954.430 23.020 ;
        RECT 672.590 22.820 672.910 22.880 ;
        RECT 954.110 22.820 954.430 22.880 ;
      LAYER via ;
        RECT 492.300 391.720 492.560 391.980 ;
        RECT 673.540 391.720 673.800 391.980 ;
        RECT 672.620 22.820 672.880 23.080 ;
        RECT 954.140 22.820 954.400 23.080 ;
      LAYER met2 ;
        RECT 493.570 400.250 493.850 404.000 ;
        RECT 492.360 400.110 493.850 400.250 ;
        RECT 492.360 392.010 492.500 400.110 ;
        RECT 493.570 400.000 493.850 400.110 ;
        RECT 492.300 391.690 492.560 392.010 ;
        RECT 673.540 391.690 673.800 392.010 ;
        RECT 673.600 324.370 673.740 391.690 ;
        RECT 672.680 324.230 673.740 324.370 ;
        RECT 672.680 23.110 672.820 324.230 ;
        RECT 672.620 22.790 672.880 23.110 ;
        RECT 954.140 22.790 954.400 23.110 ;
        RECT 954.200 2.400 954.340 22.790 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 499.170 391.240 499.490 391.300 ;
        RECT 693.290 391.240 693.610 391.300 ;
        RECT 499.170 391.100 693.610 391.240 ;
        RECT 499.170 391.040 499.490 391.100 ;
        RECT 693.290 391.040 693.610 391.100 ;
        RECT 693.290 21.660 693.610 21.720 ;
        RECT 972.050 21.660 972.370 21.720 ;
        RECT 693.290 21.520 972.370 21.660 ;
        RECT 693.290 21.460 693.610 21.520 ;
        RECT 972.050 21.460 972.370 21.520 ;
      LAYER via ;
        RECT 499.200 391.040 499.460 391.300 ;
        RECT 693.320 391.040 693.580 391.300 ;
        RECT 693.320 21.460 693.580 21.720 ;
        RECT 972.080 21.460 972.340 21.720 ;
      LAYER met2 ;
        RECT 499.090 400.180 499.370 404.000 ;
        RECT 499.090 400.000 499.400 400.180 ;
        RECT 499.260 391.330 499.400 400.000 ;
        RECT 499.200 391.010 499.460 391.330 ;
        RECT 693.320 391.010 693.580 391.330 ;
        RECT 693.380 21.750 693.520 391.010 ;
        RECT 693.320 21.430 693.580 21.750 ;
        RECT 972.080 21.430 972.340 21.750 ;
        RECT 972.140 2.400 972.280 21.430 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 393.280 400.590 393.340 ;
        RECT 401.650 393.280 401.970 393.340 ;
        RECT 400.270 393.140 401.970 393.280 ;
        RECT 400.270 393.080 400.590 393.140 ;
        RECT 401.650 393.080 401.970 393.140 ;
        RECT 401.650 39.680 401.970 39.740 ;
        RECT 652.810 39.680 653.130 39.740 ;
        RECT 401.650 39.540 653.130 39.680 ;
        RECT 401.650 39.480 401.970 39.540 ;
        RECT 652.810 39.480 653.130 39.540 ;
      LAYER via ;
        RECT 400.300 393.080 400.560 393.340 ;
        RECT 401.680 393.080 401.940 393.340 ;
        RECT 401.680 39.480 401.940 39.740 ;
        RECT 652.840 39.480 653.100 39.740 ;
      LAYER met2 ;
        RECT 400.650 400.250 400.930 404.000 ;
        RECT 400.360 400.110 400.930 400.250 ;
        RECT 400.360 393.370 400.500 400.110 ;
        RECT 400.650 400.000 400.930 400.110 ;
        RECT 400.300 393.050 400.560 393.370 ;
        RECT 401.680 393.050 401.940 393.370 ;
        RECT 401.740 39.770 401.880 393.050 ;
        RECT 401.680 39.450 401.940 39.770 ;
        RECT 652.840 39.450 653.100 39.770 ;
        RECT 652.900 2.400 653.040 39.450 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.690 61.100 505.010 61.160 ;
        RECT 989.530 61.100 989.850 61.160 ;
        RECT 504.690 60.960 989.850 61.100 ;
        RECT 504.690 60.900 505.010 60.960 ;
        RECT 989.530 60.900 989.850 60.960 ;
      LAYER via ;
        RECT 504.720 60.900 504.980 61.160 ;
        RECT 989.560 60.900 989.820 61.160 ;
      LAYER met2 ;
        RECT 504.610 400.180 504.890 404.000 ;
        RECT 504.610 400.000 504.920 400.180 ;
        RECT 504.780 61.190 504.920 400.000 ;
        RECT 504.720 60.870 504.980 61.190 ;
        RECT 989.560 60.870 989.820 61.190 ;
        RECT 989.620 2.400 989.760 60.870 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 505.150 375.600 505.470 375.660 ;
        RECT 508.830 375.600 509.150 375.660 ;
        RECT 505.150 375.460 509.150 375.600 ;
        RECT 505.150 375.400 505.470 375.460 ;
        RECT 508.830 375.400 509.150 375.460 ;
        RECT 505.150 60.080 505.470 60.140 ;
        RECT 1009.310 60.080 1009.630 60.140 ;
        RECT 505.150 59.940 1009.630 60.080 ;
        RECT 505.150 59.880 505.470 59.940 ;
        RECT 1009.310 59.880 1009.630 59.940 ;
        RECT 1007.470 20.980 1007.790 21.040 ;
        RECT 1009.310 20.980 1009.630 21.040 ;
        RECT 1007.470 20.840 1009.630 20.980 ;
        RECT 1007.470 20.780 1007.790 20.840 ;
        RECT 1009.310 20.780 1009.630 20.840 ;
      LAYER via ;
        RECT 505.180 375.400 505.440 375.660 ;
        RECT 508.860 375.400 509.120 375.660 ;
        RECT 505.180 59.880 505.440 60.140 ;
        RECT 1009.340 59.880 1009.600 60.140 ;
        RECT 1007.500 20.780 1007.760 21.040 ;
        RECT 1009.340 20.780 1009.600 21.040 ;
      LAYER met2 ;
        RECT 510.130 400.250 510.410 404.000 ;
        RECT 508.920 400.110 510.410 400.250 ;
        RECT 508.920 375.690 509.060 400.110 ;
        RECT 510.130 400.000 510.410 400.110 ;
        RECT 505.180 375.370 505.440 375.690 ;
        RECT 508.860 375.370 509.120 375.690 ;
        RECT 505.240 60.170 505.380 375.370 ;
        RECT 505.180 59.850 505.440 60.170 ;
        RECT 1009.340 59.850 1009.600 60.170 ;
        RECT 1009.400 21.070 1009.540 59.850 ;
        RECT 1007.500 20.750 1007.760 21.070 ;
        RECT 1009.340 20.750 1009.600 21.070 ;
        RECT 1007.560 2.400 1007.700 20.750 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 59.740 511.910 59.800 ;
        RECT 1025.410 59.740 1025.730 59.800 ;
        RECT 511.590 59.600 1025.730 59.740 ;
        RECT 511.590 59.540 511.910 59.600 ;
        RECT 1025.410 59.540 1025.730 59.600 ;
      LAYER via ;
        RECT 511.620 59.540 511.880 59.800 ;
        RECT 1025.440 59.540 1025.700 59.800 ;
      LAYER met2 ;
        RECT 515.650 400.250 515.930 404.000 ;
        RECT 514.440 400.110 515.930 400.250 ;
        RECT 514.440 385.970 514.580 400.110 ;
        RECT 515.650 400.000 515.930 400.110 ;
        RECT 511.680 385.830 514.580 385.970 ;
        RECT 511.680 59.830 511.820 385.830 ;
        RECT 511.620 59.510 511.880 59.830 ;
        RECT 1025.440 59.510 1025.700 59.830 ;
        RECT 1025.500 2.400 1025.640 59.510 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 521.250 391.580 521.570 391.640 ;
        RECT 708.010 391.580 708.330 391.640 ;
        RECT 521.250 391.440 708.330 391.580 ;
        RECT 521.250 391.380 521.570 391.440 ;
        RECT 708.010 391.380 708.330 391.440 ;
        RECT 707.090 22.000 707.410 22.060 ;
        RECT 1042.890 22.000 1043.210 22.060 ;
        RECT 707.090 21.860 1043.210 22.000 ;
        RECT 707.090 21.800 707.410 21.860 ;
        RECT 1042.890 21.800 1043.210 21.860 ;
      LAYER via ;
        RECT 521.280 391.380 521.540 391.640 ;
        RECT 708.040 391.380 708.300 391.640 ;
        RECT 707.120 21.800 707.380 22.060 ;
        RECT 1042.920 21.800 1043.180 22.060 ;
      LAYER met2 ;
        RECT 521.170 400.180 521.450 404.000 ;
        RECT 521.170 400.000 521.480 400.180 ;
        RECT 521.340 391.670 521.480 400.000 ;
        RECT 521.280 391.350 521.540 391.670 ;
        RECT 708.040 391.350 708.300 391.670 ;
        RECT 708.100 324.370 708.240 391.350 ;
        RECT 707.180 324.230 708.240 324.370 ;
        RECT 707.180 22.090 707.320 324.230 ;
        RECT 707.120 21.770 707.380 22.090 ;
        RECT 1042.920 21.770 1043.180 22.090 ;
        RECT 1042.980 2.400 1043.120 21.770 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 526.770 389.880 527.090 389.940 ;
        RECT 782.990 389.880 783.310 389.940 ;
        RECT 526.770 389.740 783.310 389.880 ;
        RECT 526.770 389.680 527.090 389.740 ;
        RECT 782.990 389.680 783.310 389.740 ;
        RECT 782.990 31.520 783.310 31.580 ;
        RECT 1060.830 31.520 1061.150 31.580 ;
        RECT 782.990 31.380 1061.150 31.520 ;
        RECT 782.990 31.320 783.310 31.380 ;
        RECT 1060.830 31.320 1061.150 31.380 ;
      LAYER via ;
        RECT 526.800 389.680 527.060 389.940 ;
        RECT 783.020 389.680 783.280 389.940 ;
        RECT 783.020 31.320 783.280 31.580 ;
        RECT 1060.860 31.320 1061.120 31.580 ;
      LAYER met2 ;
        RECT 526.690 400.180 526.970 404.000 ;
        RECT 526.690 400.000 527.000 400.180 ;
        RECT 526.860 389.970 527.000 400.000 ;
        RECT 526.800 389.650 527.060 389.970 ;
        RECT 783.020 389.650 783.280 389.970 ;
        RECT 783.080 31.610 783.220 389.650 ;
        RECT 783.020 31.290 783.280 31.610 ;
        RECT 1060.860 31.290 1061.120 31.610 ;
        RECT 1060.920 2.400 1061.060 31.290 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 49.880 531.690 49.940 ;
        RECT 1077.390 49.880 1077.710 49.940 ;
        RECT 531.370 49.740 1077.710 49.880 ;
        RECT 531.370 49.680 531.690 49.740 ;
        RECT 1077.390 49.680 1077.710 49.740 ;
      LAYER via ;
        RECT 531.400 49.680 531.660 49.940 ;
        RECT 1077.420 49.680 1077.680 49.940 ;
      LAYER met2 ;
        RECT 532.210 400.250 532.490 404.000 ;
        RECT 531.460 400.110 532.490 400.250 ;
        RECT 531.460 49.970 531.600 400.110 ;
        RECT 532.210 400.000 532.490 400.110 ;
        RECT 531.400 49.650 531.660 49.970 ;
        RECT 1077.420 49.650 1077.680 49.970 ;
        RECT 1077.480 1.770 1077.620 49.650 ;
        RECT 1078.190 1.770 1078.750 2.400 ;
        RECT 1077.480 1.630 1078.750 1.770 ;
        RECT 1078.190 -4.800 1078.750 1.630 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.290 386.140 532.610 386.200 ;
        RECT 535.970 386.140 536.290 386.200 ;
        RECT 532.290 386.000 536.290 386.140 ;
        RECT 532.290 385.940 532.610 386.000 ;
        RECT 535.970 385.940 536.290 386.000 ;
        RECT 532.290 57.020 532.610 57.080 ;
        RECT 1096.250 57.020 1096.570 57.080 ;
        RECT 532.290 56.880 1096.570 57.020 ;
        RECT 532.290 56.820 532.610 56.880 ;
        RECT 1096.250 56.820 1096.570 56.880 ;
      LAYER via ;
        RECT 532.320 385.940 532.580 386.200 ;
        RECT 536.000 385.940 536.260 386.200 ;
        RECT 532.320 56.820 532.580 57.080 ;
        RECT 1096.280 56.820 1096.540 57.080 ;
      LAYER met2 ;
        RECT 537.270 400.250 537.550 404.000 ;
        RECT 536.060 400.110 537.550 400.250 ;
        RECT 536.060 386.230 536.200 400.110 ;
        RECT 537.270 400.000 537.550 400.110 ;
        RECT 532.320 385.910 532.580 386.230 ;
        RECT 536.000 385.910 536.260 386.230 ;
        RECT 532.380 57.110 532.520 385.910 ;
        RECT 532.320 56.790 532.580 57.110 ;
        RECT 1096.280 56.790 1096.540 57.110 ;
        RECT 1096.340 2.400 1096.480 56.790 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 105.300 539.510 105.360 ;
        RECT 1110.970 105.300 1111.290 105.360 ;
        RECT 539.190 105.160 1111.290 105.300 ;
        RECT 539.190 105.100 539.510 105.160 ;
        RECT 1110.970 105.100 1111.290 105.160 ;
      LAYER via ;
        RECT 539.220 105.100 539.480 105.360 ;
        RECT 1111.000 105.100 1111.260 105.360 ;
      LAYER met2 ;
        RECT 542.790 400.250 543.070 404.000 ;
        RECT 541.580 400.110 543.070 400.250 ;
        RECT 541.580 324.370 541.720 400.110 ;
        RECT 542.790 400.000 543.070 400.110 ;
        RECT 539.280 324.230 541.720 324.370 ;
        RECT 539.280 105.390 539.420 324.230 ;
        RECT 539.220 105.070 539.480 105.390 ;
        RECT 1111.000 105.070 1111.260 105.390 ;
        RECT 1111.060 82.870 1111.200 105.070 ;
        RECT 1111.060 82.730 1113.960 82.870 ;
        RECT 1113.820 2.400 1113.960 82.730 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.630 112.100 545.950 112.160 ;
        RECT 1131.670 112.100 1131.990 112.160 ;
        RECT 545.630 111.960 1131.990 112.100 ;
        RECT 545.630 111.900 545.950 111.960 ;
        RECT 1131.670 111.900 1131.990 111.960 ;
      LAYER via ;
        RECT 545.660 111.900 545.920 112.160 ;
        RECT 1131.700 111.900 1131.960 112.160 ;
      LAYER met2 ;
        RECT 548.310 400.250 548.590 404.000 ;
        RECT 547.100 400.110 548.590 400.250 ;
        RECT 547.100 324.370 547.240 400.110 ;
        RECT 548.310 400.000 548.590 400.110 ;
        RECT 545.720 324.230 547.240 324.370 ;
        RECT 545.720 112.190 545.860 324.230 ;
        RECT 545.660 111.870 545.920 112.190 ;
        RECT 1131.700 111.870 1131.960 112.190 ;
        RECT 1131.760 2.400 1131.900 111.870 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.450 112.440 553.770 112.500 ;
        RECT 1145.470 112.440 1145.790 112.500 ;
        RECT 553.450 112.300 1145.790 112.440 ;
        RECT 553.450 112.240 553.770 112.300 ;
        RECT 1145.470 112.240 1145.790 112.300 ;
      LAYER via ;
        RECT 553.480 112.240 553.740 112.500 ;
        RECT 1145.500 112.240 1145.760 112.500 ;
      LAYER met2 ;
        RECT 553.830 400.180 554.110 404.000 ;
        RECT 553.830 400.000 554.140 400.180 ;
        RECT 554.000 351.970 554.140 400.000 ;
        RECT 553.540 351.830 554.140 351.970 ;
        RECT 553.540 112.530 553.680 351.830 ;
        RECT 553.480 112.210 553.740 112.530 ;
        RECT 1145.500 112.210 1145.760 112.530 ;
        RECT 1145.560 82.870 1145.700 112.210 ;
        RECT 1145.560 82.730 1147.080 82.870 ;
        RECT 1146.940 1.770 1147.080 82.730 ;
        RECT 1149.030 1.770 1149.590 2.400 ;
        RECT 1146.940 1.630 1149.590 1.770 ;
        RECT 1149.030 -4.800 1149.590 1.630 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 401.190 376.280 401.510 376.340 ;
        RECT 404.870 376.280 405.190 376.340 ;
        RECT 401.190 376.140 405.190 376.280 ;
        RECT 401.190 376.080 401.510 376.140 ;
        RECT 404.870 376.080 405.190 376.140 ;
        RECT 401.190 39.000 401.510 39.060 ;
        RECT 670.750 39.000 671.070 39.060 ;
        RECT 401.190 38.860 671.070 39.000 ;
        RECT 401.190 38.800 401.510 38.860 ;
        RECT 670.750 38.800 671.070 38.860 ;
      LAYER via ;
        RECT 401.220 376.080 401.480 376.340 ;
        RECT 404.900 376.080 405.160 376.340 ;
        RECT 401.220 38.800 401.480 39.060 ;
        RECT 670.780 38.800 671.040 39.060 ;
      LAYER met2 ;
        RECT 406.170 400.250 406.450 404.000 ;
        RECT 404.960 400.110 406.450 400.250 ;
        RECT 404.960 376.370 405.100 400.110 ;
        RECT 406.170 400.000 406.450 400.110 ;
        RECT 401.220 376.050 401.480 376.370 ;
        RECT 404.900 376.050 405.160 376.370 ;
        RECT 401.280 39.090 401.420 376.050 ;
        RECT 401.220 38.770 401.480 39.090 ;
        RECT 670.780 38.770 671.040 39.090 ;
        RECT 670.840 2.400 670.980 38.770 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.350 376.960 560.670 377.020 ;
        RECT 561.270 376.960 561.590 377.020 ;
        RECT 560.350 376.820 561.590 376.960 ;
        RECT 560.350 376.760 560.670 376.820 ;
        RECT 561.270 376.760 561.590 376.820 ;
        RECT 560.350 112.780 560.670 112.840 ;
        RECT 1166.170 112.780 1166.490 112.840 ;
        RECT 560.350 112.640 1166.490 112.780 ;
        RECT 560.350 112.580 560.670 112.640 ;
        RECT 1166.170 112.580 1166.490 112.640 ;
      LAYER via ;
        RECT 560.380 376.760 560.640 377.020 ;
        RECT 561.300 376.760 561.560 377.020 ;
        RECT 560.380 112.580 560.640 112.840 ;
        RECT 1166.200 112.580 1166.460 112.840 ;
      LAYER met2 ;
        RECT 559.350 400.250 559.630 404.000 ;
        RECT 559.350 400.110 560.580 400.250 ;
        RECT 559.350 400.000 559.630 400.110 ;
        RECT 560.440 377.050 560.580 400.110 ;
        RECT 560.380 376.730 560.640 377.050 ;
        RECT 561.300 376.730 561.560 377.050 ;
        RECT 561.360 324.370 561.500 376.730 ;
        RECT 560.440 324.230 561.500 324.370 ;
        RECT 560.440 112.870 560.580 324.230 ;
        RECT 560.380 112.550 560.640 112.870 ;
        RECT 1166.200 112.550 1166.460 112.870 ;
        RECT 1166.260 82.870 1166.400 112.550 ;
        RECT 1166.260 82.730 1167.320 82.870 ;
        RECT 1167.180 2.400 1167.320 82.730 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.890 375.940 560.210 376.000 ;
        RECT 563.570 375.940 563.890 376.000 ;
        RECT 559.890 375.800 563.890 375.940 ;
        RECT 559.890 375.740 560.210 375.800 ;
        RECT 563.570 375.740 563.890 375.800 ;
        RECT 559.890 113.120 560.210 113.180 ;
        RECT 1179.970 113.120 1180.290 113.180 ;
        RECT 559.890 112.980 1180.290 113.120 ;
        RECT 559.890 112.920 560.210 112.980 ;
        RECT 1179.970 112.920 1180.290 112.980 ;
      LAYER via ;
        RECT 559.920 375.740 560.180 376.000 ;
        RECT 563.600 375.740 563.860 376.000 ;
        RECT 559.920 112.920 560.180 113.180 ;
        RECT 1180.000 112.920 1180.260 113.180 ;
      LAYER met2 ;
        RECT 564.870 400.250 565.150 404.000 ;
        RECT 563.660 400.110 565.150 400.250 ;
        RECT 563.660 376.030 563.800 400.110 ;
        RECT 564.870 400.000 565.150 400.110 ;
        RECT 559.920 375.710 560.180 376.030 ;
        RECT 563.600 375.710 563.860 376.030 ;
        RECT 559.980 113.210 560.120 375.710 ;
        RECT 559.920 112.890 560.180 113.210 ;
        RECT 1180.000 112.890 1180.260 113.210 ;
        RECT 1180.060 82.870 1180.200 112.890 ;
        RECT 1180.060 82.730 1182.960 82.870 ;
        RECT 1182.820 1.770 1182.960 82.730 ;
        RECT 1184.910 1.770 1185.470 2.400 ;
        RECT 1182.820 1.630 1185.470 1.770 ;
        RECT 1184.910 -4.800 1185.470 1.630 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.330 375.940 566.650 376.000 ;
        RECT 569.090 375.940 569.410 376.000 ;
        RECT 566.330 375.800 569.410 375.940 ;
        RECT 566.330 375.740 566.650 375.800 ;
        RECT 569.090 375.740 569.410 375.800 ;
        RECT 566.330 63.820 566.650 63.880 ;
        RECT 1200.670 63.820 1200.990 63.880 ;
        RECT 566.330 63.680 1200.990 63.820 ;
        RECT 566.330 63.620 566.650 63.680 ;
        RECT 1200.670 63.620 1200.990 63.680 ;
      LAYER via ;
        RECT 566.360 375.740 566.620 376.000 ;
        RECT 569.120 375.740 569.380 376.000 ;
        RECT 566.360 63.620 566.620 63.880 ;
        RECT 1200.700 63.620 1200.960 63.880 ;
      LAYER met2 ;
        RECT 570.390 400.250 570.670 404.000 ;
        RECT 569.180 400.110 570.670 400.250 ;
        RECT 569.180 376.030 569.320 400.110 ;
        RECT 570.390 400.000 570.670 400.110 ;
        RECT 566.360 375.710 566.620 376.030 ;
        RECT 569.120 375.710 569.380 376.030 ;
        RECT 566.420 63.910 566.560 375.710 ;
        RECT 566.360 63.590 566.620 63.910 ;
        RECT 1200.700 63.590 1200.960 63.910 ;
        RECT 1200.760 1.770 1200.900 63.590 ;
        RECT 1202.390 1.770 1202.950 2.400 ;
        RECT 1200.760 1.630 1202.950 1.770 ;
        RECT 1202.390 -4.800 1202.950 1.630 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.230 64.160 573.550 64.220 ;
        RECT 1214.470 64.160 1214.790 64.220 ;
        RECT 573.230 64.020 1214.790 64.160 ;
        RECT 573.230 63.960 573.550 64.020 ;
        RECT 1214.470 63.960 1214.790 64.020 ;
        RECT 1214.470 15.200 1214.790 15.260 ;
        RECT 1220.450 15.200 1220.770 15.260 ;
        RECT 1214.470 15.060 1220.770 15.200 ;
        RECT 1214.470 15.000 1214.790 15.060 ;
        RECT 1220.450 15.000 1220.770 15.060 ;
      LAYER via ;
        RECT 573.260 63.960 573.520 64.220 ;
        RECT 1214.500 63.960 1214.760 64.220 ;
        RECT 1214.500 15.000 1214.760 15.260 ;
        RECT 1220.480 15.000 1220.740 15.260 ;
      LAYER met2 ;
        RECT 575.910 400.250 576.190 404.000 ;
        RECT 574.700 400.110 576.190 400.250 ;
        RECT 574.700 351.970 574.840 400.110 ;
        RECT 575.910 400.000 576.190 400.110 ;
        RECT 573.320 351.830 574.840 351.970 ;
        RECT 573.320 64.250 573.460 351.830 ;
        RECT 573.260 63.930 573.520 64.250 ;
        RECT 1214.500 63.930 1214.760 64.250 ;
        RECT 1214.560 15.290 1214.700 63.930 ;
        RECT 1214.500 14.970 1214.760 15.290 ;
        RECT 1220.480 14.970 1220.740 15.290 ;
        RECT 1220.540 2.400 1220.680 14.970 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 64.500 580.910 64.560 ;
        RECT 1237.930 64.500 1238.250 64.560 ;
        RECT 580.590 64.360 1238.250 64.500 ;
        RECT 580.590 64.300 580.910 64.360 ;
        RECT 1237.930 64.300 1238.250 64.360 ;
      LAYER via ;
        RECT 580.620 64.300 580.880 64.560 ;
        RECT 1237.960 64.300 1238.220 64.560 ;
      LAYER met2 ;
        RECT 580.970 400.250 581.250 404.000 ;
        RECT 580.680 400.110 581.250 400.250 ;
        RECT 580.680 64.590 580.820 400.110 ;
        RECT 580.970 400.000 581.250 400.110 ;
        RECT 580.620 64.270 580.880 64.590 ;
        RECT 1237.960 64.270 1238.220 64.590 ;
        RECT 1238.020 2.400 1238.160 64.270 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.030 64.840 587.350 64.900 ;
        RECT 1256.330 64.840 1256.650 64.900 ;
        RECT 587.030 64.700 1256.650 64.840 ;
        RECT 587.030 64.640 587.350 64.700 ;
        RECT 1256.330 64.640 1256.650 64.700 ;
      LAYER via ;
        RECT 587.060 64.640 587.320 64.900 ;
        RECT 1256.360 64.640 1256.620 64.900 ;
      LAYER met2 ;
        RECT 586.490 400.250 586.770 404.000 ;
        RECT 586.490 400.110 587.260 400.250 ;
        RECT 586.490 400.000 586.770 400.110 ;
        RECT 587.120 64.930 587.260 400.110 ;
        RECT 587.060 64.610 587.320 64.930 ;
        RECT 1256.360 64.610 1256.620 64.930 ;
        RECT 1256.420 17.410 1256.560 64.610 ;
        RECT 1255.960 17.270 1256.560 17.410 ;
        RECT 1255.960 2.400 1256.100 17.270 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.490 376.280 587.810 376.340 ;
        RECT 590.710 376.280 591.030 376.340 ;
        RECT 587.490 376.140 591.030 376.280 ;
        RECT 587.490 376.080 587.810 376.140 ;
        RECT 590.710 376.080 591.030 376.140 ;
        RECT 587.490 65.180 587.810 65.240 ;
        RECT 1271.050 65.180 1271.370 65.240 ;
        RECT 587.490 65.040 1271.370 65.180 ;
        RECT 587.490 64.980 587.810 65.040 ;
        RECT 1271.050 64.980 1271.370 65.040 ;
      LAYER via ;
        RECT 587.520 376.080 587.780 376.340 ;
        RECT 590.740 376.080 591.000 376.340 ;
        RECT 587.520 64.980 587.780 65.240 ;
        RECT 1271.080 64.980 1271.340 65.240 ;
      LAYER met2 ;
        RECT 592.010 400.250 592.290 404.000 ;
        RECT 590.800 400.110 592.290 400.250 ;
        RECT 590.800 376.370 590.940 400.110 ;
        RECT 592.010 400.000 592.290 400.110 ;
        RECT 587.520 376.050 587.780 376.370 ;
        RECT 590.740 376.050 591.000 376.370 ;
        RECT 587.580 65.270 587.720 376.050 ;
        RECT 587.520 64.950 587.780 65.270 ;
        RECT 1271.080 64.950 1271.340 65.270 ;
        RECT 1271.140 1.770 1271.280 64.950 ;
        RECT 1273.230 1.770 1273.790 2.400 ;
        RECT 1271.140 1.630 1273.790 1.770 ;
        RECT 1273.230 -4.800 1273.790 1.630 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 596.230 386.480 596.550 386.540 ;
        RECT 594.020 386.340 596.550 386.480 ;
        RECT 594.020 386.200 594.160 386.340 ;
        RECT 596.230 386.280 596.550 386.340 ;
        RECT 593.930 385.940 594.250 386.200 ;
        RECT 593.930 68.920 594.250 68.980 ;
        RECT 1291.290 68.920 1291.610 68.980 ;
        RECT 593.930 68.780 1291.610 68.920 ;
        RECT 593.930 68.720 594.250 68.780 ;
        RECT 1291.290 68.720 1291.610 68.780 ;
      LAYER via ;
        RECT 596.260 386.280 596.520 386.540 ;
        RECT 593.960 385.940 594.220 386.200 ;
        RECT 593.960 68.720 594.220 68.980 ;
        RECT 1291.320 68.720 1291.580 68.980 ;
      LAYER met2 ;
        RECT 597.530 400.250 597.810 404.000 ;
        RECT 596.320 400.110 597.810 400.250 ;
        RECT 596.320 386.570 596.460 400.110 ;
        RECT 597.530 400.000 597.810 400.110 ;
        RECT 596.260 386.250 596.520 386.570 ;
        RECT 593.960 385.910 594.220 386.230 ;
        RECT 594.020 69.010 594.160 385.910 ;
        RECT 593.960 68.690 594.220 69.010 ;
        RECT 1291.320 68.690 1291.580 69.010 ;
        RECT 1291.380 2.400 1291.520 68.690 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.290 68.580 601.610 68.640 ;
        RECT 1308.770 68.580 1309.090 68.640 ;
        RECT 601.290 68.440 1309.090 68.580 ;
        RECT 601.290 68.380 601.610 68.440 ;
        RECT 1308.770 68.380 1309.090 68.440 ;
      LAYER via ;
        RECT 601.320 68.380 601.580 68.640 ;
        RECT 1308.800 68.380 1309.060 68.640 ;
      LAYER met2 ;
        RECT 603.050 400.250 603.330 404.000 ;
        RECT 601.840 400.110 603.330 400.250 ;
        RECT 601.840 386.470 601.980 400.110 ;
        RECT 603.050 400.000 603.330 400.110 ;
        RECT 601.380 386.330 601.980 386.470 ;
        RECT 601.380 68.670 601.520 386.330 ;
        RECT 601.320 68.350 601.580 68.670 ;
        RECT 1308.800 68.350 1309.060 68.670 ;
        RECT 1308.860 2.400 1309.000 68.350 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 68.240 608.050 68.300 ;
        RECT 1324.870 68.240 1325.190 68.300 ;
        RECT 607.730 68.100 1325.190 68.240 ;
        RECT 607.730 68.040 608.050 68.100 ;
        RECT 1324.870 68.040 1325.190 68.100 ;
      LAYER via ;
        RECT 607.760 68.040 608.020 68.300 ;
        RECT 1324.900 68.040 1325.160 68.300 ;
      LAYER met2 ;
        RECT 608.570 400.250 608.850 404.000 ;
        RECT 607.820 400.110 608.850 400.250 ;
        RECT 607.820 68.330 607.960 400.110 ;
        RECT 608.570 400.000 608.850 400.110 ;
        RECT 607.760 68.010 608.020 68.330 ;
        RECT 1324.900 68.010 1325.160 68.330 ;
        RECT 1324.960 1.770 1325.100 68.010 ;
        RECT 1326.590 1.770 1327.150 2.400 ;
        RECT 1324.960 1.630 1327.150 1.770 ;
        RECT 1326.590 -4.800 1327.150 1.630 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.630 398.720 407.950 398.780 ;
        RECT 410.390 398.720 410.710 398.780 ;
        RECT 407.630 398.580 410.710 398.720 ;
        RECT 407.630 398.520 407.950 398.580 ;
        RECT 410.390 398.520 410.710 398.580 ;
        RECT 407.630 38.660 407.950 38.720 ;
        RECT 688.230 38.660 688.550 38.720 ;
        RECT 407.630 38.520 688.550 38.660 ;
        RECT 407.630 38.460 407.950 38.520 ;
        RECT 688.230 38.460 688.550 38.520 ;
      LAYER via ;
        RECT 407.660 398.520 407.920 398.780 ;
        RECT 410.420 398.520 410.680 398.780 ;
        RECT 407.660 38.460 407.920 38.720 ;
        RECT 688.260 38.460 688.520 38.720 ;
      LAYER met2 ;
        RECT 411.690 400.250 411.970 404.000 ;
        RECT 410.480 400.110 411.970 400.250 ;
        RECT 410.480 398.810 410.620 400.110 ;
        RECT 411.690 400.000 411.970 400.110 ;
        RECT 407.660 398.490 407.920 398.810 ;
        RECT 410.420 398.490 410.680 398.810 ;
        RECT 407.720 38.750 407.860 398.490 ;
        RECT 407.660 38.430 407.920 38.750 ;
        RECT 688.260 38.430 688.520 38.750 ;
        RECT 688.320 2.400 688.460 38.430 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.630 67.900 614.950 67.960 ;
        RECT 1341.890 67.900 1342.210 67.960 ;
        RECT 614.630 67.760 1342.210 67.900 ;
        RECT 614.630 67.700 614.950 67.760 ;
        RECT 1341.890 67.700 1342.210 67.760 ;
      LAYER via ;
        RECT 614.660 67.700 614.920 67.960 ;
        RECT 1341.920 67.700 1342.180 67.960 ;
      LAYER met2 ;
        RECT 614.090 400.250 614.370 404.000 ;
        RECT 614.090 400.110 614.860 400.250 ;
        RECT 614.090 400.000 614.370 400.110 ;
        RECT 614.720 67.990 614.860 400.110 ;
        RECT 614.660 67.670 614.920 67.990 ;
        RECT 1341.920 67.670 1342.180 67.990 ;
        RECT 1341.980 1.770 1342.120 67.670 ;
        RECT 1344.070 1.770 1344.630 2.400 ;
        RECT 1341.980 1.630 1344.630 1.770 ;
        RECT 1344.070 -4.800 1344.630 1.630 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 386.480 614.490 386.540 ;
        RECT 618.310 386.480 618.630 386.540 ;
        RECT 614.170 386.340 618.630 386.480 ;
        RECT 614.170 386.280 614.490 386.340 ;
        RECT 618.310 386.280 618.630 386.340 ;
        RECT 614.170 67.560 614.490 67.620 ;
        RECT 1362.130 67.560 1362.450 67.620 ;
        RECT 614.170 67.420 1362.450 67.560 ;
        RECT 614.170 67.360 614.490 67.420 ;
        RECT 1362.130 67.360 1362.450 67.420 ;
      LAYER via ;
        RECT 614.200 386.280 614.460 386.540 ;
        RECT 618.340 386.280 618.600 386.540 ;
        RECT 614.200 67.360 614.460 67.620 ;
        RECT 1362.160 67.360 1362.420 67.620 ;
      LAYER met2 ;
        RECT 619.610 400.250 619.890 404.000 ;
        RECT 618.400 400.110 619.890 400.250 ;
        RECT 618.400 386.570 618.540 400.110 ;
        RECT 619.610 400.000 619.890 400.110 ;
        RECT 614.200 386.250 614.460 386.570 ;
        RECT 618.340 386.250 618.600 386.570 ;
        RECT 614.260 67.650 614.400 386.250 ;
        RECT 614.200 67.330 614.460 67.650 ;
        RECT 1362.160 67.330 1362.420 67.650 ;
        RECT 1362.220 2.400 1362.360 67.330 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 386.140 621.390 386.200 ;
        RECT 623.830 386.140 624.150 386.200 ;
        RECT 621.070 386.000 624.150 386.140 ;
        RECT 621.070 385.940 621.390 386.000 ;
        RECT 623.830 385.940 624.150 386.000 ;
        RECT 621.070 67.220 621.390 67.280 ;
        RECT 1380.530 67.220 1380.850 67.280 ;
        RECT 621.070 67.080 1380.850 67.220 ;
        RECT 621.070 67.020 621.390 67.080 ;
        RECT 1380.530 67.020 1380.850 67.080 ;
      LAYER via ;
        RECT 621.100 385.940 621.360 386.200 ;
        RECT 623.860 385.940 624.120 386.200 ;
        RECT 621.100 67.020 621.360 67.280 ;
        RECT 1380.560 67.020 1380.820 67.280 ;
      LAYER met2 ;
        RECT 625.130 400.250 625.410 404.000 ;
        RECT 623.920 400.110 625.410 400.250 ;
        RECT 623.920 386.230 624.060 400.110 ;
        RECT 625.130 400.000 625.410 400.110 ;
        RECT 621.100 385.910 621.360 386.230 ;
        RECT 623.860 385.910 624.120 386.230 ;
        RECT 621.160 67.310 621.300 385.910 ;
        RECT 621.100 66.990 621.360 67.310 ;
        RECT 1380.560 66.990 1380.820 67.310 ;
        RECT 1380.620 17.410 1380.760 66.990 ;
        RECT 1380.160 17.270 1380.760 17.410 ;
        RECT 1380.160 2.400 1380.300 17.270 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.970 387.160 628.290 387.220 ;
        RECT 629.350 387.160 629.670 387.220 ;
        RECT 627.970 387.020 629.670 387.160 ;
        RECT 627.970 386.960 628.290 387.020 ;
        RECT 629.350 386.960 629.670 387.020 ;
        RECT 627.970 66.880 628.290 66.940 ;
        RECT 1395.250 66.880 1395.570 66.940 ;
        RECT 627.970 66.740 1395.570 66.880 ;
        RECT 627.970 66.680 628.290 66.740 ;
        RECT 1395.250 66.680 1395.570 66.740 ;
      LAYER via ;
        RECT 628.000 386.960 628.260 387.220 ;
        RECT 629.380 386.960 629.640 387.220 ;
        RECT 628.000 66.680 628.260 66.940 ;
        RECT 1395.280 66.680 1395.540 66.940 ;
      LAYER met2 ;
        RECT 630.190 400.250 630.470 404.000 ;
        RECT 629.440 400.110 630.470 400.250 ;
        RECT 629.440 387.250 629.580 400.110 ;
        RECT 630.190 400.000 630.470 400.110 ;
        RECT 628.000 386.930 628.260 387.250 ;
        RECT 629.380 386.930 629.640 387.250 ;
        RECT 628.060 66.970 628.200 386.930 ;
        RECT 628.000 66.650 628.260 66.970 ;
        RECT 1395.280 66.650 1395.540 66.970 ;
        RECT 1395.340 1.770 1395.480 66.650 ;
        RECT 1397.430 1.770 1397.990 2.400 ;
        RECT 1395.340 1.630 1397.990 1.770 ;
        RECT 1397.430 -4.800 1397.990 1.630 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.870 66.540 635.190 66.600 ;
        RECT 1415.490 66.540 1415.810 66.600 ;
        RECT 634.870 66.400 1415.810 66.540 ;
        RECT 634.870 66.340 635.190 66.400 ;
        RECT 1415.490 66.340 1415.810 66.400 ;
      LAYER via ;
        RECT 634.900 66.340 635.160 66.600 ;
        RECT 1415.520 66.340 1415.780 66.600 ;
      LAYER met2 ;
        RECT 635.710 400.250 635.990 404.000 ;
        RECT 634.960 400.110 635.990 400.250 ;
        RECT 634.960 66.630 635.100 400.110 ;
        RECT 635.710 400.000 635.990 400.110 ;
        RECT 634.900 66.310 635.160 66.630 ;
        RECT 1415.520 66.310 1415.780 66.630 ;
        RECT 1415.580 2.400 1415.720 66.310 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.330 386.480 635.650 386.540 ;
        RECT 639.930 386.480 640.250 386.540 ;
        RECT 635.330 386.340 640.250 386.480 ;
        RECT 635.330 386.280 635.650 386.340 ;
        RECT 639.930 386.280 640.250 386.340 ;
        RECT 635.330 66.200 635.650 66.260 ;
        RECT 1432.970 66.200 1433.290 66.260 ;
        RECT 635.330 66.060 1433.290 66.200 ;
        RECT 635.330 66.000 635.650 66.060 ;
        RECT 1432.970 66.000 1433.290 66.060 ;
      LAYER via ;
        RECT 635.360 386.280 635.620 386.540 ;
        RECT 639.960 386.280 640.220 386.540 ;
        RECT 635.360 66.000 635.620 66.260 ;
        RECT 1433.000 66.000 1433.260 66.260 ;
      LAYER met2 ;
        RECT 641.230 400.250 641.510 404.000 ;
        RECT 640.020 400.110 641.510 400.250 ;
        RECT 640.020 386.570 640.160 400.110 ;
        RECT 641.230 400.000 641.510 400.110 ;
        RECT 635.360 386.250 635.620 386.570 ;
        RECT 639.960 386.250 640.220 386.570 ;
        RECT 635.420 66.290 635.560 386.250 ;
        RECT 635.360 65.970 635.620 66.290 ;
        RECT 1433.000 65.970 1433.260 66.290 ;
        RECT 1433.060 2.400 1433.200 65.970 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.230 386.140 642.550 386.200 ;
        RECT 645.450 386.140 645.770 386.200 ;
        RECT 642.230 386.000 645.770 386.140 ;
        RECT 642.230 385.940 642.550 386.000 ;
        RECT 645.450 385.940 645.770 386.000 ;
        RECT 642.230 65.860 642.550 65.920 ;
        RECT 1449.070 65.860 1449.390 65.920 ;
        RECT 642.230 65.720 1449.390 65.860 ;
        RECT 642.230 65.660 642.550 65.720 ;
        RECT 1449.070 65.660 1449.390 65.720 ;
      LAYER via ;
        RECT 642.260 385.940 642.520 386.200 ;
        RECT 645.480 385.940 645.740 386.200 ;
        RECT 642.260 65.660 642.520 65.920 ;
        RECT 1449.100 65.660 1449.360 65.920 ;
      LAYER met2 ;
        RECT 646.750 400.250 647.030 404.000 ;
        RECT 645.540 400.110 647.030 400.250 ;
        RECT 645.540 386.230 645.680 400.110 ;
        RECT 646.750 400.000 647.030 400.110 ;
        RECT 642.260 385.910 642.520 386.230 ;
        RECT 645.480 385.910 645.740 386.230 ;
        RECT 642.320 65.950 642.460 385.910 ;
        RECT 642.260 65.630 642.520 65.950 ;
        RECT 1449.100 65.630 1449.360 65.950 ;
        RECT 1449.160 1.770 1449.300 65.630 ;
        RECT 1450.790 1.770 1451.350 2.400 ;
        RECT 1449.160 1.630 1451.350 1.770 ;
        RECT 1450.790 -4.800 1451.350 1.630 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.130 65.520 649.450 65.580 ;
        RECT 1466.090 65.520 1466.410 65.580 ;
        RECT 649.130 65.380 1466.410 65.520 ;
        RECT 649.130 65.320 649.450 65.380 ;
        RECT 1466.090 65.320 1466.410 65.380 ;
      LAYER via ;
        RECT 649.160 65.320 649.420 65.580 ;
        RECT 1466.120 65.320 1466.380 65.580 ;
      LAYER met2 ;
        RECT 652.270 400.250 652.550 404.000 ;
        RECT 651.060 400.110 652.550 400.250 ;
        RECT 651.060 386.650 651.200 400.110 ;
        RECT 652.270 400.000 652.550 400.110 ;
        RECT 649.220 386.510 651.200 386.650 ;
        RECT 649.220 65.610 649.360 386.510 ;
        RECT 649.160 65.290 649.420 65.610 ;
        RECT 1466.120 65.290 1466.380 65.610 ;
        RECT 1466.180 1.770 1466.320 65.290 ;
        RECT 1468.270 1.770 1468.830 2.400 ;
        RECT 1466.180 1.630 1468.830 1.770 ;
        RECT 1468.270 -4.800 1468.830 1.630 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.790 400.250 658.070 404.000 ;
        RECT 656.580 400.110 658.070 400.250 ;
        RECT 656.580 65.805 656.720 400.110 ;
        RECT 657.790 400.000 658.070 400.110 ;
        RECT 656.510 65.435 656.790 65.805 ;
        RECT 1486.350 65.435 1486.630 65.805 ;
        RECT 1486.420 2.400 1486.560 65.435 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
      LAYER via2 ;
        RECT 656.510 65.480 656.790 65.760 ;
        RECT 1486.350 65.480 1486.630 65.760 ;
      LAYER met3 ;
        RECT 656.485 65.770 656.815 65.785 ;
        RECT 1486.325 65.770 1486.655 65.785 ;
        RECT 656.485 65.470 1486.655 65.770 ;
        RECT 656.485 65.455 656.815 65.470 ;
        RECT 1486.325 65.455 1486.655 65.470 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.850 113.460 664.170 113.520 ;
        RECT 1497.370 113.460 1497.690 113.520 ;
        RECT 663.850 113.320 1497.690 113.460 ;
        RECT 663.850 113.260 664.170 113.320 ;
        RECT 1497.370 113.260 1497.690 113.320 ;
        RECT 1497.370 15.200 1497.690 15.260 ;
        RECT 1503.810 15.200 1504.130 15.260 ;
        RECT 1497.370 15.060 1504.130 15.200 ;
        RECT 1497.370 15.000 1497.690 15.060 ;
        RECT 1503.810 15.000 1504.130 15.060 ;
      LAYER via ;
        RECT 663.880 113.260 664.140 113.520 ;
        RECT 1497.400 113.260 1497.660 113.520 ;
        RECT 1497.400 15.000 1497.660 15.260 ;
        RECT 1503.840 15.000 1504.100 15.260 ;
      LAYER met2 ;
        RECT 663.310 400.250 663.590 404.000 ;
        RECT 663.310 400.110 664.080 400.250 ;
        RECT 663.310 400.000 663.590 400.110 ;
        RECT 663.940 113.550 664.080 400.110 ;
        RECT 663.880 113.230 664.140 113.550 ;
        RECT 1497.400 113.230 1497.660 113.550 ;
        RECT 1497.460 15.290 1497.600 113.230 ;
        RECT 1497.400 14.970 1497.660 15.290 ;
        RECT 1503.840 14.970 1504.100 15.290 ;
        RECT 1503.900 2.400 1504.040 14.970 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.990 37.980 415.310 38.040 ;
        RECT 706.170 37.980 706.490 38.040 ;
        RECT 414.990 37.840 706.490 37.980 ;
        RECT 414.990 37.780 415.310 37.840 ;
        RECT 706.170 37.780 706.490 37.840 ;
      LAYER via ;
        RECT 415.020 37.780 415.280 38.040 ;
        RECT 706.200 37.780 706.460 38.040 ;
      LAYER met2 ;
        RECT 417.210 400.250 417.490 404.000 ;
        RECT 416.000 400.110 417.490 400.250 ;
        RECT 416.000 324.370 416.140 400.110 ;
        RECT 417.210 400.000 417.490 400.110 ;
        RECT 415.080 324.230 416.140 324.370 ;
        RECT 415.080 38.070 415.220 324.230 ;
        RECT 415.020 37.750 415.280 38.070 ;
        RECT 706.200 37.750 706.460 38.070 ;
        RECT 706.260 2.400 706.400 37.750 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 386.140 663.710 386.200 ;
        RECT 667.530 386.140 667.850 386.200 ;
        RECT 663.390 386.000 667.850 386.140 ;
        RECT 663.390 385.940 663.710 386.000 ;
        RECT 667.530 385.940 667.850 386.000 ;
        RECT 663.390 117.200 663.710 117.260 ;
        RECT 1518.070 117.200 1518.390 117.260 ;
        RECT 663.390 117.060 1518.390 117.200 ;
        RECT 663.390 117.000 663.710 117.060 ;
        RECT 1518.070 117.000 1518.390 117.060 ;
      LAYER via ;
        RECT 663.420 385.940 663.680 386.200 ;
        RECT 667.560 385.940 667.820 386.200 ;
        RECT 663.420 117.000 663.680 117.260 ;
        RECT 1518.100 117.000 1518.360 117.260 ;
      LAYER met2 ;
        RECT 668.830 400.250 669.110 404.000 ;
        RECT 667.620 400.110 669.110 400.250 ;
        RECT 667.620 386.230 667.760 400.110 ;
        RECT 668.830 400.000 669.110 400.110 ;
        RECT 663.420 385.910 663.680 386.230 ;
        RECT 667.560 385.910 667.820 386.230 ;
        RECT 663.480 117.290 663.620 385.910 ;
        RECT 663.420 116.970 663.680 117.290 ;
        RECT 1518.100 116.970 1518.360 117.290 ;
        RECT 1518.160 82.870 1518.300 116.970 ;
        RECT 1518.160 82.730 1519.680 82.870 ;
        RECT 1519.540 1.770 1519.680 82.730 ;
        RECT 1521.630 1.770 1522.190 2.400 ;
        RECT 1519.540 1.630 1522.190 1.770 ;
        RECT 1521.630 -4.800 1522.190 1.630 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.750 116.860 671.070 116.920 ;
        RECT 1538.770 116.860 1539.090 116.920 ;
        RECT 670.750 116.720 1539.090 116.860 ;
        RECT 670.750 116.660 671.070 116.720 ;
        RECT 1538.770 116.660 1539.090 116.720 ;
      LAYER via ;
        RECT 670.780 116.660 671.040 116.920 ;
        RECT 1538.800 116.660 1539.060 116.920 ;
      LAYER met2 ;
        RECT 674.350 400.250 674.630 404.000 ;
        RECT 673.140 400.110 674.630 400.250 ;
        RECT 673.140 386.470 673.280 400.110 ;
        RECT 674.350 400.000 674.630 400.110 ;
        RECT 670.840 386.330 673.280 386.470 ;
        RECT 670.840 116.950 670.980 386.330 ;
        RECT 670.780 116.630 671.040 116.950 ;
        RECT 1538.800 116.630 1539.060 116.950 ;
        RECT 1538.860 17.410 1539.000 116.630 ;
        RECT 1538.860 17.270 1539.920 17.410 ;
        RECT 1539.780 2.400 1539.920 17.270 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 677.190 118.900 677.510 118.960 ;
        RECT 1552.570 118.900 1552.890 118.960 ;
        RECT 677.190 118.760 1552.890 118.900 ;
        RECT 677.190 118.700 677.510 118.760 ;
        RECT 1552.570 118.700 1552.890 118.760 ;
      LAYER via ;
        RECT 677.220 118.700 677.480 118.960 ;
        RECT 1552.600 118.700 1552.860 118.960 ;
      LAYER met2 ;
        RECT 679.410 400.250 679.690 404.000 ;
        RECT 678.200 400.110 679.690 400.250 ;
        RECT 678.200 324.370 678.340 400.110 ;
        RECT 679.410 400.000 679.690 400.110 ;
        RECT 677.280 324.230 678.340 324.370 ;
        RECT 677.280 118.990 677.420 324.230 ;
        RECT 677.220 118.670 677.480 118.990 ;
        RECT 1552.600 118.670 1552.860 118.990 ;
        RECT 1552.660 82.870 1552.800 118.670 ;
        RECT 1552.660 82.730 1557.400 82.870 ;
        RECT 1557.260 2.400 1557.400 82.730 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.090 119.240 684.410 119.300 ;
        RECT 1573.270 119.240 1573.590 119.300 ;
        RECT 684.090 119.100 1573.590 119.240 ;
        RECT 684.090 119.040 684.410 119.100 ;
        RECT 1573.270 119.040 1573.590 119.100 ;
      LAYER via ;
        RECT 684.120 119.040 684.380 119.300 ;
        RECT 1573.300 119.040 1573.560 119.300 ;
      LAYER met2 ;
        RECT 684.930 400.250 685.210 404.000 ;
        RECT 684.180 400.110 685.210 400.250 ;
        RECT 684.180 119.330 684.320 400.110 ;
        RECT 684.930 400.000 685.210 400.110 ;
        RECT 684.120 119.010 684.380 119.330 ;
        RECT 1573.300 119.010 1573.560 119.330 ;
        RECT 1573.360 1.770 1573.500 119.010 ;
        RECT 1574.990 1.770 1575.550 2.400 ;
        RECT 1573.360 1.630 1575.550 1.770 ;
        RECT 1574.990 -4.800 1575.550 1.630 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.990 70.620 691.310 70.680 ;
        RECT 1590.290 70.620 1590.610 70.680 ;
        RECT 690.990 70.480 1590.610 70.620 ;
        RECT 690.990 70.420 691.310 70.480 ;
        RECT 1590.290 70.420 1590.610 70.480 ;
      LAYER via ;
        RECT 691.020 70.420 691.280 70.680 ;
        RECT 1590.320 70.420 1590.580 70.680 ;
      LAYER met2 ;
        RECT 690.450 400.250 690.730 404.000 ;
        RECT 690.450 400.110 691.220 400.250 ;
        RECT 690.450 400.000 690.730 400.110 ;
        RECT 691.080 70.710 691.220 400.110 ;
        RECT 691.020 70.390 691.280 70.710 ;
        RECT 1590.320 70.390 1590.580 70.710 ;
        RECT 1590.380 1.770 1590.520 70.390 ;
        RECT 1592.470 1.770 1593.030 2.400 ;
        RECT 1590.380 1.630 1593.030 1.770 ;
        RECT 1592.470 -4.800 1593.030 1.630 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.530 376.280 690.850 376.340 ;
        RECT 694.670 376.280 694.990 376.340 ;
        RECT 690.530 376.140 694.990 376.280 ;
        RECT 690.530 376.080 690.850 376.140 ;
        RECT 694.670 376.080 694.990 376.140 ;
        RECT 690.530 70.960 690.850 71.020 ;
        RECT 1610.530 70.960 1610.850 71.020 ;
        RECT 690.530 70.820 1610.850 70.960 ;
        RECT 690.530 70.760 690.850 70.820 ;
        RECT 1610.530 70.760 1610.850 70.820 ;
      LAYER via ;
        RECT 690.560 376.080 690.820 376.340 ;
        RECT 694.700 376.080 694.960 376.340 ;
        RECT 690.560 70.760 690.820 71.020 ;
        RECT 1610.560 70.760 1610.820 71.020 ;
      LAYER met2 ;
        RECT 695.970 400.250 696.250 404.000 ;
        RECT 694.760 400.110 696.250 400.250 ;
        RECT 694.760 376.370 694.900 400.110 ;
        RECT 695.970 400.000 696.250 400.110 ;
        RECT 690.560 376.050 690.820 376.370 ;
        RECT 694.700 376.050 694.960 376.370 ;
        RECT 690.620 71.050 690.760 376.050 ;
        RECT 690.560 70.730 690.820 71.050 ;
        RECT 1610.560 70.730 1610.820 71.050 ;
        RECT 1610.620 2.400 1610.760 70.730 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.430 375.940 697.750 376.000 ;
        RECT 700.190 375.940 700.510 376.000 ;
        RECT 697.430 375.800 700.510 375.940 ;
        RECT 697.430 375.740 697.750 375.800 ;
        RECT 700.190 375.740 700.510 375.800 ;
        RECT 697.430 71.300 697.750 71.360 ;
        RECT 1621.570 71.300 1621.890 71.360 ;
        RECT 697.430 71.160 1621.890 71.300 ;
        RECT 697.430 71.100 697.750 71.160 ;
        RECT 1621.570 71.100 1621.890 71.160 ;
        RECT 1621.570 15.200 1621.890 15.260 ;
        RECT 1628.010 15.200 1628.330 15.260 ;
        RECT 1621.570 15.060 1628.330 15.200 ;
        RECT 1621.570 15.000 1621.890 15.060 ;
        RECT 1628.010 15.000 1628.330 15.060 ;
      LAYER via ;
        RECT 697.460 375.740 697.720 376.000 ;
        RECT 700.220 375.740 700.480 376.000 ;
        RECT 697.460 71.100 697.720 71.360 ;
        RECT 1621.600 71.100 1621.860 71.360 ;
        RECT 1621.600 15.000 1621.860 15.260 ;
        RECT 1628.040 15.000 1628.300 15.260 ;
      LAYER met2 ;
        RECT 701.490 400.250 701.770 404.000 ;
        RECT 700.280 400.110 701.770 400.250 ;
        RECT 700.280 376.030 700.420 400.110 ;
        RECT 701.490 400.000 701.770 400.110 ;
        RECT 697.460 375.710 697.720 376.030 ;
        RECT 700.220 375.710 700.480 376.030 ;
        RECT 697.520 71.390 697.660 375.710 ;
        RECT 697.460 71.070 697.720 71.390 ;
        RECT 1621.600 71.070 1621.860 71.390 ;
        RECT 1621.660 15.290 1621.800 71.070 ;
        RECT 1621.600 14.970 1621.860 15.290 ;
        RECT 1628.040 14.970 1628.300 15.290 ;
        RECT 1628.100 2.400 1628.240 14.970 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.330 71.640 704.650 71.700 ;
        RECT 1643.650 71.640 1643.970 71.700 ;
        RECT 704.330 71.500 1643.970 71.640 ;
        RECT 704.330 71.440 704.650 71.500 ;
        RECT 1643.650 71.440 1643.970 71.500 ;
      LAYER via ;
        RECT 704.360 71.440 704.620 71.700 ;
        RECT 1643.680 71.440 1643.940 71.700 ;
      LAYER met2 ;
        RECT 707.010 400.250 707.290 404.000 ;
        RECT 705.800 400.110 707.290 400.250 ;
        RECT 705.800 399.570 705.940 400.110 ;
        RECT 707.010 400.000 707.290 400.110 ;
        RECT 704.420 399.430 705.940 399.570 ;
        RECT 704.420 71.730 704.560 399.430 ;
        RECT 704.360 71.410 704.620 71.730 ;
        RECT 1643.680 71.410 1643.940 71.730 ;
        RECT 1643.740 1.770 1643.880 71.410 ;
        RECT 1645.830 1.770 1646.390 2.400 ;
        RECT 1643.740 1.630 1646.390 1.770 ;
        RECT 1645.830 -4.800 1646.390 1.630 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.690 71.980 712.010 72.040 ;
        RECT 1663.430 71.980 1663.750 72.040 ;
        RECT 711.690 71.840 1663.750 71.980 ;
        RECT 711.690 71.780 712.010 71.840 ;
        RECT 1663.430 71.780 1663.750 71.840 ;
      LAYER via ;
        RECT 711.720 71.780 711.980 72.040 ;
        RECT 1663.460 71.780 1663.720 72.040 ;
      LAYER met2 ;
        RECT 712.530 400.250 712.810 404.000 ;
        RECT 711.780 400.110 712.810 400.250 ;
        RECT 711.780 72.070 711.920 400.110 ;
        RECT 712.530 400.000 712.810 400.110 ;
        RECT 711.720 71.750 711.980 72.070 ;
        RECT 1663.460 71.750 1663.720 72.070 ;
        RECT 1663.520 2.400 1663.660 71.750 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.130 75.720 718.450 75.780 ;
        RECT 1681.370 75.720 1681.690 75.780 ;
        RECT 718.130 75.580 1681.690 75.720 ;
        RECT 718.130 75.520 718.450 75.580 ;
        RECT 1681.370 75.520 1681.690 75.580 ;
      LAYER via ;
        RECT 718.160 75.520 718.420 75.780 ;
        RECT 1681.400 75.520 1681.660 75.780 ;
      LAYER met2 ;
        RECT 718.050 400.180 718.330 404.000 ;
        RECT 718.050 400.000 718.360 400.180 ;
        RECT 718.220 75.810 718.360 400.000 ;
        RECT 718.160 75.490 718.420 75.810 ;
        RECT 1681.400 75.490 1681.660 75.810 ;
        RECT 1681.460 2.400 1681.600 75.490 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 422.350 36.280 422.670 36.340 ;
        RECT 723.650 36.280 723.970 36.340 ;
        RECT 422.350 36.140 723.970 36.280 ;
        RECT 422.350 36.080 422.670 36.140 ;
        RECT 723.650 36.080 723.970 36.140 ;
      LAYER via ;
        RECT 422.380 36.080 422.640 36.340 ;
        RECT 723.680 36.080 723.940 36.340 ;
      LAYER met2 ;
        RECT 422.730 400.250 423.010 404.000 ;
        RECT 422.440 400.110 423.010 400.250 ;
        RECT 422.440 36.370 422.580 400.110 ;
        RECT 422.730 400.000 423.010 400.110 ;
        RECT 422.380 36.050 422.640 36.370 ;
        RECT 723.680 36.050 723.940 36.370 ;
        RECT 723.740 2.400 723.880 36.050 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.590 376.280 718.910 376.340 ;
        RECT 722.270 376.280 722.590 376.340 ;
        RECT 718.590 376.140 722.590 376.280 ;
        RECT 718.590 376.080 718.910 376.140 ;
        RECT 722.270 376.080 722.590 376.140 ;
        RECT 718.590 75.380 718.910 75.440 ;
        RECT 1697.470 75.380 1697.790 75.440 ;
        RECT 718.590 75.240 1697.790 75.380 ;
        RECT 718.590 75.180 718.910 75.240 ;
        RECT 1697.470 75.180 1697.790 75.240 ;
      LAYER via ;
        RECT 718.620 376.080 718.880 376.340 ;
        RECT 722.300 376.080 722.560 376.340 ;
        RECT 718.620 75.180 718.880 75.440 ;
        RECT 1697.500 75.180 1697.760 75.440 ;
      LAYER met2 ;
        RECT 723.110 400.250 723.390 404.000 ;
        RECT 722.360 400.110 723.390 400.250 ;
        RECT 722.360 376.370 722.500 400.110 ;
        RECT 723.110 400.000 723.390 400.110 ;
        RECT 718.620 376.050 718.880 376.370 ;
        RECT 722.300 376.050 722.560 376.370 ;
        RECT 718.680 75.470 718.820 376.050 ;
        RECT 718.620 75.150 718.880 75.470 ;
        RECT 1697.500 75.150 1697.760 75.470 ;
        RECT 1697.560 1.770 1697.700 75.150 ;
        RECT 1699.190 1.770 1699.750 2.400 ;
        RECT 1697.560 1.630 1699.750 1.770 ;
        RECT 1699.190 -4.800 1699.750 1.630 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.030 375.940 725.350 376.000 ;
        RECT 727.330 375.940 727.650 376.000 ;
        RECT 725.030 375.800 727.650 375.940 ;
        RECT 725.030 375.740 725.350 375.800 ;
        RECT 727.330 375.740 727.650 375.800 ;
        RECT 725.030 75.040 725.350 75.100 ;
        RECT 1714.490 75.040 1714.810 75.100 ;
        RECT 725.030 74.900 1714.810 75.040 ;
        RECT 725.030 74.840 725.350 74.900 ;
        RECT 1714.490 74.840 1714.810 74.900 ;
      LAYER via ;
        RECT 725.060 375.740 725.320 376.000 ;
        RECT 727.360 375.740 727.620 376.000 ;
        RECT 725.060 74.840 725.320 75.100 ;
        RECT 1714.520 74.840 1714.780 75.100 ;
      LAYER met2 ;
        RECT 728.630 400.250 728.910 404.000 ;
        RECT 727.420 400.110 728.910 400.250 ;
        RECT 727.420 376.030 727.560 400.110 ;
        RECT 728.630 400.000 728.910 400.110 ;
        RECT 725.060 375.710 725.320 376.030 ;
        RECT 727.360 375.710 727.620 376.030 ;
        RECT 725.120 75.130 725.260 375.710 ;
        RECT 725.060 74.810 725.320 75.130 ;
        RECT 1714.520 74.810 1714.780 75.130 ;
        RECT 1714.580 1.770 1714.720 74.810 ;
        RECT 1716.670 1.770 1717.230 2.400 ;
        RECT 1714.580 1.630 1717.230 1.770 ;
        RECT 1716.670 -4.800 1717.230 1.630 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.930 74.700 732.250 74.760 ;
        RECT 1734.730 74.700 1735.050 74.760 ;
        RECT 731.930 74.560 1735.050 74.700 ;
        RECT 731.930 74.500 732.250 74.560 ;
        RECT 1734.730 74.500 1735.050 74.560 ;
      LAYER via ;
        RECT 731.960 74.500 732.220 74.760 ;
        RECT 1734.760 74.500 1735.020 74.760 ;
      LAYER met2 ;
        RECT 734.150 400.250 734.430 404.000 ;
        RECT 732.940 400.110 734.430 400.250 ;
        RECT 732.940 399.570 733.080 400.110 ;
        RECT 734.150 400.000 734.430 400.110 ;
        RECT 732.020 399.430 733.080 399.570 ;
        RECT 732.020 74.790 732.160 399.430 ;
        RECT 731.960 74.470 732.220 74.790 ;
        RECT 1734.760 74.470 1735.020 74.790 ;
        RECT 1734.820 2.400 1734.960 74.470 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.370 74.360 738.690 74.420 ;
        RECT 1746.230 74.360 1746.550 74.420 ;
        RECT 738.370 74.220 1746.550 74.360 ;
        RECT 738.370 74.160 738.690 74.220 ;
        RECT 1746.230 74.160 1746.550 74.220 ;
        RECT 1746.230 15.200 1746.550 15.260 ;
        RECT 1752.210 15.200 1752.530 15.260 ;
        RECT 1746.230 15.060 1752.530 15.200 ;
        RECT 1746.230 15.000 1746.550 15.060 ;
        RECT 1752.210 15.000 1752.530 15.060 ;
      LAYER via ;
        RECT 738.400 74.160 738.660 74.420 ;
        RECT 1746.260 74.160 1746.520 74.420 ;
        RECT 1746.260 15.000 1746.520 15.260 ;
        RECT 1752.240 15.000 1752.500 15.260 ;
      LAYER met2 ;
        RECT 739.670 400.250 739.950 404.000 ;
        RECT 738.460 400.110 739.950 400.250 ;
        RECT 738.460 74.450 738.600 400.110 ;
        RECT 739.670 400.000 739.950 400.110 ;
        RECT 738.400 74.130 738.660 74.450 ;
        RECT 1746.260 74.130 1746.520 74.450 ;
        RECT 1746.320 15.290 1746.460 74.130 ;
        RECT 1746.260 14.970 1746.520 15.290 ;
        RECT 1752.240 14.970 1752.500 15.290 ;
        RECT 1752.300 2.400 1752.440 14.970 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.730 74.020 746.050 74.080 ;
        RECT 1767.850 74.020 1768.170 74.080 ;
        RECT 745.730 73.880 1768.170 74.020 ;
        RECT 745.730 73.820 746.050 73.880 ;
        RECT 1767.850 73.820 1768.170 73.880 ;
      LAYER via ;
        RECT 745.760 73.820 746.020 74.080 ;
        RECT 1767.880 73.820 1768.140 74.080 ;
      LAYER met2 ;
        RECT 745.190 400.250 745.470 404.000 ;
        RECT 745.190 400.110 745.960 400.250 ;
        RECT 745.190 400.000 745.470 400.110 ;
        RECT 745.820 74.110 745.960 400.110 ;
        RECT 745.760 73.790 746.020 74.110 ;
        RECT 1767.880 73.790 1768.140 74.110 ;
        RECT 1767.940 1.770 1768.080 73.790 ;
        RECT 1770.030 1.770 1770.590 2.400 ;
        RECT 1767.940 1.630 1770.590 1.770 ;
        RECT 1770.030 -4.800 1770.590 1.630 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.270 376.280 745.590 376.340 ;
        RECT 749.410 376.280 749.730 376.340 ;
        RECT 745.270 376.140 749.730 376.280 ;
        RECT 745.270 376.080 745.590 376.140 ;
        RECT 749.410 376.080 749.730 376.140 ;
        RECT 745.270 73.680 745.590 73.740 ;
        RECT 1787.630 73.680 1787.950 73.740 ;
        RECT 745.270 73.540 1787.950 73.680 ;
        RECT 745.270 73.480 745.590 73.540 ;
        RECT 1787.630 73.480 1787.950 73.540 ;
      LAYER via ;
        RECT 745.300 376.080 745.560 376.340 ;
        RECT 749.440 376.080 749.700 376.340 ;
        RECT 745.300 73.480 745.560 73.740 ;
        RECT 1787.660 73.480 1787.920 73.740 ;
      LAYER met2 ;
        RECT 750.710 400.250 750.990 404.000 ;
        RECT 749.500 400.110 750.990 400.250 ;
        RECT 749.500 376.370 749.640 400.110 ;
        RECT 750.710 400.000 750.990 400.110 ;
        RECT 745.300 376.050 745.560 376.370 ;
        RECT 749.440 376.050 749.700 376.370 ;
        RECT 745.360 73.770 745.500 376.050 ;
        RECT 745.300 73.450 745.560 73.770 ;
        RECT 1787.660 73.450 1787.920 73.770 ;
        RECT 1787.720 2.400 1787.860 73.450 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.170 376.280 752.490 376.340 ;
        RECT 754.930 376.280 755.250 376.340 ;
        RECT 752.170 376.140 755.250 376.280 ;
        RECT 752.170 376.080 752.490 376.140 ;
        RECT 754.930 376.080 755.250 376.140 ;
        RECT 752.170 73.340 752.490 73.400 ;
        RECT 1805.570 73.340 1805.890 73.400 ;
        RECT 752.170 73.200 1805.890 73.340 ;
        RECT 752.170 73.140 752.490 73.200 ;
        RECT 1805.570 73.140 1805.890 73.200 ;
      LAYER via ;
        RECT 752.200 376.080 752.460 376.340 ;
        RECT 754.960 376.080 755.220 376.340 ;
        RECT 752.200 73.140 752.460 73.400 ;
        RECT 1805.600 73.140 1805.860 73.400 ;
      LAYER met2 ;
        RECT 756.230 400.250 756.510 404.000 ;
        RECT 755.020 400.110 756.510 400.250 ;
        RECT 755.020 376.370 755.160 400.110 ;
        RECT 756.230 400.000 756.510 400.110 ;
        RECT 752.200 376.050 752.460 376.370 ;
        RECT 754.960 376.050 755.220 376.370 ;
        RECT 752.260 73.430 752.400 376.050 ;
        RECT 752.200 73.110 752.460 73.430 ;
        RECT 1805.600 73.110 1805.860 73.430 ;
        RECT 1805.660 2.400 1805.800 73.110 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.530 376.280 759.850 376.340 ;
        RECT 760.450 376.280 760.770 376.340 ;
        RECT 759.530 376.140 760.770 376.280 ;
        RECT 759.530 376.080 759.850 376.140 ;
        RECT 760.450 376.080 760.770 376.140 ;
        RECT 759.530 73.000 759.850 73.060 ;
        RECT 1823.050 73.000 1823.370 73.060 ;
        RECT 759.530 72.860 1823.370 73.000 ;
        RECT 759.530 72.800 759.850 72.860 ;
        RECT 1823.050 72.800 1823.370 72.860 ;
      LAYER via ;
        RECT 759.560 376.080 759.820 376.340 ;
        RECT 760.480 376.080 760.740 376.340 ;
        RECT 759.560 72.800 759.820 73.060 ;
        RECT 1823.080 72.800 1823.340 73.060 ;
      LAYER met2 ;
        RECT 761.750 400.250 762.030 404.000 ;
        RECT 760.540 400.110 762.030 400.250 ;
        RECT 760.540 376.370 760.680 400.110 ;
        RECT 761.750 400.000 762.030 400.110 ;
        RECT 759.560 376.050 759.820 376.370 ;
        RECT 760.480 376.050 760.740 376.370 ;
        RECT 759.620 73.090 759.760 376.050 ;
        RECT 759.560 72.770 759.820 73.090 ;
        RECT 1823.080 72.770 1823.340 73.090 ;
        RECT 1823.140 2.400 1823.280 72.770 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.890 72.660 767.210 72.720 ;
        RECT 1838.690 72.660 1839.010 72.720 ;
        RECT 766.890 72.520 1839.010 72.660 ;
        RECT 766.890 72.460 767.210 72.520 ;
        RECT 1838.690 72.460 1839.010 72.520 ;
      LAYER via ;
        RECT 766.920 72.460 767.180 72.720 ;
        RECT 1838.720 72.460 1838.980 72.720 ;
      LAYER met2 ;
        RECT 767.270 400.250 767.550 404.000 ;
        RECT 766.980 400.110 767.550 400.250 ;
        RECT 766.980 72.750 767.120 400.110 ;
        RECT 767.270 400.000 767.550 400.110 ;
        RECT 766.920 72.430 767.180 72.750 ;
        RECT 1838.720 72.430 1838.980 72.750 ;
        RECT 1838.780 1.770 1838.920 72.430 ;
        RECT 1840.870 1.770 1841.430 2.400 ;
        RECT 1838.780 1.630 1841.430 1.770 ;
        RECT 1840.870 -4.800 1841.430 1.630 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.430 375.940 766.750 376.000 ;
        RECT 771.030 375.940 771.350 376.000 ;
        RECT 766.430 375.800 771.350 375.940 ;
        RECT 766.430 375.740 766.750 375.800 ;
        RECT 771.030 375.740 771.350 375.800 ;
        RECT 766.430 72.320 766.750 72.380 ;
        RECT 1856.170 72.320 1856.490 72.380 ;
        RECT 766.430 72.180 1856.490 72.320 ;
        RECT 766.430 72.120 766.750 72.180 ;
        RECT 1856.170 72.120 1856.490 72.180 ;
      LAYER via ;
        RECT 766.460 375.740 766.720 376.000 ;
        RECT 771.060 375.740 771.320 376.000 ;
        RECT 766.460 72.120 766.720 72.380 ;
        RECT 1856.200 72.120 1856.460 72.380 ;
      LAYER met2 ;
        RECT 772.330 400.250 772.610 404.000 ;
        RECT 771.120 400.110 772.610 400.250 ;
        RECT 771.120 376.030 771.260 400.110 ;
        RECT 772.330 400.000 772.610 400.110 ;
        RECT 766.460 375.710 766.720 376.030 ;
        RECT 771.060 375.710 771.320 376.030 ;
        RECT 766.520 72.410 766.660 375.710 ;
        RECT 766.460 72.090 766.720 72.410 ;
        RECT 1856.200 72.090 1856.460 72.410 ;
        RECT 1856.260 1.770 1856.400 72.090 ;
        RECT 1858.350 1.770 1858.910 2.400 ;
        RECT 1856.260 1.630 1858.910 1.770 ;
        RECT 1858.350 -4.800 1858.910 1.630 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.330 46.140 428.650 46.200 ;
        RECT 741.590 46.140 741.910 46.200 ;
        RECT 428.330 46.000 741.910 46.140 ;
        RECT 428.330 45.940 428.650 46.000 ;
        RECT 741.590 45.940 741.910 46.000 ;
      LAYER via ;
        RECT 428.360 45.940 428.620 46.200 ;
        RECT 741.620 45.940 741.880 46.200 ;
      LAYER met2 ;
        RECT 428.250 400.180 428.530 404.000 ;
        RECT 428.250 400.000 428.560 400.180 ;
        RECT 428.420 46.230 428.560 400.000 ;
        RECT 428.360 45.910 428.620 46.230 ;
        RECT 741.620 45.910 741.880 46.230 ;
        RECT 741.680 2.400 741.820 45.910 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.330 375.940 773.650 376.000 ;
        RECT 776.550 375.940 776.870 376.000 ;
        RECT 773.330 375.800 776.870 375.940 ;
        RECT 773.330 375.740 773.650 375.800 ;
        RECT 776.550 375.740 776.870 375.800 ;
        RECT 1869.970 15.200 1870.290 15.260 ;
        RECT 1876.410 15.200 1876.730 15.260 ;
        RECT 1869.970 15.060 1876.730 15.200 ;
        RECT 1869.970 15.000 1870.290 15.060 ;
        RECT 1876.410 15.000 1876.730 15.060 ;
      LAYER via ;
        RECT 773.360 375.740 773.620 376.000 ;
        RECT 776.580 375.740 776.840 376.000 ;
        RECT 1870.000 15.000 1870.260 15.260 ;
        RECT 1876.440 15.000 1876.700 15.260 ;
      LAYER met2 ;
        RECT 777.850 400.250 778.130 404.000 ;
        RECT 776.640 400.110 778.130 400.250 ;
        RECT 776.640 376.030 776.780 400.110 ;
        RECT 777.850 400.000 778.130 400.110 ;
        RECT 773.360 375.710 773.620 376.030 ;
        RECT 776.580 375.710 776.840 376.030 ;
        RECT 773.420 72.605 773.560 375.710 ;
        RECT 773.350 72.235 773.630 72.605 ;
        RECT 1869.990 72.235 1870.270 72.605 ;
        RECT 1870.060 15.290 1870.200 72.235 ;
        RECT 1870.000 14.970 1870.260 15.290 ;
        RECT 1876.440 14.970 1876.700 15.290 ;
        RECT 1876.500 2.400 1876.640 14.970 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
      LAYER via2 ;
        RECT 773.350 72.280 773.630 72.560 ;
        RECT 1869.990 72.280 1870.270 72.560 ;
      LAYER met3 ;
        RECT 773.325 72.570 773.655 72.585 ;
        RECT 1869.965 72.570 1870.295 72.585 ;
        RECT 773.325 72.270 1870.295 72.570 ;
        RECT 773.325 72.255 773.655 72.270 ;
        RECT 1869.965 72.255 1870.295 72.270 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.230 120.260 780.550 120.320 ;
        RECT 1890.670 120.260 1890.990 120.320 ;
        RECT 780.230 120.120 1890.990 120.260 ;
        RECT 780.230 120.060 780.550 120.120 ;
        RECT 1890.670 120.060 1890.990 120.120 ;
      LAYER via ;
        RECT 780.260 120.060 780.520 120.320 ;
        RECT 1890.700 120.060 1890.960 120.320 ;
      LAYER met2 ;
        RECT 783.370 400.250 783.650 404.000 ;
        RECT 782.160 400.110 783.650 400.250 ;
        RECT 782.160 351.970 782.300 400.110 ;
        RECT 783.370 400.000 783.650 400.110 ;
        RECT 780.320 351.830 782.300 351.970 ;
        RECT 780.320 120.350 780.460 351.830 ;
        RECT 780.260 120.030 780.520 120.350 ;
        RECT 1890.700 120.030 1890.960 120.350 ;
        RECT 1890.760 82.870 1890.900 120.030 ;
        RECT 1890.760 82.730 1892.280 82.870 ;
        RECT 1892.140 1.770 1892.280 82.730 ;
        RECT 1894.230 1.770 1894.790 2.400 ;
        RECT 1892.140 1.630 1894.790 1.770 ;
        RECT 1894.230 -4.800 1894.790 1.630 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.590 124.000 787.910 124.060 ;
        RECT 1911.830 124.000 1912.150 124.060 ;
        RECT 787.590 123.860 1912.150 124.000 ;
        RECT 787.590 123.800 787.910 123.860 ;
        RECT 1911.830 123.800 1912.150 123.860 ;
      LAYER via ;
        RECT 787.620 123.800 787.880 124.060 ;
        RECT 1911.860 123.800 1912.120 124.060 ;
      LAYER met2 ;
        RECT 788.890 400.250 789.170 404.000 ;
        RECT 787.680 400.110 789.170 400.250 ;
        RECT 787.680 124.090 787.820 400.110 ;
        RECT 788.890 400.000 789.170 400.110 ;
        RECT 787.620 123.770 787.880 124.090 ;
        RECT 1911.860 123.770 1912.120 124.090 ;
        RECT 1911.920 2.400 1912.060 123.770 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.490 123.660 794.810 123.720 ;
        RECT 1925.170 123.660 1925.490 123.720 ;
        RECT 794.490 123.520 1925.490 123.660 ;
        RECT 794.490 123.460 794.810 123.520 ;
        RECT 1925.170 123.460 1925.490 123.520 ;
      LAYER via ;
        RECT 794.520 123.460 794.780 123.720 ;
        RECT 1925.200 123.460 1925.460 123.720 ;
      LAYER met2 ;
        RECT 794.410 400.180 794.690 404.000 ;
        RECT 794.410 400.000 794.720 400.180 ;
        RECT 794.580 123.750 794.720 400.000 ;
        RECT 794.520 123.430 794.780 123.750 ;
        RECT 1925.200 123.430 1925.460 123.750 ;
        RECT 1925.260 82.870 1925.400 123.430 ;
        RECT 1925.260 82.730 1930.000 82.870 ;
        RECT 1929.860 2.400 1930.000 82.730 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.030 375.940 794.350 376.000 ;
        RECT 798.630 375.940 798.950 376.000 ;
        RECT 794.030 375.800 798.950 375.940 ;
        RECT 794.030 375.740 794.350 375.800 ;
        RECT 798.630 375.740 798.950 375.800 ;
        RECT 794.030 123.320 794.350 123.380 ;
        RECT 1945.870 123.320 1946.190 123.380 ;
        RECT 794.030 123.180 1946.190 123.320 ;
        RECT 794.030 123.120 794.350 123.180 ;
        RECT 1945.870 123.120 1946.190 123.180 ;
      LAYER via ;
        RECT 794.060 375.740 794.320 376.000 ;
        RECT 798.660 375.740 798.920 376.000 ;
        RECT 794.060 123.120 794.320 123.380 ;
        RECT 1945.900 123.120 1946.160 123.380 ;
      LAYER met2 ;
        RECT 799.930 400.250 800.210 404.000 ;
        RECT 798.720 400.110 800.210 400.250 ;
        RECT 798.720 376.030 798.860 400.110 ;
        RECT 799.930 400.000 800.210 400.110 ;
        RECT 794.060 375.710 794.320 376.030 ;
        RECT 798.660 375.710 798.920 376.030 ;
        RECT 794.120 123.410 794.260 375.710 ;
        RECT 794.060 123.090 794.320 123.410 ;
        RECT 1945.900 123.090 1946.160 123.410 ;
        RECT 1945.960 82.870 1946.100 123.090 ;
        RECT 1945.960 82.730 1947.480 82.870 ;
        RECT 1947.340 2.400 1947.480 82.730 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.930 122.980 801.250 123.040 ;
        RECT 1959.670 122.980 1959.990 123.040 ;
        RECT 800.930 122.840 1959.990 122.980 ;
        RECT 800.930 122.780 801.250 122.840 ;
        RECT 1959.670 122.780 1959.990 122.840 ;
      LAYER via ;
        RECT 800.960 122.780 801.220 123.040 ;
        RECT 1959.700 122.780 1959.960 123.040 ;
      LAYER met2 ;
        RECT 805.450 400.250 805.730 404.000 ;
        RECT 804.240 400.110 805.730 400.250 ;
        RECT 804.240 324.370 804.380 400.110 ;
        RECT 805.450 400.000 805.730 400.110 ;
        RECT 801.020 324.230 804.380 324.370 ;
        RECT 801.020 123.070 801.160 324.230 ;
        RECT 800.960 122.750 801.220 123.070 ;
        RECT 1959.700 122.750 1959.960 123.070 ;
        RECT 1959.760 82.870 1959.900 122.750 ;
        RECT 1959.760 82.730 1963.120 82.870 ;
        RECT 1962.980 1.770 1963.120 82.730 ;
        RECT 1965.070 1.770 1965.630 2.400 ;
        RECT 1962.980 1.630 1965.630 1.770 ;
        RECT 1965.070 -4.800 1965.630 1.630 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.830 376.280 808.150 376.340 ;
        RECT 809.670 376.280 809.990 376.340 ;
        RECT 807.830 376.140 809.990 376.280 ;
        RECT 807.830 376.080 808.150 376.140 ;
        RECT 809.670 376.080 809.990 376.140 ;
        RECT 807.830 78.100 808.150 78.160 ;
        RECT 1980.370 78.100 1980.690 78.160 ;
        RECT 807.830 77.960 1980.690 78.100 ;
        RECT 807.830 77.900 808.150 77.960 ;
        RECT 1980.370 77.900 1980.690 77.960 ;
      LAYER via ;
        RECT 807.860 376.080 808.120 376.340 ;
        RECT 809.700 376.080 809.960 376.340 ;
        RECT 807.860 77.900 808.120 78.160 ;
        RECT 1980.400 77.900 1980.660 78.160 ;
      LAYER met2 ;
        RECT 810.970 400.250 811.250 404.000 ;
        RECT 809.760 400.110 811.250 400.250 ;
        RECT 809.760 376.370 809.900 400.110 ;
        RECT 810.970 400.000 811.250 400.110 ;
        RECT 807.860 376.050 808.120 376.370 ;
        RECT 809.700 376.050 809.960 376.370 ;
        RECT 807.920 78.190 808.060 376.050 ;
        RECT 807.860 77.870 808.120 78.190 ;
        RECT 1980.400 77.870 1980.660 78.190 ;
        RECT 1980.460 1.770 1980.600 77.870 ;
        RECT 1982.550 1.770 1983.110 2.400 ;
        RECT 1980.460 1.630 1983.110 1.770 ;
        RECT 1982.550 -4.800 1983.110 1.630 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 815.190 78.440 815.510 78.500 ;
        RECT 1994.170 78.440 1994.490 78.500 ;
        RECT 815.190 78.300 1994.490 78.440 ;
        RECT 815.190 78.240 815.510 78.300 ;
        RECT 1994.170 78.240 1994.490 78.300 ;
        RECT 1994.170 15.200 1994.490 15.260 ;
        RECT 2000.610 15.200 2000.930 15.260 ;
        RECT 1994.170 15.060 2000.930 15.200 ;
        RECT 1994.170 15.000 1994.490 15.060 ;
        RECT 2000.610 15.000 2000.930 15.060 ;
      LAYER via ;
        RECT 815.220 78.240 815.480 78.500 ;
        RECT 1994.200 78.240 1994.460 78.500 ;
        RECT 1994.200 15.000 1994.460 15.260 ;
        RECT 2000.640 15.000 2000.900 15.260 ;
      LAYER met2 ;
        RECT 816.490 400.250 816.770 404.000 ;
        RECT 815.280 400.110 816.770 400.250 ;
        RECT 815.280 78.530 815.420 400.110 ;
        RECT 816.490 400.000 816.770 400.110 ;
        RECT 815.220 78.210 815.480 78.530 ;
        RECT 1994.200 78.210 1994.460 78.530 ;
        RECT 1994.260 15.290 1994.400 78.210 ;
        RECT 1994.200 14.970 1994.460 15.290 ;
        RECT 2000.640 14.970 2000.900 15.290 ;
        RECT 2000.700 2.400 2000.840 14.970 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.630 78.780 821.950 78.840 ;
        RECT 2018.090 78.780 2018.410 78.840 ;
        RECT 821.630 78.640 2018.410 78.780 ;
        RECT 821.630 78.580 821.950 78.640 ;
        RECT 2018.090 78.580 2018.410 78.640 ;
      LAYER via ;
        RECT 821.660 78.580 821.920 78.840 ;
        RECT 2018.120 78.580 2018.380 78.840 ;
      LAYER met2 ;
        RECT 821.550 400.180 821.830 404.000 ;
        RECT 821.550 400.000 821.860 400.180 ;
        RECT 821.720 78.870 821.860 400.000 ;
        RECT 821.660 78.550 821.920 78.870 ;
        RECT 2018.120 78.550 2018.380 78.870 ;
        RECT 2018.180 2.400 2018.320 78.550 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 822.090 79.120 822.410 79.180 ;
        RECT 2036.030 79.120 2036.350 79.180 ;
        RECT 822.090 78.980 2036.350 79.120 ;
        RECT 822.090 78.920 822.410 78.980 ;
        RECT 2036.030 78.920 2036.350 78.980 ;
      LAYER via ;
        RECT 822.120 78.920 822.380 79.180 ;
        RECT 2036.060 78.920 2036.320 79.180 ;
      LAYER met2 ;
        RECT 827.070 400.250 827.350 404.000 ;
        RECT 825.860 400.110 827.350 400.250 ;
        RECT 825.860 324.370 826.000 400.110 ;
        RECT 827.070 400.000 827.350 400.110 ;
        RECT 822.180 324.230 826.000 324.370 ;
        RECT 822.180 79.210 822.320 324.230 ;
        RECT 822.120 78.890 822.380 79.210 ;
        RECT 2036.060 78.890 2036.320 79.210 ;
        RECT 2036.120 2.400 2036.260 78.890 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.790 45.800 429.110 45.860 ;
        RECT 759.070 45.800 759.390 45.860 ;
        RECT 428.790 45.660 759.390 45.800 ;
        RECT 428.790 45.600 429.110 45.660 ;
        RECT 759.070 45.600 759.390 45.660 ;
      LAYER via ;
        RECT 428.820 45.600 429.080 45.860 ;
        RECT 759.100 45.600 759.360 45.860 ;
      LAYER met2 ;
        RECT 433.770 400.250 434.050 404.000 ;
        RECT 432.560 400.110 434.050 400.250 ;
        RECT 432.560 324.370 432.700 400.110 ;
        RECT 433.770 400.000 434.050 400.110 ;
        RECT 428.880 324.230 432.700 324.370 ;
        RECT 428.880 45.890 429.020 324.230 ;
        RECT 428.820 45.570 429.080 45.890 ;
        RECT 759.100 45.570 759.360 45.890 ;
        RECT 759.160 2.400 759.300 45.570 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.530 375.940 828.850 376.000 ;
        RECT 831.290 375.940 831.610 376.000 ;
        RECT 828.530 375.800 831.610 375.940 ;
        RECT 828.530 375.740 828.850 375.800 ;
        RECT 831.290 375.740 831.610 375.800 ;
        RECT 828.530 82.860 828.850 82.920 ;
        RECT 2053.970 82.860 2054.290 82.920 ;
        RECT 828.530 82.720 2054.290 82.860 ;
        RECT 828.530 82.660 828.850 82.720 ;
        RECT 2053.970 82.660 2054.290 82.720 ;
      LAYER via ;
        RECT 828.560 375.740 828.820 376.000 ;
        RECT 831.320 375.740 831.580 376.000 ;
        RECT 828.560 82.660 828.820 82.920 ;
        RECT 2054.000 82.660 2054.260 82.920 ;
      LAYER met2 ;
        RECT 832.590 400.250 832.870 404.000 ;
        RECT 831.380 400.110 832.870 400.250 ;
        RECT 831.380 376.030 831.520 400.110 ;
        RECT 832.590 400.000 832.870 400.110 ;
        RECT 828.560 375.710 828.820 376.030 ;
        RECT 831.320 375.710 831.580 376.030 ;
        RECT 828.620 82.950 828.760 375.710 ;
        RECT 828.560 82.630 828.820 82.950 ;
        RECT 2054.000 82.630 2054.260 82.950 ;
        RECT 2054.060 2.400 2054.200 82.630 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.430 82.520 835.750 82.580 ;
        RECT 2071.450 82.520 2071.770 82.580 ;
        RECT 835.430 82.380 2071.770 82.520 ;
        RECT 835.430 82.320 835.750 82.380 ;
        RECT 2071.450 82.320 2071.770 82.380 ;
      LAYER via ;
        RECT 835.460 82.320 835.720 82.580 ;
        RECT 2071.480 82.320 2071.740 82.580 ;
      LAYER met2 ;
        RECT 838.110 400.250 838.390 404.000 ;
        RECT 836.900 400.110 838.390 400.250 ;
        RECT 836.900 386.480 837.040 400.110 ;
        RECT 838.110 400.000 838.390 400.110 ;
        RECT 835.520 386.340 837.040 386.480 ;
        RECT 835.520 82.610 835.660 386.340 ;
        RECT 835.460 82.290 835.720 82.610 ;
        RECT 2071.480 82.290 2071.740 82.610 ;
        RECT 2071.540 2.400 2071.680 82.290 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.790 82.180 843.110 82.240 ;
        RECT 2087.090 82.180 2087.410 82.240 ;
        RECT 842.790 82.040 2087.410 82.180 ;
        RECT 842.790 81.980 843.110 82.040 ;
        RECT 2087.090 81.980 2087.410 82.040 ;
      LAYER via ;
        RECT 842.820 81.980 843.080 82.240 ;
        RECT 2087.120 81.980 2087.380 82.240 ;
      LAYER met2 ;
        RECT 843.630 400.250 843.910 404.000 ;
        RECT 842.880 400.110 843.910 400.250 ;
        RECT 842.880 82.270 843.020 400.110 ;
        RECT 843.630 400.000 843.910 400.110 ;
        RECT 842.820 81.950 843.080 82.270 ;
        RECT 2087.120 81.950 2087.380 82.270 ;
        RECT 2087.180 1.770 2087.320 81.950 ;
        RECT 2089.270 1.770 2089.830 2.400 ;
        RECT 2087.180 1.630 2089.830 1.770 ;
        RECT 2089.270 -4.800 2089.830 1.630 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 849.230 81.840 849.550 81.900 ;
        RECT 2104.570 81.840 2104.890 81.900 ;
        RECT 849.230 81.700 2104.890 81.840 ;
        RECT 849.230 81.640 849.550 81.700 ;
        RECT 2104.570 81.640 2104.890 81.700 ;
      LAYER via ;
        RECT 849.260 81.640 849.520 81.900 ;
        RECT 2104.600 81.640 2104.860 81.900 ;
      LAYER met2 ;
        RECT 849.150 400.180 849.430 404.000 ;
        RECT 849.150 400.000 849.460 400.180 ;
        RECT 849.320 81.930 849.460 400.000 ;
        RECT 849.260 81.610 849.520 81.930 ;
        RECT 2104.600 81.610 2104.860 81.930 ;
        RECT 2104.660 1.770 2104.800 81.610 ;
        RECT 2106.750 1.770 2107.310 2.400 ;
        RECT 2104.660 1.630 2107.310 1.770 ;
        RECT 2106.750 -4.800 2107.310 1.630 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 849.690 386.480 850.010 386.540 ;
        RECT 853.370 386.480 853.690 386.540 ;
        RECT 849.690 386.340 853.690 386.480 ;
        RECT 849.690 386.280 850.010 386.340 ;
        RECT 853.370 386.280 853.690 386.340 ;
        RECT 849.690 81.500 850.010 81.560 ;
        RECT 2118.370 81.500 2118.690 81.560 ;
        RECT 849.690 81.360 2118.690 81.500 ;
        RECT 849.690 81.300 850.010 81.360 ;
        RECT 2118.370 81.300 2118.690 81.360 ;
        RECT 2118.370 15.880 2118.690 15.940 ;
        RECT 2124.810 15.880 2125.130 15.940 ;
        RECT 2118.370 15.740 2125.130 15.880 ;
        RECT 2118.370 15.680 2118.690 15.740 ;
        RECT 2124.810 15.680 2125.130 15.740 ;
      LAYER via ;
        RECT 849.720 386.280 849.980 386.540 ;
        RECT 853.400 386.280 853.660 386.540 ;
        RECT 849.720 81.300 849.980 81.560 ;
        RECT 2118.400 81.300 2118.660 81.560 ;
        RECT 2118.400 15.680 2118.660 15.940 ;
        RECT 2124.840 15.680 2125.100 15.940 ;
      LAYER met2 ;
        RECT 854.670 400.250 854.950 404.000 ;
        RECT 853.460 400.110 854.950 400.250 ;
        RECT 853.460 386.570 853.600 400.110 ;
        RECT 854.670 400.000 854.950 400.110 ;
        RECT 849.720 386.250 849.980 386.570 ;
        RECT 853.400 386.250 853.660 386.570 ;
        RECT 849.780 81.590 849.920 386.250 ;
        RECT 849.720 81.270 849.980 81.590 ;
        RECT 2118.400 81.270 2118.660 81.590 ;
        RECT 2118.460 15.970 2118.600 81.270 ;
        RECT 2118.400 15.650 2118.660 15.970 ;
        RECT 2124.840 15.650 2125.100 15.970 ;
        RECT 2124.900 2.400 2125.040 15.650 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.590 386.480 856.910 386.540 ;
        RECT 858.890 386.480 859.210 386.540 ;
        RECT 856.590 386.340 859.210 386.480 ;
        RECT 856.590 386.280 856.910 386.340 ;
        RECT 858.890 386.280 859.210 386.340 ;
        RECT 856.590 81.160 856.910 81.220 ;
        RECT 2142.290 81.160 2142.610 81.220 ;
        RECT 856.590 81.020 2142.610 81.160 ;
        RECT 856.590 80.960 856.910 81.020 ;
        RECT 2142.290 80.960 2142.610 81.020 ;
      LAYER via ;
        RECT 856.620 386.280 856.880 386.540 ;
        RECT 858.920 386.280 859.180 386.540 ;
        RECT 856.620 80.960 856.880 81.220 ;
        RECT 2142.320 80.960 2142.580 81.220 ;
      LAYER met2 ;
        RECT 860.190 400.250 860.470 404.000 ;
        RECT 858.980 400.110 860.470 400.250 ;
        RECT 858.980 386.570 859.120 400.110 ;
        RECT 860.190 400.000 860.470 400.110 ;
        RECT 856.620 386.250 856.880 386.570 ;
        RECT 858.920 386.250 859.180 386.570 ;
        RECT 856.680 81.250 856.820 386.250 ;
        RECT 856.620 80.930 856.880 81.250 ;
        RECT 2142.320 80.930 2142.580 81.250 ;
        RECT 2142.380 2.400 2142.520 80.930 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.030 386.480 863.350 386.540 ;
        RECT 864.410 386.480 864.730 386.540 ;
        RECT 863.030 386.340 864.730 386.480 ;
        RECT 863.030 386.280 863.350 386.340 ;
        RECT 864.410 386.280 864.730 386.340 ;
        RECT 863.030 80.820 863.350 80.880 ;
        RECT 2160.230 80.820 2160.550 80.880 ;
        RECT 863.030 80.680 2160.550 80.820 ;
        RECT 863.030 80.620 863.350 80.680 ;
        RECT 2160.230 80.620 2160.550 80.680 ;
      LAYER via ;
        RECT 863.060 386.280 863.320 386.540 ;
        RECT 864.440 386.280 864.700 386.540 ;
        RECT 863.060 80.620 863.320 80.880 ;
        RECT 2160.260 80.620 2160.520 80.880 ;
      LAYER met2 ;
        RECT 865.250 400.250 865.530 404.000 ;
        RECT 864.500 400.110 865.530 400.250 ;
        RECT 864.500 386.570 864.640 400.110 ;
        RECT 865.250 400.000 865.530 400.110 ;
        RECT 863.060 386.250 863.320 386.570 ;
        RECT 864.440 386.250 864.700 386.570 ;
        RECT 863.120 80.910 863.260 386.250 ;
        RECT 863.060 80.590 863.320 80.910 ;
        RECT 2160.260 80.590 2160.520 80.910 ;
        RECT 2160.320 2.400 2160.460 80.590 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.930 80.480 870.250 80.540 ;
        RECT 2175.410 80.480 2175.730 80.540 ;
        RECT 869.930 80.340 2175.730 80.480 ;
        RECT 869.930 80.280 870.250 80.340 ;
        RECT 2175.410 80.280 2175.730 80.340 ;
      LAYER via ;
        RECT 869.960 80.280 870.220 80.540 ;
        RECT 2175.440 80.280 2175.700 80.540 ;
      LAYER met2 ;
        RECT 870.770 400.250 871.050 404.000 ;
        RECT 870.020 400.110 871.050 400.250 ;
        RECT 870.020 80.570 870.160 400.110 ;
        RECT 870.770 400.000 871.050 400.110 ;
        RECT 869.960 80.250 870.220 80.570 ;
        RECT 2175.440 80.250 2175.700 80.570 ;
        RECT 2175.500 1.770 2175.640 80.250 ;
        RECT 2177.590 1.770 2178.150 2.400 ;
        RECT 2175.500 1.630 2178.150 1.770 ;
        RECT 2177.590 -4.800 2178.150 1.630 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 877.290 80.140 877.610 80.200 ;
        RECT 2195.650 80.140 2195.970 80.200 ;
        RECT 877.290 80.000 2195.970 80.140 ;
        RECT 877.290 79.940 877.610 80.000 ;
        RECT 2195.650 79.940 2195.970 80.000 ;
      LAYER via ;
        RECT 877.320 79.940 877.580 80.200 ;
        RECT 2195.680 79.940 2195.940 80.200 ;
      LAYER met2 ;
        RECT 876.290 400.250 876.570 404.000 ;
        RECT 876.290 400.110 877.520 400.250 ;
        RECT 876.290 400.000 876.570 400.110 ;
        RECT 877.380 80.230 877.520 400.110 ;
        RECT 877.320 79.910 877.580 80.230 ;
        RECT 2195.680 79.910 2195.940 80.230 ;
        RECT 2195.740 2.400 2195.880 79.910 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.830 386.140 877.150 386.200 ;
        RECT 880.510 386.140 880.830 386.200 ;
        RECT 876.830 386.000 880.830 386.140 ;
        RECT 876.830 385.940 877.150 386.000 ;
        RECT 880.510 385.940 880.830 386.000 ;
        RECT 876.830 79.800 877.150 79.860 ;
        RECT 2213.130 79.800 2213.450 79.860 ;
        RECT 876.830 79.660 2213.450 79.800 ;
        RECT 876.830 79.600 877.150 79.660 ;
        RECT 2213.130 79.600 2213.450 79.660 ;
      LAYER via ;
        RECT 876.860 385.940 877.120 386.200 ;
        RECT 880.540 385.940 880.800 386.200 ;
        RECT 876.860 79.600 877.120 79.860 ;
        RECT 2213.160 79.600 2213.420 79.860 ;
      LAYER met2 ;
        RECT 881.810 400.250 882.090 404.000 ;
        RECT 880.600 400.110 882.090 400.250 ;
        RECT 880.600 386.230 880.740 400.110 ;
        RECT 881.810 400.000 882.090 400.110 ;
        RECT 876.860 385.910 877.120 386.230 ;
        RECT 880.540 385.910 880.800 386.230 ;
        RECT 876.920 79.890 877.060 385.910 ;
        RECT 876.860 79.570 877.120 79.890 ;
        RECT 2213.160 79.570 2213.420 79.890 ;
        RECT 2213.220 2.400 2213.360 79.570 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 436.150 45.460 436.470 45.520 ;
        RECT 777.010 45.460 777.330 45.520 ;
        RECT 436.150 45.320 777.330 45.460 ;
        RECT 436.150 45.260 436.470 45.320 ;
        RECT 777.010 45.260 777.330 45.320 ;
      LAYER via ;
        RECT 436.180 45.260 436.440 45.520 ;
        RECT 777.040 45.260 777.300 45.520 ;
      LAYER met2 ;
        RECT 438.830 400.250 439.110 404.000 ;
        RECT 438.080 400.110 439.110 400.250 ;
        RECT 438.080 324.370 438.220 400.110 ;
        RECT 438.830 400.000 439.110 400.110 ;
        RECT 436.240 324.230 438.220 324.370 ;
        RECT 436.240 45.550 436.380 324.230 ;
        RECT 436.180 45.230 436.440 45.550 ;
        RECT 777.040 45.230 777.300 45.550 ;
        RECT 777.100 2.400 777.240 45.230 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 884.650 79.460 884.970 79.520 ;
        RECT 2228.770 79.460 2229.090 79.520 ;
        RECT 884.650 79.320 2229.090 79.460 ;
        RECT 884.650 79.260 884.970 79.320 ;
        RECT 2228.770 79.260 2229.090 79.320 ;
      LAYER via ;
        RECT 884.680 79.260 884.940 79.520 ;
        RECT 2228.800 79.260 2229.060 79.520 ;
      LAYER met2 ;
        RECT 887.330 400.250 887.610 404.000 ;
        RECT 886.120 400.110 887.610 400.250 ;
        RECT 886.120 324.370 886.260 400.110 ;
        RECT 887.330 400.000 887.610 400.110 ;
        RECT 884.740 324.230 886.260 324.370 ;
        RECT 884.740 79.550 884.880 324.230 ;
        RECT 884.680 79.230 884.940 79.550 ;
        RECT 2228.800 79.230 2229.060 79.550 ;
        RECT 2228.860 1.770 2229.000 79.230 ;
        RECT 2230.950 1.770 2231.510 2.400 ;
        RECT 2228.860 1.630 2231.510 1.770 ;
        RECT 2230.950 -4.800 2231.510 1.630 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2242.570 16.900 2242.890 16.960 ;
        RECT 2249.010 16.900 2249.330 16.960 ;
        RECT 2242.570 16.760 2249.330 16.900 ;
        RECT 2242.570 16.700 2242.890 16.760 ;
        RECT 2249.010 16.700 2249.330 16.760 ;
      LAYER via ;
        RECT 2242.600 16.700 2242.860 16.960 ;
        RECT 2249.040 16.700 2249.300 16.960 ;
      LAYER met2 ;
        RECT 892.850 400.250 893.130 404.000 ;
        RECT 891.640 400.110 893.130 400.250 ;
        RECT 891.640 80.085 891.780 400.110 ;
        RECT 892.850 400.000 893.130 400.110 ;
        RECT 891.570 79.715 891.850 80.085 ;
        RECT 2242.590 79.715 2242.870 80.085 ;
        RECT 2242.660 16.990 2242.800 79.715 ;
        RECT 2242.600 16.670 2242.860 16.990 ;
        RECT 2249.040 16.670 2249.300 16.990 ;
        RECT 2249.100 2.400 2249.240 16.670 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
      LAYER via2 ;
        RECT 891.570 79.760 891.850 80.040 ;
        RECT 2242.590 79.760 2242.870 80.040 ;
      LAYER met3 ;
        RECT 891.545 80.050 891.875 80.065 ;
        RECT 2242.565 80.050 2242.895 80.065 ;
        RECT 891.545 79.750 2242.895 80.050 ;
        RECT 891.545 79.735 891.875 79.750 ;
        RECT 2242.565 79.735 2242.895 79.750 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.370 400.180 898.650 404.000 ;
        RECT 898.370 400.000 898.680 400.180 ;
        RECT 898.540 324.370 898.680 400.000 ;
        RECT 898.080 324.230 898.680 324.370 ;
        RECT 898.080 79.405 898.220 324.230 ;
        RECT 898.010 79.035 898.290 79.405 ;
        RECT 2266.510 79.035 2266.790 79.405 ;
        RECT 2266.580 2.400 2266.720 79.035 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
      LAYER via2 ;
        RECT 898.010 79.080 898.290 79.360 ;
        RECT 2266.510 79.080 2266.790 79.360 ;
      LAYER met3 ;
        RECT 897.985 79.370 898.315 79.385 ;
        RECT 2266.485 79.370 2266.815 79.385 ;
        RECT 897.985 79.070 2266.815 79.370 ;
        RECT 897.985 79.055 898.315 79.070 ;
        RECT 2266.485 79.055 2266.815 79.070 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.890 122.640 905.210 122.700 ;
        RECT 2284.430 122.640 2284.750 122.700 ;
        RECT 904.890 122.500 2284.750 122.640 ;
        RECT 904.890 122.440 905.210 122.500 ;
        RECT 2284.430 122.440 2284.750 122.500 ;
      LAYER via ;
        RECT 904.920 122.440 905.180 122.700 ;
        RECT 2284.460 122.440 2284.720 122.700 ;
      LAYER met2 ;
        RECT 903.890 400.250 904.170 404.000 ;
        RECT 903.890 400.110 905.120 400.250 ;
        RECT 903.890 400.000 904.170 400.110 ;
        RECT 904.980 122.730 905.120 400.110 ;
        RECT 904.920 122.410 905.180 122.730 ;
        RECT 2284.460 122.410 2284.720 122.730 ;
        RECT 2284.520 2.400 2284.660 122.410 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 905.350 122.300 905.670 122.360 ;
        RECT 2297.770 122.300 2298.090 122.360 ;
        RECT 905.350 122.160 2298.090 122.300 ;
        RECT 905.350 122.100 905.670 122.160 ;
        RECT 2297.770 122.100 2298.090 122.160 ;
      LAYER via ;
        RECT 905.380 122.100 905.640 122.360 ;
        RECT 2297.800 122.100 2298.060 122.360 ;
      LAYER met2 ;
        RECT 909.410 400.250 909.690 404.000 ;
        RECT 908.200 400.110 909.690 400.250 ;
        RECT 908.200 324.370 908.340 400.110 ;
        RECT 909.410 400.000 909.690 400.110 ;
        RECT 905.440 324.230 908.340 324.370 ;
        RECT 905.440 122.390 905.580 324.230 ;
        RECT 905.380 122.070 905.640 122.390 ;
        RECT 2297.800 122.070 2298.060 122.390 ;
        RECT 2297.860 82.870 2298.000 122.070 ;
        RECT 2297.860 82.730 2299.840 82.870 ;
        RECT 2299.700 1.770 2299.840 82.730 ;
        RECT 2301.790 1.770 2302.350 2.400 ;
        RECT 2299.700 1.630 2302.350 1.770 ;
        RECT 2301.790 -4.800 2302.350 1.630 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 912.250 121.960 912.570 122.020 ;
        RECT 2318.470 121.960 2318.790 122.020 ;
        RECT 912.250 121.820 2318.790 121.960 ;
        RECT 912.250 121.760 912.570 121.820 ;
        RECT 2318.470 121.760 2318.790 121.820 ;
      LAYER via ;
        RECT 912.280 121.760 912.540 122.020 ;
        RECT 2318.500 121.760 2318.760 122.020 ;
      LAYER met2 ;
        RECT 914.470 400.250 914.750 404.000 ;
        RECT 913.260 400.110 914.750 400.250 ;
        RECT 913.260 324.370 913.400 400.110 ;
        RECT 914.470 400.000 914.750 400.110 ;
        RECT 912.340 324.230 913.400 324.370 ;
        RECT 912.340 122.050 912.480 324.230 ;
        RECT 912.280 121.730 912.540 122.050 ;
        RECT 2318.500 121.730 2318.760 122.050 ;
        RECT 2318.560 82.870 2318.700 121.730 ;
        RECT 2318.560 82.730 2320.080 82.870 ;
        RECT 2319.940 2.400 2320.080 82.730 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 919.150 121.620 919.470 121.680 ;
        RECT 2332.270 121.620 2332.590 121.680 ;
        RECT 919.150 121.480 2332.590 121.620 ;
        RECT 919.150 121.420 919.470 121.480 ;
        RECT 2332.270 121.420 2332.590 121.480 ;
      LAYER via ;
        RECT 919.180 121.420 919.440 121.680 ;
        RECT 2332.300 121.420 2332.560 121.680 ;
      LAYER met2 ;
        RECT 919.990 400.250 920.270 404.000 ;
        RECT 919.240 400.110 920.270 400.250 ;
        RECT 919.240 121.710 919.380 400.110 ;
        RECT 919.990 400.000 920.270 400.110 ;
        RECT 919.180 121.390 919.440 121.710 ;
        RECT 2332.300 121.390 2332.560 121.710 ;
        RECT 2332.360 82.870 2332.500 121.390 ;
        RECT 2332.360 82.730 2337.560 82.870 ;
        RECT 2337.420 2.400 2337.560 82.730 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 926.050 121.280 926.370 121.340 ;
        RECT 2352.970 121.280 2353.290 121.340 ;
        RECT 926.050 121.140 2353.290 121.280 ;
        RECT 926.050 121.080 926.370 121.140 ;
        RECT 2352.970 121.080 2353.290 121.140 ;
      LAYER via ;
        RECT 926.080 121.080 926.340 121.340 ;
        RECT 2353.000 121.080 2353.260 121.340 ;
      LAYER met2 ;
        RECT 925.510 400.250 925.790 404.000 ;
        RECT 925.510 400.110 926.280 400.250 ;
        RECT 925.510 400.000 925.790 400.110 ;
        RECT 926.140 121.370 926.280 400.110 ;
        RECT 926.080 121.050 926.340 121.370 ;
        RECT 2353.000 121.050 2353.260 121.370 ;
        RECT 2353.060 1.770 2353.200 121.050 ;
        RECT 2355.150 1.770 2355.710 2.400 ;
        RECT 2353.060 1.630 2355.710 1.770 ;
        RECT 2355.150 -4.800 2355.710 1.630 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.590 386.820 925.910 386.880 ;
        RECT 929.730 386.820 930.050 386.880 ;
        RECT 925.590 386.680 930.050 386.820 ;
        RECT 925.590 386.620 925.910 386.680 ;
        RECT 929.730 386.620 930.050 386.680 ;
        RECT 925.590 84.900 925.910 84.960 ;
        RECT 2366.770 84.900 2367.090 84.960 ;
        RECT 925.590 84.760 2367.090 84.900 ;
        RECT 925.590 84.700 925.910 84.760 ;
        RECT 2366.770 84.700 2367.090 84.760 ;
        RECT 2366.770 17.580 2367.090 17.640 ;
        RECT 2370.910 17.580 2371.230 17.640 ;
        RECT 2366.770 17.440 2371.230 17.580 ;
        RECT 2366.770 17.380 2367.090 17.440 ;
        RECT 2370.910 17.380 2371.230 17.440 ;
      LAYER via ;
        RECT 925.620 386.620 925.880 386.880 ;
        RECT 929.760 386.620 930.020 386.880 ;
        RECT 925.620 84.700 925.880 84.960 ;
        RECT 2366.800 84.700 2367.060 84.960 ;
        RECT 2366.800 17.380 2367.060 17.640 ;
        RECT 2370.940 17.380 2371.200 17.640 ;
      LAYER met2 ;
        RECT 931.030 400.250 931.310 404.000 ;
        RECT 929.820 400.110 931.310 400.250 ;
        RECT 929.820 386.910 929.960 400.110 ;
        RECT 931.030 400.000 931.310 400.110 ;
        RECT 925.620 386.590 925.880 386.910 ;
        RECT 929.760 386.590 930.020 386.910 ;
        RECT 925.680 84.990 925.820 386.590 ;
        RECT 925.620 84.670 925.880 84.990 ;
        RECT 2366.800 84.670 2367.060 84.990 ;
        RECT 2366.860 17.670 2367.000 84.670 ;
        RECT 2366.800 17.350 2367.060 17.670 ;
        RECT 2370.940 17.350 2371.200 17.670 ;
        RECT 2371.000 1.770 2371.140 17.350 ;
        RECT 2372.630 1.770 2373.190 2.400 ;
        RECT 2371.000 1.630 2373.190 1.770 ;
        RECT 2372.630 -4.800 2373.190 1.630 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.490 85.240 932.810 85.300 ;
        RECT 2387.470 85.240 2387.790 85.300 ;
        RECT 932.490 85.100 2387.790 85.240 ;
        RECT 932.490 85.040 932.810 85.100 ;
        RECT 2387.470 85.040 2387.790 85.100 ;
      LAYER via ;
        RECT 932.520 85.040 932.780 85.300 ;
        RECT 2387.500 85.040 2387.760 85.300 ;
      LAYER met2 ;
        RECT 936.550 400.250 936.830 404.000 ;
        RECT 935.340 400.110 936.830 400.250 ;
        RECT 935.340 324.370 935.480 400.110 ;
        RECT 936.550 400.000 936.830 400.110 ;
        RECT 932.580 324.230 935.480 324.370 ;
        RECT 932.580 85.330 932.720 324.230 ;
        RECT 932.520 85.010 932.780 85.330 ;
        RECT 2387.500 85.010 2387.760 85.330 ;
        RECT 2387.560 82.870 2387.700 85.010 ;
        RECT 2387.560 82.730 2390.920 82.870 ;
        RECT 2390.780 2.400 2390.920 82.730 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.590 45.120 442.910 45.180 ;
        RECT 794.490 45.120 794.810 45.180 ;
        RECT 442.590 44.980 794.810 45.120 ;
        RECT 442.590 44.920 442.910 44.980 ;
        RECT 794.490 44.920 794.810 44.980 ;
      LAYER via ;
        RECT 442.620 44.920 442.880 45.180 ;
        RECT 794.520 44.920 794.780 45.180 ;
      LAYER met2 ;
        RECT 444.350 400.250 444.630 404.000 ;
        RECT 443.140 400.110 444.630 400.250 ;
        RECT 443.140 324.370 443.280 400.110 ;
        RECT 444.350 400.000 444.630 400.110 ;
        RECT 442.680 324.230 443.280 324.370 ;
        RECT 442.680 45.210 442.820 324.230 ;
        RECT 442.620 44.890 442.880 45.210 ;
        RECT 794.520 44.890 794.780 45.210 ;
        RECT 794.580 2.400 794.720 44.890 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.750 40.020 395.070 40.080 ;
        RECT 640.850 40.020 641.170 40.080 ;
        RECT 394.750 39.880 641.170 40.020 ;
        RECT 394.750 39.820 395.070 39.880 ;
        RECT 640.850 39.820 641.170 39.880 ;
      LAYER via ;
        RECT 394.780 39.820 395.040 40.080 ;
        RECT 640.880 39.820 641.140 40.080 ;
      LAYER met2 ;
        RECT 396.970 400.250 397.250 404.000 ;
        RECT 395.760 400.110 397.250 400.250 ;
        RECT 395.760 324.370 395.900 400.110 ;
        RECT 396.970 400.000 397.250 400.110 ;
        RECT 394.840 324.230 395.900 324.370 ;
        RECT 394.840 40.110 394.980 324.230 ;
        RECT 394.780 39.790 395.040 40.110 ;
        RECT 640.880 39.790 641.140 40.110 ;
        RECT 640.940 2.400 641.080 39.790 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 939.390 376.280 939.710 376.340 ;
        RECT 942.610 376.280 942.930 376.340 ;
        RECT 939.390 376.140 942.930 376.280 ;
        RECT 939.390 376.080 939.710 376.140 ;
        RECT 942.610 376.080 942.930 376.140 ;
        RECT 939.390 85.580 939.710 85.640 ;
        RECT 2408.170 85.580 2408.490 85.640 ;
        RECT 939.390 85.440 2408.490 85.580 ;
        RECT 939.390 85.380 939.710 85.440 ;
        RECT 2408.170 85.380 2408.490 85.440 ;
        RECT 2408.170 17.580 2408.490 17.640 ;
        RECT 2412.310 17.580 2412.630 17.640 ;
        RECT 2408.170 17.440 2412.630 17.580 ;
        RECT 2408.170 17.380 2408.490 17.440 ;
        RECT 2412.310 17.380 2412.630 17.440 ;
      LAYER via ;
        RECT 939.420 376.080 939.680 376.340 ;
        RECT 942.640 376.080 942.900 376.340 ;
        RECT 939.420 85.380 939.680 85.640 ;
        RECT 2408.200 85.380 2408.460 85.640 ;
        RECT 2408.200 17.380 2408.460 17.640 ;
        RECT 2412.340 17.380 2412.600 17.640 ;
      LAYER met2 ;
        RECT 943.910 400.250 944.190 404.000 ;
        RECT 942.700 400.110 944.190 400.250 ;
        RECT 942.700 376.370 942.840 400.110 ;
        RECT 943.910 400.000 944.190 400.110 ;
        RECT 939.420 376.050 939.680 376.370 ;
        RECT 942.640 376.050 942.900 376.370 ;
        RECT 939.480 85.670 939.620 376.050 ;
        RECT 939.420 85.350 939.680 85.670 ;
        RECT 2408.200 85.350 2408.460 85.670 ;
        RECT 2408.260 17.670 2408.400 85.350 ;
        RECT 2408.200 17.350 2408.460 17.670 ;
        RECT 2412.340 17.350 2412.600 17.670 ;
        RECT 2412.400 1.770 2412.540 17.350 ;
        RECT 2414.030 1.770 2414.590 2.400 ;
        RECT 2412.400 1.630 2414.590 1.770 ;
        RECT 2414.030 -4.800 2414.590 1.630 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.830 376.620 946.150 376.680 ;
        RECT 948.130 376.620 948.450 376.680 ;
        RECT 945.830 376.480 948.450 376.620 ;
        RECT 945.830 376.420 946.150 376.480 ;
        RECT 948.130 376.420 948.450 376.480 ;
        RECT 945.830 85.920 946.150 85.980 ;
        RECT 2428.870 85.920 2429.190 85.980 ;
        RECT 945.830 85.780 2429.190 85.920 ;
        RECT 945.830 85.720 946.150 85.780 ;
        RECT 2428.870 85.720 2429.190 85.780 ;
      LAYER via ;
        RECT 945.860 376.420 946.120 376.680 ;
        RECT 948.160 376.420 948.420 376.680 ;
        RECT 945.860 85.720 946.120 85.980 ;
        RECT 2428.900 85.720 2429.160 85.980 ;
      LAYER met2 ;
        RECT 949.430 400.250 949.710 404.000 ;
        RECT 948.220 400.110 949.710 400.250 ;
        RECT 948.220 376.710 948.360 400.110 ;
        RECT 949.430 400.000 949.710 400.110 ;
        RECT 945.860 376.390 946.120 376.710 ;
        RECT 948.160 376.390 948.420 376.710 ;
        RECT 945.920 86.010 946.060 376.390 ;
        RECT 945.860 85.690 946.120 86.010 ;
        RECT 2428.900 85.690 2429.160 86.010 ;
        RECT 2428.960 82.870 2429.100 85.690 ;
        RECT 2428.960 82.730 2432.320 82.870 ;
        RECT 2432.180 2.400 2432.320 82.730 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 953.190 89.660 953.510 89.720 ;
        RECT 2450.030 89.660 2450.350 89.720 ;
        RECT 953.190 89.520 2450.350 89.660 ;
        RECT 953.190 89.460 953.510 89.520 ;
        RECT 2450.030 89.460 2450.350 89.520 ;
      LAYER via ;
        RECT 953.220 89.460 953.480 89.720 ;
        RECT 2450.060 89.460 2450.320 89.720 ;
      LAYER met2 ;
        RECT 954.950 400.250 955.230 404.000 ;
        RECT 953.740 400.110 955.230 400.250 ;
        RECT 953.740 351.970 953.880 400.110 ;
        RECT 954.950 400.000 955.230 400.110 ;
        RECT 953.280 351.830 953.880 351.970 ;
        RECT 953.280 89.750 953.420 351.830 ;
        RECT 953.220 89.430 953.480 89.750 ;
        RECT 2450.060 89.430 2450.320 89.750 ;
        RECT 2450.120 16.730 2450.260 89.430 ;
        RECT 2449.660 16.590 2450.260 16.730 ;
        RECT 2449.660 2.400 2449.800 16.590 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.630 89.320 959.950 89.380 ;
        RECT 2463.370 89.320 2463.690 89.380 ;
        RECT 959.630 89.180 2463.690 89.320 ;
        RECT 959.630 89.120 959.950 89.180 ;
        RECT 2463.370 89.120 2463.690 89.180 ;
      LAYER via ;
        RECT 959.660 89.120 959.920 89.380 ;
        RECT 2463.400 89.120 2463.660 89.380 ;
      LAYER met2 ;
        RECT 960.010 400.250 960.290 404.000 ;
        RECT 959.720 400.110 960.290 400.250 ;
        RECT 959.720 89.410 959.860 400.110 ;
        RECT 960.010 400.000 960.290 400.110 ;
        RECT 959.660 89.090 959.920 89.410 ;
        RECT 2463.400 89.090 2463.660 89.410 ;
        RECT 2463.460 82.870 2463.600 89.090 ;
        RECT 2463.460 82.730 2465.440 82.870 ;
        RECT 2465.300 1.770 2465.440 82.730 ;
        RECT 2467.390 1.770 2467.950 2.400 ;
        RECT 2465.300 1.630 2467.950 1.770 ;
        RECT 2467.390 -4.800 2467.950 1.630 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.090 376.280 960.410 376.340 ;
        RECT 964.230 376.280 964.550 376.340 ;
        RECT 960.090 376.140 964.550 376.280 ;
        RECT 960.090 376.080 960.410 376.140 ;
        RECT 964.230 376.080 964.550 376.140 ;
        RECT 960.090 88.980 960.410 89.040 ;
        RECT 2484.070 88.980 2484.390 89.040 ;
        RECT 960.090 88.840 2484.390 88.980 ;
        RECT 960.090 88.780 960.410 88.840 ;
        RECT 2484.070 88.780 2484.390 88.840 ;
      LAYER via ;
        RECT 960.120 376.080 960.380 376.340 ;
        RECT 964.260 376.080 964.520 376.340 ;
        RECT 960.120 88.780 960.380 89.040 ;
        RECT 2484.100 88.780 2484.360 89.040 ;
      LAYER met2 ;
        RECT 965.530 400.250 965.810 404.000 ;
        RECT 964.320 400.110 965.810 400.250 ;
        RECT 964.320 376.370 964.460 400.110 ;
        RECT 965.530 400.000 965.810 400.110 ;
        RECT 960.120 376.050 960.380 376.370 ;
        RECT 964.260 376.050 964.520 376.370 ;
        RECT 960.180 89.070 960.320 376.050 ;
        RECT 960.120 88.750 960.380 89.070 ;
        RECT 2484.100 88.750 2484.360 89.070 ;
        RECT 2484.160 82.870 2484.300 88.750 ;
        RECT 2484.160 82.730 2485.680 82.870 ;
        RECT 2485.540 2.400 2485.680 82.730 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.990 88.640 967.310 88.700 ;
        RECT 2497.870 88.640 2498.190 88.700 ;
        RECT 966.990 88.500 2498.190 88.640 ;
        RECT 966.990 88.440 967.310 88.500 ;
        RECT 2497.870 88.440 2498.190 88.500 ;
      LAYER via ;
        RECT 967.020 88.440 967.280 88.700 ;
        RECT 2497.900 88.440 2498.160 88.700 ;
      LAYER met2 ;
        RECT 971.050 400.250 971.330 404.000 ;
        RECT 969.840 400.110 971.330 400.250 ;
        RECT 969.840 324.370 969.980 400.110 ;
        RECT 971.050 400.000 971.330 400.110 ;
        RECT 967.080 324.230 969.980 324.370 ;
        RECT 967.080 88.730 967.220 324.230 ;
        RECT 967.020 88.410 967.280 88.730 ;
        RECT 2497.900 88.410 2498.160 88.730 ;
        RECT 2497.960 82.870 2498.100 88.410 ;
        RECT 2497.960 82.730 2503.160 82.870 ;
        RECT 2503.020 2.400 2503.160 82.730 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 974.350 88.300 974.670 88.360 ;
        RECT 2518.570 88.300 2518.890 88.360 ;
        RECT 974.350 88.160 2518.890 88.300 ;
        RECT 974.350 88.100 974.670 88.160 ;
        RECT 2518.570 88.100 2518.890 88.160 ;
      LAYER via ;
        RECT 974.380 88.100 974.640 88.360 ;
        RECT 2518.600 88.100 2518.860 88.360 ;
      LAYER met2 ;
        RECT 976.570 400.250 976.850 404.000 ;
        RECT 975.360 400.110 976.850 400.250 ;
        RECT 975.360 324.370 975.500 400.110 ;
        RECT 976.570 400.000 976.850 400.110 ;
        RECT 974.440 324.230 975.500 324.370 ;
        RECT 974.440 88.390 974.580 324.230 ;
        RECT 974.380 88.070 974.640 88.390 ;
        RECT 2518.600 88.070 2518.860 88.390 ;
        RECT 2518.660 1.770 2518.800 88.070 ;
        RECT 2520.750 1.770 2521.310 2.400 ;
        RECT 2518.660 1.630 2521.310 1.770 ;
        RECT 2520.750 -4.800 2521.310 1.630 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.330 376.280 980.650 376.340 ;
        RECT 981.250 376.280 981.570 376.340 ;
        RECT 980.330 376.140 981.570 376.280 ;
        RECT 980.330 376.080 980.650 376.140 ;
        RECT 981.250 376.080 981.570 376.140 ;
        RECT 980.330 87.960 980.650 88.020 ;
        RECT 2532.830 87.960 2533.150 88.020 ;
        RECT 980.330 87.820 2533.150 87.960 ;
        RECT 980.330 87.760 980.650 87.820 ;
        RECT 2532.830 87.760 2533.150 87.820 ;
      LAYER via ;
        RECT 980.360 376.080 980.620 376.340 ;
        RECT 981.280 376.080 981.540 376.340 ;
        RECT 980.360 87.760 980.620 88.020 ;
        RECT 2532.860 87.760 2533.120 88.020 ;
      LAYER met2 ;
        RECT 982.090 400.250 982.370 404.000 ;
        RECT 981.340 400.110 982.370 400.250 ;
        RECT 981.340 376.370 981.480 400.110 ;
        RECT 982.090 400.000 982.370 400.110 ;
        RECT 980.360 376.050 980.620 376.370 ;
        RECT 981.280 376.050 981.540 376.370 ;
        RECT 980.420 88.050 980.560 376.050 ;
        RECT 980.360 87.730 980.620 88.050 ;
        RECT 2532.860 87.730 2533.120 88.050 ;
        RECT 2532.920 82.870 2533.060 87.730 ;
        RECT 2532.920 82.730 2536.280 82.870 ;
        RECT 2536.140 1.770 2536.280 82.730 ;
        RECT 2538.230 1.770 2538.790 2.400 ;
        RECT 2536.140 1.630 2538.790 1.770 ;
        RECT 2538.230 -4.800 2538.790 1.630 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.230 87.620 987.550 87.680 ;
        RECT 2553.070 87.620 2553.390 87.680 ;
        RECT 987.230 87.480 2553.390 87.620 ;
        RECT 987.230 87.420 987.550 87.480 ;
        RECT 2553.070 87.420 2553.390 87.480 ;
      LAYER via ;
        RECT 987.260 87.420 987.520 87.680 ;
        RECT 2553.100 87.420 2553.360 87.680 ;
      LAYER met2 ;
        RECT 987.610 400.250 987.890 404.000 ;
        RECT 987.320 400.110 987.890 400.250 ;
        RECT 987.320 87.710 987.460 400.110 ;
        RECT 987.610 400.000 987.890 400.110 ;
        RECT 987.260 87.390 987.520 87.710 ;
        RECT 2553.100 87.390 2553.360 87.710 ;
        RECT 2553.160 82.870 2553.300 87.390 ;
        RECT 2553.160 82.730 2556.520 82.870 ;
        RECT 2556.380 2.400 2556.520 82.730 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.690 375.940 988.010 376.000 ;
        RECT 991.830 375.940 992.150 376.000 ;
        RECT 987.690 375.800 992.150 375.940 ;
        RECT 987.690 375.740 988.010 375.800 ;
        RECT 991.830 375.740 992.150 375.800 ;
        RECT 987.690 87.280 988.010 87.340 ;
        RECT 2573.770 87.280 2574.090 87.340 ;
        RECT 987.690 87.140 2574.090 87.280 ;
        RECT 987.690 87.080 988.010 87.140 ;
        RECT 2573.770 87.080 2574.090 87.140 ;
      LAYER via ;
        RECT 987.720 375.740 987.980 376.000 ;
        RECT 991.860 375.740 992.120 376.000 ;
        RECT 987.720 87.080 987.980 87.340 ;
        RECT 2573.800 87.080 2574.060 87.340 ;
      LAYER met2 ;
        RECT 993.130 400.250 993.410 404.000 ;
        RECT 991.920 400.110 993.410 400.250 ;
        RECT 991.920 376.030 992.060 400.110 ;
        RECT 993.130 400.000 993.410 400.110 ;
        RECT 987.720 375.710 987.980 376.030 ;
        RECT 991.860 375.710 992.120 376.030 ;
        RECT 987.780 87.370 987.920 375.710 ;
        RECT 987.720 87.050 987.980 87.370 ;
        RECT 2573.800 87.050 2574.060 87.370 ;
        RECT 2573.860 2.400 2574.000 87.050 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 44.780 449.350 44.840 ;
        RECT 818.410 44.780 818.730 44.840 ;
        RECT 449.030 44.640 818.730 44.780 ;
        RECT 449.030 44.580 449.350 44.640 ;
        RECT 818.410 44.580 818.730 44.640 ;
      LAYER via ;
        RECT 449.060 44.580 449.320 44.840 ;
        RECT 818.440 44.580 818.700 44.840 ;
      LAYER met2 ;
        RECT 451.710 400.250 451.990 404.000 ;
        RECT 450.500 400.110 451.990 400.250 ;
        RECT 450.500 324.370 450.640 400.110 ;
        RECT 451.710 400.000 451.990 400.110 ;
        RECT 449.120 324.230 450.640 324.370 ;
        RECT 449.120 44.870 449.260 324.230 ;
        RECT 449.060 44.550 449.320 44.870 ;
        RECT 818.440 44.550 818.700 44.870 ;
        RECT 818.500 2.400 818.640 44.550 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.130 376.280 994.450 376.340 ;
        RECT 997.350 376.280 997.670 376.340 ;
        RECT 994.130 376.140 997.670 376.280 ;
        RECT 994.130 376.080 994.450 376.140 ;
        RECT 997.350 376.080 997.670 376.140 ;
        RECT 994.130 86.940 994.450 87.000 ;
        RECT 2587.570 86.940 2587.890 87.000 ;
        RECT 994.130 86.800 2587.890 86.940 ;
        RECT 994.130 86.740 994.450 86.800 ;
        RECT 2587.570 86.740 2587.890 86.800 ;
      LAYER via ;
        RECT 994.160 376.080 994.420 376.340 ;
        RECT 997.380 376.080 997.640 376.340 ;
        RECT 994.160 86.740 994.420 87.000 ;
        RECT 2587.600 86.740 2587.860 87.000 ;
      LAYER met2 ;
        RECT 998.650 400.250 998.930 404.000 ;
        RECT 997.440 400.110 998.930 400.250 ;
        RECT 997.440 376.370 997.580 400.110 ;
        RECT 998.650 400.000 998.930 400.110 ;
        RECT 994.160 376.050 994.420 376.370 ;
        RECT 997.380 376.050 997.640 376.370 ;
        RECT 994.220 87.030 994.360 376.050 ;
        RECT 994.160 86.710 994.420 87.030 ;
        RECT 2587.600 86.710 2587.860 87.030 ;
        RECT 2587.660 82.870 2587.800 86.710 ;
        RECT 2587.660 82.730 2589.640 82.870 ;
        RECT 2589.500 1.770 2589.640 82.730 ;
        RECT 2591.590 1.770 2592.150 2.400 ;
        RECT 2589.500 1.630 2592.150 1.770 ;
        RECT 2591.590 -4.800 2592.150 1.630 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.950 86.600 1002.270 86.660 ;
        RECT 2608.270 86.600 2608.590 86.660 ;
        RECT 1001.950 86.460 2608.590 86.600 ;
        RECT 1001.950 86.400 1002.270 86.460 ;
        RECT 2608.270 86.400 2608.590 86.460 ;
      LAYER via ;
        RECT 1001.980 86.400 1002.240 86.660 ;
        RECT 2608.300 86.400 2608.560 86.660 ;
      LAYER met2 ;
        RECT 1004.170 400.250 1004.450 404.000 ;
        RECT 1002.960 400.110 1004.450 400.250 ;
        RECT 1002.960 324.370 1003.100 400.110 ;
        RECT 1004.170 400.000 1004.450 400.110 ;
        RECT 1002.040 324.230 1003.100 324.370 ;
        RECT 1002.040 86.690 1002.180 324.230 ;
        RECT 1001.980 86.370 1002.240 86.690 ;
        RECT 2608.300 86.370 2608.560 86.690 ;
        RECT 2608.360 1.770 2608.500 86.370 ;
        RECT 2609.070 1.770 2609.630 2.400 ;
        RECT 2608.360 1.630 2609.630 1.770 ;
        RECT 2609.070 -4.800 2609.630 1.630 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1008.850 86.260 1009.170 86.320 ;
        RECT 2622.070 86.260 2622.390 86.320 ;
        RECT 1008.850 86.120 2622.390 86.260 ;
        RECT 1008.850 86.060 1009.170 86.120 ;
        RECT 2622.070 86.060 2622.390 86.120 ;
      LAYER via ;
        RECT 1008.880 86.060 1009.140 86.320 ;
        RECT 2622.100 86.060 2622.360 86.320 ;
      LAYER met2 ;
        RECT 1009.230 400.250 1009.510 404.000 ;
        RECT 1008.940 400.110 1009.510 400.250 ;
        RECT 1008.940 86.350 1009.080 400.110 ;
        RECT 1009.230 400.000 1009.510 400.110 ;
        RECT 1008.880 86.030 1009.140 86.350 ;
        RECT 2622.100 86.030 2622.360 86.350 ;
        RECT 2622.160 82.870 2622.300 86.030 ;
        RECT 2622.160 82.730 2627.360 82.870 ;
        RECT 2627.220 2.400 2627.360 82.730 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.750 400.180 1015.030 404.000 ;
        RECT 1014.750 400.000 1015.060 400.180 ;
        RECT 1014.920 377.130 1015.060 400.000 ;
        RECT 1014.920 376.990 1015.520 377.130 ;
        RECT 1015.380 86.885 1015.520 376.990 ;
        RECT 1015.310 86.515 1015.590 86.885 ;
        RECT 2642.790 86.515 2643.070 86.885 ;
        RECT 2642.860 1.770 2643.000 86.515 ;
        RECT 2644.950 1.770 2645.510 2.400 ;
        RECT 2642.860 1.630 2645.510 1.770 ;
        RECT 2644.950 -4.800 2645.510 1.630 ;
      LAYER via2 ;
        RECT 1015.310 86.560 1015.590 86.840 ;
        RECT 2642.790 86.560 2643.070 86.840 ;
      LAYER met3 ;
        RECT 1015.285 86.850 1015.615 86.865 ;
        RECT 2642.765 86.850 2643.095 86.865 ;
        RECT 1015.285 86.550 2643.095 86.850 ;
        RECT 1015.285 86.535 1015.615 86.550 ;
        RECT 2642.765 86.535 2643.095 86.550 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2656.570 17.580 2656.890 17.640 ;
        RECT 2660.710 17.580 2661.030 17.640 ;
        RECT 2656.570 17.440 2661.030 17.580 ;
        RECT 2656.570 17.380 2656.890 17.440 ;
        RECT 2660.710 17.380 2661.030 17.440 ;
      LAYER via ;
        RECT 2656.600 17.380 2656.860 17.640 ;
        RECT 2660.740 17.380 2661.000 17.640 ;
      LAYER met2 ;
        RECT 1020.270 400.250 1020.550 404.000 ;
        RECT 1019.060 400.110 1020.550 400.250 ;
        RECT 1019.060 324.370 1019.200 400.110 ;
        RECT 1020.270 400.000 1020.550 400.110 ;
        RECT 1016.300 324.230 1019.200 324.370 ;
        RECT 1016.300 86.205 1016.440 324.230 ;
        RECT 1016.230 85.835 1016.510 86.205 ;
        RECT 2656.590 85.835 2656.870 86.205 ;
        RECT 2656.660 17.670 2656.800 85.835 ;
        RECT 2656.600 17.350 2656.860 17.670 ;
        RECT 2660.740 17.350 2661.000 17.670 ;
        RECT 2660.800 1.770 2660.940 17.350 ;
        RECT 2662.430 1.770 2662.990 2.400 ;
        RECT 2660.800 1.630 2662.990 1.770 ;
        RECT 2662.430 -4.800 2662.990 1.630 ;
      LAYER via2 ;
        RECT 1016.230 85.880 1016.510 86.160 ;
        RECT 2656.590 85.880 2656.870 86.160 ;
      LAYER met3 ;
        RECT 1016.205 86.170 1016.535 86.185 ;
        RECT 2656.565 86.170 2656.895 86.185 ;
        RECT 1016.205 85.870 2656.895 86.170 ;
        RECT 1016.205 85.855 1016.535 85.870 ;
        RECT 2656.565 85.855 2656.895 85.870 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.650 120.940 1022.970 121.000 ;
        RECT 2677.270 120.940 2677.590 121.000 ;
        RECT 1022.650 120.800 2677.590 120.940 ;
        RECT 1022.650 120.740 1022.970 120.800 ;
        RECT 2677.270 120.740 2677.590 120.800 ;
      LAYER via ;
        RECT 1022.680 120.740 1022.940 121.000 ;
        RECT 2677.300 120.740 2677.560 121.000 ;
      LAYER met2 ;
        RECT 1025.790 400.250 1026.070 404.000 ;
        RECT 1024.580 400.110 1026.070 400.250 ;
        RECT 1024.580 324.370 1024.720 400.110 ;
        RECT 1025.790 400.000 1026.070 400.110 ;
        RECT 1022.740 324.230 1024.720 324.370 ;
        RECT 1022.740 121.030 1022.880 324.230 ;
        RECT 1022.680 120.710 1022.940 121.030 ;
        RECT 2677.300 120.710 2677.560 121.030 ;
        RECT 2677.360 82.870 2677.500 120.710 ;
        RECT 2677.360 82.730 2680.720 82.870 ;
        RECT 2680.580 2.400 2680.720 82.730 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1029.090 120.600 1029.410 120.660 ;
        RECT 2697.970 120.600 2698.290 120.660 ;
        RECT 1029.090 120.460 2698.290 120.600 ;
        RECT 1029.090 120.400 1029.410 120.460 ;
        RECT 2697.970 120.400 2698.290 120.460 ;
      LAYER via ;
        RECT 1029.120 120.400 1029.380 120.660 ;
        RECT 2698.000 120.400 2698.260 120.660 ;
      LAYER met2 ;
        RECT 1031.310 400.250 1031.590 404.000 ;
        RECT 1030.100 400.110 1031.590 400.250 ;
        RECT 1030.100 324.370 1030.240 400.110 ;
        RECT 1031.310 400.000 1031.590 400.110 ;
        RECT 1029.180 324.230 1030.240 324.370 ;
        RECT 1029.180 120.690 1029.320 324.230 ;
        RECT 1029.120 120.370 1029.380 120.690 ;
        RECT 2698.000 120.370 2698.260 120.690 ;
        RECT 2698.060 2.400 2698.200 120.370 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.830 400.250 1037.110 404.000 ;
        RECT 1036.540 400.110 1037.110 400.250 ;
        RECT 1036.540 121.565 1036.680 400.110 ;
        RECT 1036.830 400.000 1037.110 400.110 ;
        RECT 1036.470 121.195 1036.750 121.565 ;
        RECT 2711.790 121.195 2712.070 121.565 ;
        RECT 2711.860 82.870 2712.000 121.195 ;
        RECT 2711.860 82.730 2713.840 82.870 ;
        RECT 2713.700 1.770 2713.840 82.730 ;
        RECT 2715.790 1.770 2716.350 2.400 ;
        RECT 2713.700 1.630 2716.350 1.770 ;
        RECT 2715.790 -4.800 2716.350 1.630 ;
      LAYER via2 ;
        RECT 1036.470 121.240 1036.750 121.520 ;
        RECT 2711.790 121.240 2712.070 121.520 ;
      LAYER met3 ;
        RECT 1036.445 121.530 1036.775 121.545 ;
        RECT 2711.765 121.530 2712.095 121.545 ;
        RECT 1036.445 121.230 2712.095 121.530 ;
        RECT 1036.445 121.215 1036.775 121.230 ;
        RECT 2711.765 121.215 2712.095 121.230 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.350 400.250 1042.630 404.000 ;
        RECT 1042.350 400.110 1044.040 400.250 ;
        RECT 1042.350 400.000 1042.630 400.110 ;
        RECT 1043.900 351.970 1044.040 400.110 ;
        RECT 1043.900 351.830 1044.500 351.970 ;
        RECT 1044.360 324.370 1044.500 351.830 ;
        RECT 1043.440 324.230 1044.500 324.370 ;
        RECT 1043.440 120.885 1043.580 324.230 ;
        RECT 1043.370 120.515 1043.650 120.885 ;
        RECT 2732.490 120.515 2732.770 120.885 ;
        RECT 2732.560 1.770 2732.700 120.515 ;
        RECT 2733.270 1.770 2733.830 2.400 ;
        RECT 2732.560 1.630 2733.830 1.770 ;
        RECT 2733.270 -4.800 2733.830 1.630 ;
      LAYER via2 ;
        RECT 1043.370 120.560 1043.650 120.840 ;
        RECT 2732.490 120.560 2732.770 120.840 ;
      LAYER met3 ;
        RECT 1043.345 120.850 1043.675 120.865 ;
        RECT 2732.465 120.850 2732.795 120.865 ;
        RECT 1043.345 120.550 2732.795 120.850 ;
        RECT 1043.345 120.535 1043.675 120.550 ;
        RECT 2732.465 120.535 2732.795 120.550 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.890 376.280 1043.210 376.340 ;
        RECT 1046.570 376.280 1046.890 376.340 ;
        RECT 1042.890 376.140 1046.890 376.280 ;
        RECT 1042.890 376.080 1043.210 376.140 ;
        RECT 1046.570 376.080 1046.890 376.140 ;
        RECT 1042.890 94.760 1043.210 94.820 ;
        RECT 2746.270 94.760 2746.590 94.820 ;
        RECT 1042.890 94.620 2746.590 94.760 ;
        RECT 1042.890 94.560 1043.210 94.620 ;
        RECT 2746.270 94.560 2746.590 94.620 ;
      LAYER via ;
        RECT 1042.920 376.080 1043.180 376.340 ;
        RECT 1046.600 376.080 1046.860 376.340 ;
        RECT 1042.920 94.560 1043.180 94.820 ;
        RECT 2746.300 94.560 2746.560 94.820 ;
      LAYER met2 ;
        RECT 1047.870 400.250 1048.150 404.000 ;
        RECT 1046.660 400.110 1048.150 400.250 ;
        RECT 1046.660 376.370 1046.800 400.110 ;
        RECT 1047.870 400.000 1048.150 400.110 ;
        RECT 1042.920 376.050 1043.180 376.370 ;
        RECT 1046.600 376.050 1046.860 376.370 ;
        RECT 1042.980 94.850 1043.120 376.050 ;
        RECT 1042.920 94.530 1043.180 94.850 ;
        RECT 2746.300 94.530 2746.560 94.850 ;
        RECT 2746.360 82.870 2746.500 94.530 ;
        RECT 2746.360 82.730 2751.560 82.870 ;
        RECT 2751.420 2.400 2751.560 82.730 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 42.740 456.710 42.800 ;
        RECT 835.890 42.740 836.210 42.800 ;
        RECT 456.390 42.600 836.210 42.740 ;
        RECT 456.390 42.540 456.710 42.600 ;
        RECT 835.890 42.540 836.210 42.600 ;
      LAYER via ;
        RECT 456.420 42.540 456.680 42.800 ;
        RECT 835.920 42.540 836.180 42.800 ;
      LAYER met2 ;
        RECT 457.230 400.250 457.510 404.000 ;
        RECT 456.480 400.110 457.510 400.250 ;
        RECT 456.480 42.830 456.620 400.110 ;
        RECT 457.230 400.000 457.510 400.110 ;
        RECT 456.420 42.510 456.680 42.830 ;
        RECT 835.920 42.510 836.180 42.830 ;
        RECT 835.980 2.400 836.120 42.510 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1050.250 94.420 1050.570 94.480 ;
        RECT 2766.970 94.420 2767.290 94.480 ;
        RECT 1050.250 94.280 2767.290 94.420 ;
        RECT 1050.250 94.220 1050.570 94.280 ;
        RECT 2766.970 94.220 2767.290 94.280 ;
      LAYER via ;
        RECT 1050.280 94.220 1050.540 94.480 ;
        RECT 2767.000 94.220 2767.260 94.480 ;
      LAYER met2 ;
        RECT 1053.390 400.250 1053.670 404.000 ;
        RECT 1052.180 400.110 1053.670 400.250 ;
        RECT 1052.180 351.970 1052.320 400.110 ;
        RECT 1053.390 400.000 1053.670 400.110 ;
        RECT 1050.340 351.830 1052.320 351.970 ;
        RECT 1050.340 94.510 1050.480 351.830 ;
        RECT 1050.280 94.190 1050.540 94.510 ;
        RECT 2767.000 94.190 2767.260 94.510 ;
        RECT 2767.060 82.870 2767.200 94.190 ;
        RECT 2767.060 82.730 2769.040 82.870 ;
        RECT 2768.900 2.400 2769.040 82.730 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1056.690 94.080 1057.010 94.140 ;
        RECT 2780.770 94.080 2781.090 94.140 ;
        RECT 1056.690 93.940 2781.090 94.080 ;
        RECT 1056.690 93.880 1057.010 93.940 ;
        RECT 2780.770 93.880 2781.090 93.940 ;
        RECT 2780.770 17.580 2781.090 17.640 ;
        RECT 2784.910 17.580 2785.230 17.640 ;
        RECT 2780.770 17.440 2785.230 17.580 ;
        RECT 2780.770 17.380 2781.090 17.440 ;
        RECT 2784.910 17.380 2785.230 17.440 ;
      LAYER via ;
        RECT 1056.720 93.880 1056.980 94.140 ;
        RECT 2780.800 93.880 2781.060 94.140 ;
        RECT 2780.800 17.380 2781.060 17.640 ;
        RECT 2784.940 17.380 2785.200 17.640 ;
      LAYER met2 ;
        RECT 1058.450 400.250 1058.730 404.000 ;
        RECT 1057.240 400.110 1058.730 400.250 ;
        RECT 1057.240 351.970 1057.380 400.110 ;
        RECT 1058.450 400.000 1058.730 400.110 ;
        RECT 1056.780 351.830 1057.380 351.970 ;
        RECT 1056.780 94.170 1056.920 351.830 ;
        RECT 1056.720 93.850 1056.980 94.170 ;
        RECT 2780.800 93.850 2781.060 94.170 ;
        RECT 2780.860 17.670 2781.000 93.850 ;
        RECT 2780.800 17.350 2781.060 17.670 ;
        RECT 2784.940 17.350 2785.200 17.670 ;
        RECT 2785.000 1.770 2785.140 17.350 ;
        RECT 2786.630 1.770 2787.190 2.400 ;
        RECT 2785.000 1.630 2787.190 1.770 ;
        RECT 2786.630 -4.800 2787.190 1.630 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.130 93.740 1063.450 93.800 ;
        RECT 2801.470 93.740 2801.790 93.800 ;
        RECT 1063.130 93.600 2801.790 93.740 ;
        RECT 1063.130 93.540 1063.450 93.600 ;
        RECT 2801.470 93.540 2801.790 93.600 ;
      LAYER via ;
        RECT 1063.160 93.540 1063.420 93.800 ;
        RECT 2801.500 93.540 2801.760 93.800 ;
      LAYER met2 ;
        RECT 1063.970 400.250 1064.250 404.000 ;
        RECT 1063.220 400.110 1064.250 400.250 ;
        RECT 1063.220 93.830 1063.360 400.110 ;
        RECT 1063.970 400.000 1064.250 400.110 ;
        RECT 1063.160 93.510 1063.420 93.830 ;
        RECT 2801.500 93.510 2801.760 93.830 ;
        RECT 2801.560 82.870 2801.700 93.510 ;
        RECT 2801.560 82.730 2802.160 82.870 ;
        RECT 2802.020 1.770 2802.160 82.730 ;
        RECT 2804.110 1.770 2804.670 2.400 ;
        RECT 2802.020 1.630 2804.670 1.770 ;
        RECT 2804.110 -4.800 2804.670 1.630 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.490 93.400 1070.810 93.460 ;
        RECT 2822.630 93.400 2822.950 93.460 ;
        RECT 1070.490 93.260 2822.950 93.400 ;
        RECT 1070.490 93.200 1070.810 93.260 ;
        RECT 2822.630 93.200 2822.950 93.260 ;
      LAYER via ;
        RECT 1070.520 93.200 1070.780 93.460 ;
        RECT 2822.660 93.200 2822.920 93.460 ;
      LAYER met2 ;
        RECT 1069.490 400.250 1069.770 404.000 ;
        RECT 1069.490 400.110 1070.720 400.250 ;
        RECT 1069.490 400.000 1069.770 400.110 ;
        RECT 1070.580 93.490 1070.720 400.110 ;
        RECT 1070.520 93.170 1070.780 93.490 ;
        RECT 2822.660 93.170 2822.920 93.490 ;
        RECT 2822.720 16.730 2822.860 93.170 ;
        RECT 2822.260 16.590 2822.860 16.730 ;
        RECT 2822.260 2.400 2822.400 16.590 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.030 376.280 1070.350 376.340 ;
        RECT 1073.710 376.280 1074.030 376.340 ;
        RECT 1070.030 376.140 1074.030 376.280 ;
        RECT 1070.030 376.080 1070.350 376.140 ;
        RECT 1073.710 376.080 1074.030 376.140 ;
        RECT 1070.030 93.060 1070.350 93.120 ;
        RECT 2835.970 93.060 2836.290 93.120 ;
        RECT 1070.030 92.920 2836.290 93.060 ;
        RECT 1070.030 92.860 1070.350 92.920 ;
        RECT 2835.970 92.860 2836.290 92.920 ;
      LAYER via ;
        RECT 1070.060 376.080 1070.320 376.340 ;
        RECT 1073.740 376.080 1074.000 376.340 ;
        RECT 1070.060 92.860 1070.320 93.120 ;
        RECT 2836.000 92.860 2836.260 93.120 ;
      LAYER met2 ;
        RECT 1075.010 400.250 1075.290 404.000 ;
        RECT 1073.800 400.110 1075.290 400.250 ;
        RECT 1073.800 376.370 1073.940 400.110 ;
        RECT 1075.010 400.000 1075.290 400.110 ;
        RECT 1070.060 376.050 1070.320 376.370 ;
        RECT 1073.740 376.050 1074.000 376.370 ;
        RECT 1070.120 93.150 1070.260 376.050 ;
        RECT 1070.060 92.830 1070.320 93.150 ;
        RECT 2836.000 92.830 2836.260 93.150 ;
        RECT 2836.060 82.870 2836.200 92.830 ;
        RECT 2836.060 82.730 2838.040 82.870 ;
        RECT 2837.900 1.770 2838.040 82.730 ;
        RECT 2839.990 1.770 2840.550 2.400 ;
        RECT 2837.900 1.630 2840.550 1.770 ;
        RECT 2839.990 -4.800 2840.550 1.630 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.530 400.250 1080.810 404.000 ;
        RECT 1079.320 400.110 1080.810 400.250 ;
        RECT 1079.320 324.370 1079.460 400.110 ;
        RECT 1080.530 400.000 1080.810 400.110 ;
        RECT 1077.940 324.230 1079.460 324.370 ;
        RECT 1077.940 93.685 1078.080 324.230 ;
        RECT 1077.870 93.315 1078.150 93.685 ;
        RECT 2856.690 93.315 2856.970 93.685 ;
        RECT 2856.760 1.770 2856.900 93.315 ;
        RECT 2857.470 1.770 2858.030 2.400 ;
        RECT 2856.760 1.630 2858.030 1.770 ;
        RECT 2857.470 -4.800 2858.030 1.630 ;
      LAYER via2 ;
        RECT 1077.870 93.360 1078.150 93.640 ;
        RECT 2856.690 93.360 2856.970 93.640 ;
      LAYER met3 ;
        RECT 1077.845 93.650 1078.175 93.665 ;
        RECT 2856.665 93.650 2856.995 93.665 ;
        RECT 1077.845 93.350 2856.995 93.650 ;
        RECT 1077.845 93.335 1078.175 93.350 ;
        RECT 2856.665 93.335 2856.995 93.350 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.050 400.250 1086.330 404.000 ;
        RECT 1084.840 400.110 1086.330 400.250 ;
        RECT 1084.840 93.005 1084.980 400.110 ;
        RECT 1086.050 400.000 1086.330 400.110 ;
        RECT 1084.770 92.635 1085.050 93.005 ;
        RECT 2870.490 92.635 2870.770 93.005 ;
        RECT 2870.560 82.870 2870.700 92.635 ;
        RECT 2870.560 82.730 2875.760 82.870 ;
        RECT 2875.620 2.400 2875.760 82.730 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
      LAYER via2 ;
        RECT 1084.770 92.680 1085.050 92.960 ;
        RECT 2870.490 92.680 2870.770 92.960 ;
      LAYER met3 ;
        RECT 1084.745 92.970 1085.075 92.985 ;
        RECT 2870.465 92.970 2870.795 92.985 ;
        RECT 1084.745 92.670 2870.795 92.970 ;
        RECT 1084.745 92.655 1085.075 92.670 ;
        RECT 2870.465 92.655 2870.795 92.670 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1090.270 30.840 1090.590 30.900 ;
        RECT 2893.010 30.840 2893.330 30.900 ;
        RECT 1090.270 30.700 2893.330 30.840 ;
        RECT 1090.270 30.640 1090.590 30.700 ;
        RECT 2893.010 30.640 2893.330 30.700 ;
      LAYER via ;
        RECT 1090.300 30.640 1090.560 30.900 ;
        RECT 2893.040 30.640 2893.300 30.900 ;
      LAYER met2 ;
        RECT 1091.570 400.250 1091.850 404.000 ;
        RECT 1090.360 400.110 1091.850 400.250 ;
        RECT 1090.360 30.930 1090.500 400.110 ;
        RECT 1091.570 400.000 1091.850 400.110 ;
        RECT 1090.300 30.610 1090.560 30.930 ;
        RECT 2893.040 30.610 2893.300 30.930 ;
        RECT 2893.100 2.400 2893.240 30.610 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 35.940 462.690 36.000 ;
        RECT 744.810 35.940 745.130 36.000 ;
        RECT 462.370 35.800 745.130 35.940 ;
        RECT 462.370 35.740 462.690 35.800 ;
        RECT 744.810 35.740 745.130 35.800 ;
        RECT 744.810 16.560 745.130 16.620 ;
        RECT 853.830 16.560 854.150 16.620 ;
        RECT 744.810 16.420 854.150 16.560 ;
        RECT 744.810 16.360 745.130 16.420 ;
        RECT 853.830 16.360 854.150 16.420 ;
      LAYER via ;
        RECT 462.400 35.740 462.660 36.000 ;
        RECT 744.840 35.740 745.100 36.000 ;
        RECT 744.840 16.360 745.100 16.620 ;
        RECT 853.860 16.360 854.120 16.620 ;
      LAYER met2 ;
        RECT 462.750 400.250 463.030 404.000 ;
        RECT 462.460 400.110 463.030 400.250 ;
        RECT 462.460 36.030 462.600 400.110 ;
        RECT 462.750 400.000 463.030 400.110 ;
        RECT 462.400 35.710 462.660 36.030 ;
        RECT 744.840 35.710 745.100 36.030 ;
        RECT 744.900 16.650 745.040 35.710 ;
        RECT 744.840 16.330 745.100 16.650 ;
        RECT 853.860 16.330 854.120 16.650 ;
        RECT 853.920 2.400 854.060 16.330 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 52.940 463.610 53.000 ;
        RECT 869.930 52.940 870.250 53.000 ;
        RECT 463.290 52.800 870.250 52.940 ;
        RECT 463.290 52.740 463.610 52.800 ;
        RECT 869.930 52.740 870.250 52.800 ;
      LAYER via ;
        RECT 463.320 52.740 463.580 53.000 ;
        RECT 869.960 52.740 870.220 53.000 ;
      LAYER met2 ;
        RECT 468.270 400.250 468.550 404.000 ;
        RECT 467.060 400.110 468.550 400.250 ;
        RECT 467.060 399.570 467.200 400.110 ;
        RECT 468.270 400.000 468.550 400.110 ;
        RECT 465.220 399.430 467.200 399.570 ;
        RECT 465.220 351.970 465.360 399.430 ;
        RECT 463.380 351.830 465.360 351.970 ;
        RECT 463.380 53.030 463.520 351.830 ;
        RECT 463.320 52.710 463.580 53.030 ;
        RECT 869.960 52.710 870.220 53.030 ;
        RECT 870.020 1.770 870.160 52.710 ;
        RECT 871.190 1.770 871.750 2.400 ;
        RECT 870.020 1.630 871.750 1.770 ;
        RECT 871.190 -4.800 871.750 1.630 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.730 52.600 470.050 52.660 ;
        RECT 889.250 52.600 889.570 52.660 ;
        RECT 469.730 52.460 889.570 52.600 ;
        RECT 469.730 52.400 470.050 52.460 ;
        RECT 889.250 52.400 889.570 52.460 ;
      LAYER via ;
        RECT 469.760 52.400 470.020 52.660 ;
        RECT 889.280 52.400 889.540 52.660 ;
      LAYER met2 ;
        RECT 473.790 400.250 474.070 404.000 ;
        RECT 472.580 400.110 474.070 400.250 ;
        RECT 472.580 324.370 472.720 400.110 ;
        RECT 473.790 400.000 474.070 400.110 ;
        RECT 469.820 324.230 472.720 324.370 ;
        RECT 469.820 52.690 469.960 324.230 ;
        RECT 469.760 52.370 470.020 52.690 ;
        RECT 889.280 52.370 889.540 52.690 ;
        RECT 889.340 2.400 889.480 52.370 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.090 51.920 477.410 51.980 ;
        RECT 904.890 51.920 905.210 51.980 ;
        RECT 477.090 51.780 905.210 51.920 ;
        RECT 477.090 51.720 477.410 51.780 ;
        RECT 904.890 51.720 905.210 51.780 ;
      LAYER via ;
        RECT 477.120 51.720 477.380 51.980 ;
        RECT 904.920 51.720 905.180 51.980 ;
      LAYER met2 ;
        RECT 479.310 400.250 479.590 404.000 ;
        RECT 478.100 400.110 479.590 400.250 ;
        RECT 478.100 324.370 478.240 400.110 ;
        RECT 479.310 400.000 479.590 400.110 ;
        RECT 477.180 324.230 478.240 324.370 ;
        RECT 477.180 52.010 477.320 324.230 ;
        RECT 477.120 51.690 477.380 52.010 ;
        RECT 904.920 51.690 905.180 52.010 ;
        RECT 904.980 1.770 905.120 51.690 ;
        RECT 907.070 1.770 907.630 2.400 ;
        RECT 904.980 1.630 907.630 1.770 ;
        RECT 907.070 -4.800 907.630 1.630 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 51.580 483.850 51.640 ;
        RECT 925.130 51.580 925.450 51.640 ;
        RECT 483.530 51.440 925.450 51.580 ;
        RECT 483.530 51.380 483.850 51.440 ;
        RECT 925.130 51.380 925.450 51.440 ;
      LAYER via ;
        RECT 483.560 51.380 483.820 51.640 ;
        RECT 925.160 51.380 925.420 51.640 ;
      LAYER met2 ;
        RECT 484.830 400.250 485.110 404.000 ;
        RECT 483.620 400.110 485.110 400.250 ;
        RECT 483.620 51.670 483.760 400.110 ;
        RECT 484.830 400.000 485.110 400.110 ;
        RECT 483.560 51.350 483.820 51.670 ;
        RECT 925.160 51.350 925.420 51.670 ;
        RECT 925.220 17.410 925.360 51.350 ;
        RECT 924.760 17.270 925.360 17.410 ;
        RECT 924.760 2.400 924.900 17.270 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 43.080 490.750 43.140 ;
        RECT 942.610 43.080 942.930 43.140 ;
        RECT 490.430 42.940 942.930 43.080 ;
        RECT 490.430 42.880 490.750 42.940 ;
        RECT 942.610 42.880 942.930 42.940 ;
      LAYER via ;
        RECT 490.460 42.880 490.720 43.140 ;
        RECT 942.640 42.880 942.900 43.140 ;
      LAYER met2 ;
        RECT 489.890 400.250 490.170 404.000 ;
        RECT 489.890 400.110 490.660 400.250 ;
        RECT 489.890 400.000 490.170 400.110 ;
        RECT 490.520 43.170 490.660 400.110 ;
        RECT 490.460 42.850 490.720 43.170 ;
        RECT 942.640 42.850 942.900 43.170 ;
        RECT 942.700 2.400 942.840 42.850 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.890 49.540 491.210 49.600 ;
        RECT 960.090 49.540 960.410 49.600 ;
        RECT 490.890 49.400 960.410 49.540 ;
        RECT 490.890 49.340 491.210 49.400 ;
        RECT 960.090 49.340 960.410 49.400 ;
      LAYER via ;
        RECT 490.920 49.340 491.180 49.600 ;
        RECT 960.120 49.340 960.380 49.600 ;
      LAYER met2 ;
        RECT 495.410 400.250 495.690 404.000 ;
        RECT 494.200 400.110 495.690 400.250 ;
        RECT 494.200 399.570 494.340 400.110 ;
        RECT 495.410 400.000 495.690 400.110 ;
        RECT 492.820 399.430 494.340 399.570 ;
        RECT 492.820 351.970 492.960 399.430 ;
        RECT 491.440 351.830 492.960 351.970 ;
        RECT 491.440 324.370 491.580 351.830 ;
        RECT 490.980 324.230 491.580 324.370 ;
        RECT 490.980 49.630 491.120 324.230 ;
        RECT 490.920 49.310 491.180 49.630 ;
        RECT 960.120 49.310 960.380 49.630 ;
        RECT 960.180 2.400 960.320 49.310 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 501.010 390.900 501.330 390.960 ;
        RECT 501.010 390.760 518.260 390.900 ;
        RECT 501.010 390.700 501.330 390.760 ;
        RECT 518.120 390.220 518.260 390.760 ;
        RECT 727.790 390.220 728.110 390.280 ;
        RECT 518.120 390.080 728.110 390.220 ;
        RECT 727.790 390.020 728.110 390.080 ;
        RECT 727.790 27.440 728.110 27.500 ;
        RECT 978.030 27.440 978.350 27.500 ;
        RECT 727.790 27.300 978.350 27.440 ;
        RECT 727.790 27.240 728.110 27.300 ;
        RECT 978.030 27.240 978.350 27.300 ;
      LAYER via ;
        RECT 501.040 390.700 501.300 390.960 ;
        RECT 727.820 390.020 728.080 390.280 ;
        RECT 727.820 27.240 728.080 27.500 ;
        RECT 978.060 27.240 978.320 27.500 ;
      LAYER met2 ;
        RECT 500.930 400.180 501.210 404.000 ;
        RECT 500.930 400.000 501.240 400.180 ;
        RECT 501.100 390.990 501.240 400.000 ;
        RECT 501.040 390.670 501.300 390.990 ;
        RECT 727.820 389.990 728.080 390.310 ;
        RECT 727.880 27.530 728.020 389.990 ;
        RECT 727.820 27.210 728.080 27.530 ;
        RECT 978.060 27.210 978.320 27.530 ;
        RECT 978.120 2.400 978.260 27.210 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.730 29.480 401.050 29.540 ;
        RECT 600.370 29.480 600.690 29.540 ;
        RECT 400.730 29.340 600.690 29.480 ;
        RECT 400.730 29.280 401.050 29.340 ;
        RECT 600.370 29.280 600.690 29.340 ;
        RECT 600.370 15.540 600.690 15.600 ;
        RECT 658.790 15.540 659.110 15.600 ;
        RECT 600.370 15.400 659.110 15.540 ;
        RECT 600.370 15.340 600.690 15.400 ;
        RECT 658.790 15.340 659.110 15.400 ;
      LAYER via ;
        RECT 400.760 29.280 401.020 29.540 ;
        RECT 600.400 29.280 600.660 29.540 ;
        RECT 600.400 15.340 600.660 15.600 ;
        RECT 658.820 15.340 659.080 15.600 ;
      LAYER met2 ;
        RECT 402.490 400.250 402.770 404.000 ;
        RECT 401.280 400.110 402.770 400.250 ;
        RECT 401.280 386.470 401.420 400.110 ;
        RECT 402.490 400.000 402.770 400.110 ;
        RECT 400.820 386.330 401.420 386.470 ;
        RECT 400.820 29.570 400.960 386.330 ;
        RECT 400.760 29.250 401.020 29.570 ;
        RECT 600.400 29.250 600.660 29.570 ;
        RECT 600.460 15.630 600.600 29.250 ;
        RECT 600.400 15.310 600.660 15.630 ;
        RECT 658.820 15.310 659.080 15.630 ;
        RECT 658.880 2.400 659.020 15.310 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 376.280 504.550 376.340 ;
        RECT 505.150 376.280 505.470 376.340 ;
        RECT 504.230 376.140 505.470 376.280 ;
        RECT 504.230 376.080 504.550 376.140 ;
        RECT 505.150 376.080 505.470 376.140 ;
        RECT 504.230 60.760 504.550 60.820 ;
        RECT 994.130 60.760 994.450 60.820 ;
        RECT 504.230 60.620 994.450 60.760 ;
        RECT 504.230 60.560 504.550 60.620 ;
        RECT 994.130 60.560 994.450 60.620 ;
      LAYER via ;
        RECT 504.260 376.080 504.520 376.340 ;
        RECT 505.180 376.080 505.440 376.340 ;
        RECT 504.260 60.560 504.520 60.820 ;
        RECT 994.160 60.560 994.420 60.820 ;
      LAYER met2 ;
        RECT 506.450 400.250 506.730 404.000 ;
        RECT 505.240 400.110 506.730 400.250 ;
        RECT 505.240 376.370 505.380 400.110 ;
        RECT 506.450 400.000 506.730 400.110 ;
        RECT 504.260 376.050 504.520 376.370 ;
        RECT 505.180 376.050 505.440 376.370 ;
        RECT 504.320 60.850 504.460 376.050 ;
        RECT 504.260 60.530 504.520 60.850 ;
        RECT 994.160 60.530 994.420 60.850 ;
        RECT 994.220 1.770 994.360 60.530 ;
        RECT 995.390 1.770 995.950 2.400 ;
        RECT 994.220 1.630 995.950 1.770 ;
        RECT 995.390 -4.800 995.950 1.630 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 60.420 511.450 60.480 ;
        RECT 1008.850 60.420 1009.170 60.480 ;
        RECT 511.130 60.280 1009.170 60.420 ;
        RECT 511.130 60.220 511.450 60.280 ;
        RECT 1008.850 60.220 1009.170 60.280 ;
      LAYER via ;
        RECT 511.160 60.220 511.420 60.480 ;
        RECT 1008.880 60.220 1009.140 60.480 ;
      LAYER met2 ;
        RECT 511.970 400.250 512.250 404.000 ;
        RECT 511.220 400.110 512.250 400.250 ;
        RECT 511.220 60.510 511.360 400.110 ;
        RECT 511.970 400.000 512.250 400.110 ;
        RECT 511.160 60.190 511.420 60.510 ;
        RECT 1008.880 60.190 1009.140 60.510 ;
        RECT 1008.940 17.410 1009.080 60.190 ;
        RECT 1008.940 17.270 1013.680 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.490 59.400 518.810 59.460 ;
        RECT 1030.930 59.400 1031.250 59.460 ;
        RECT 518.490 59.260 1031.250 59.400 ;
        RECT 518.490 59.200 518.810 59.260 ;
        RECT 1030.930 59.200 1031.250 59.260 ;
      LAYER via ;
        RECT 518.520 59.200 518.780 59.460 ;
        RECT 1030.960 59.200 1031.220 59.460 ;
      LAYER met2 ;
        RECT 517.490 400.250 517.770 404.000 ;
        RECT 517.490 400.110 518.720 400.250 ;
        RECT 517.490 400.000 517.770 400.110 ;
        RECT 518.580 59.490 518.720 400.110 ;
        RECT 518.520 59.170 518.780 59.490 ;
        RECT 1030.960 59.170 1031.220 59.490 ;
        RECT 1031.020 2.400 1031.160 59.170 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 386.140 518.350 386.200 ;
        RECT 521.710 386.140 522.030 386.200 ;
        RECT 518.030 386.000 522.030 386.140 ;
        RECT 518.030 385.940 518.350 386.000 ;
        RECT 521.710 385.940 522.030 386.000 ;
        RECT 518.030 59.060 518.350 59.120 ;
        RECT 1048.870 59.060 1049.190 59.120 ;
        RECT 518.030 58.920 1049.190 59.060 ;
        RECT 518.030 58.860 518.350 58.920 ;
        RECT 1048.870 58.860 1049.190 58.920 ;
      LAYER via ;
        RECT 518.060 385.940 518.320 386.200 ;
        RECT 521.740 385.940 522.000 386.200 ;
        RECT 518.060 58.860 518.320 59.120 ;
        RECT 1048.900 58.860 1049.160 59.120 ;
      LAYER met2 ;
        RECT 523.010 400.250 523.290 404.000 ;
        RECT 521.800 400.110 523.290 400.250 ;
        RECT 521.800 386.230 521.940 400.110 ;
        RECT 523.010 400.000 523.290 400.110 ;
        RECT 518.060 385.910 518.320 386.230 ;
        RECT 521.740 385.910 522.000 386.230 ;
        RECT 518.120 59.150 518.260 385.910 ;
        RECT 518.060 58.830 518.320 59.150 ;
        RECT 1048.900 58.830 1049.160 59.150 ;
        RECT 1048.960 2.400 1049.100 58.830 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 58.720 525.250 58.780 ;
        RECT 1066.810 58.720 1067.130 58.780 ;
        RECT 524.930 58.580 1067.130 58.720 ;
        RECT 524.930 58.520 525.250 58.580 ;
        RECT 1066.810 58.520 1067.130 58.580 ;
      LAYER via ;
        RECT 524.960 58.520 525.220 58.780 ;
        RECT 1066.840 58.520 1067.100 58.780 ;
      LAYER met2 ;
        RECT 528.530 400.250 528.810 404.000 ;
        RECT 527.320 400.110 528.810 400.250 ;
        RECT 527.320 387.330 527.460 400.110 ;
        RECT 528.530 400.000 528.810 400.110 ;
        RECT 525.020 387.190 527.460 387.330 ;
        RECT 525.020 58.810 525.160 387.190 ;
        RECT 524.960 58.490 525.220 58.810 ;
        RECT 1066.840 58.490 1067.100 58.810 ;
        RECT 1066.900 2.400 1067.040 58.490 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 56.680 532.150 56.740 ;
        RECT 1084.290 56.680 1084.610 56.740 ;
        RECT 531.830 56.540 1084.610 56.680 ;
        RECT 531.830 56.480 532.150 56.540 ;
        RECT 1084.290 56.480 1084.610 56.540 ;
      LAYER via ;
        RECT 531.860 56.480 532.120 56.740 ;
        RECT 1084.320 56.480 1084.580 56.740 ;
      LAYER met2 ;
        RECT 533.590 400.250 533.870 404.000 ;
        RECT 532.840 400.110 533.870 400.250 ;
        RECT 532.840 386.650 532.980 400.110 ;
        RECT 533.590 400.000 533.870 400.110 ;
        RECT 531.920 386.510 532.980 386.650 ;
        RECT 531.920 56.770 532.060 386.510 ;
        RECT 531.860 56.450 532.120 56.770 ;
        RECT 1084.320 56.450 1084.580 56.770 ;
        RECT 1084.380 2.400 1084.520 56.450 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 77.760 538.590 77.820 ;
        RECT 1099.930 77.760 1100.250 77.820 ;
        RECT 538.270 77.620 1100.250 77.760 ;
        RECT 538.270 77.560 538.590 77.620 ;
        RECT 1099.930 77.560 1100.250 77.620 ;
      LAYER via ;
        RECT 538.300 77.560 538.560 77.820 ;
        RECT 1099.960 77.560 1100.220 77.820 ;
      LAYER met2 ;
        RECT 539.110 400.250 539.390 404.000 ;
        RECT 538.360 400.110 539.390 400.250 ;
        RECT 538.360 77.850 538.500 400.110 ;
        RECT 539.110 400.000 539.390 400.110 ;
        RECT 538.300 77.530 538.560 77.850 ;
        RECT 1099.960 77.530 1100.220 77.850 ;
        RECT 1100.020 1.770 1100.160 77.530 ;
        RECT 1102.110 1.770 1102.670 2.400 ;
        RECT 1100.020 1.630 1102.670 1.770 ;
        RECT 1102.110 -4.800 1102.670 1.630 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 386.480 539.050 386.540 ;
        RECT 543.330 386.480 543.650 386.540 ;
        RECT 538.730 386.340 543.650 386.480 ;
        RECT 538.730 386.280 539.050 386.340 ;
        RECT 543.330 386.280 543.650 386.340 ;
        RECT 538.730 84.560 539.050 84.620 ;
        RECT 1117.870 84.560 1118.190 84.620 ;
        RECT 538.730 84.420 1118.190 84.560 ;
        RECT 538.730 84.360 539.050 84.420 ;
        RECT 1117.870 84.360 1118.190 84.420 ;
      LAYER via ;
        RECT 538.760 386.280 539.020 386.540 ;
        RECT 543.360 386.280 543.620 386.540 ;
        RECT 538.760 84.360 539.020 84.620 ;
        RECT 1117.900 84.360 1118.160 84.620 ;
      LAYER met2 ;
        RECT 544.630 400.250 544.910 404.000 ;
        RECT 543.420 400.110 544.910 400.250 ;
        RECT 543.420 386.570 543.560 400.110 ;
        RECT 544.630 400.000 544.910 400.110 ;
        RECT 538.760 386.250 539.020 386.570 ;
        RECT 543.360 386.250 543.620 386.570 ;
        RECT 538.820 84.650 538.960 386.250 ;
        RECT 538.760 84.330 539.020 84.650 ;
        RECT 1117.900 84.330 1118.160 84.650 ;
        RECT 1117.960 1.770 1118.100 84.330 ;
        RECT 1119.590 1.770 1120.150 2.400 ;
        RECT 1117.960 1.630 1120.150 1.770 ;
        RECT 1119.590 -4.800 1120.150 1.630 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 376.280 545.490 376.340 ;
        RECT 548.850 376.280 549.170 376.340 ;
        RECT 545.170 376.140 549.170 376.280 ;
        RECT 545.170 376.080 545.490 376.140 ;
        RECT 548.850 376.080 549.170 376.140 ;
        RECT 545.170 91.360 545.490 91.420 ;
        RECT 1132.130 91.360 1132.450 91.420 ;
        RECT 545.170 91.220 1132.450 91.360 ;
        RECT 545.170 91.160 545.490 91.220 ;
        RECT 1132.130 91.160 1132.450 91.220 ;
      LAYER via ;
        RECT 545.200 376.080 545.460 376.340 ;
        RECT 548.880 376.080 549.140 376.340 ;
        RECT 545.200 91.160 545.460 91.420 ;
        RECT 1132.160 91.160 1132.420 91.420 ;
      LAYER met2 ;
        RECT 550.150 400.250 550.430 404.000 ;
        RECT 548.940 400.110 550.430 400.250 ;
        RECT 548.940 376.370 549.080 400.110 ;
        RECT 550.150 400.000 550.430 400.110 ;
        RECT 545.200 376.050 545.460 376.370 ;
        RECT 548.880 376.050 549.140 376.370 ;
        RECT 545.260 91.450 545.400 376.050 ;
        RECT 545.200 91.130 545.460 91.450 ;
        RECT 1132.160 91.130 1132.420 91.450 ;
        RECT 1132.220 82.870 1132.360 91.130 ;
        RECT 1132.220 82.730 1137.880 82.870 ;
        RECT 1137.740 2.400 1137.880 82.730 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.990 375.940 553.310 376.000 ;
        RECT 554.370 375.940 554.690 376.000 ;
        RECT 552.990 375.800 554.690 375.940 ;
        RECT 552.990 375.740 553.310 375.800 ;
        RECT 554.370 375.740 554.690 375.800 ;
        RECT 552.990 91.700 553.310 91.760 ;
        RECT 1152.370 91.700 1152.690 91.760 ;
        RECT 552.990 91.560 1152.690 91.700 ;
        RECT 552.990 91.500 553.310 91.560 ;
        RECT 1152.370 91.500 1152.690 91.560 ;
      LAYER via ;
        RECT 553.020 375.740 553.280 376.000 ;
        RECT 554.400 375.740 554.660 376.000 ;
        RECT 553.020 91.500 553.280 91.760 ;
        RECT 1152.400 91.500 1152.660 91.760 ;
      LAYER met2 ;
        RECT 555.670 400.250 555.950 404.000 ;
        RECT 554.460 400.110 555.950 400.250 ;
        RECT 554.460 376.030 554.600 400.110 ;
        RECT 555.670 400.000 555.950 400.110 ;
        RECT 553.020 375.710 553.280 376.030 ;
        RECT 554.400 375.710 554.660 376.030 ;
        RECT 553.080 91.790 553.220 375.710 ;
        RECT 553.020 91.470 553.280 91.790 ;
        RECT 1152.400 91.470 1152.660 91.790 ;
        RECT 1152.460 82.870 1152.600 91.470 ;
        RECT 1152.460 82.730 1155.360 82.870 ;
        RECT 1155.220 2.400 1155.360 82.730 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.090 39.340 408.410 39.400 ;
        RECT 676.270 39.340 676.590 39.400 ;
        RECT 408.090 39.200 676.590 39.340 ;
        RECT 408.090 39.140 408.410 39.200 ;
        RECT 676.270 39.140 676.590 39.200 ;
      LAYER via ;
        RECT 408.120 39.140 408.380 39.400 ;
        RECT 676.300 39.140 676.560 39.400 ;
      LAYER met2 ;
        RECT 408.010 400.180 408.290 404.000 ;
        RECT 408.010 400.000 408.320 400.180 ;
        RECT 408.180 39.430 408.320 400.000 ;
        RECT 408.120 39.110 408.380 39.430 ;
        RECT 676.300 39.110 676.560 39.430 ;
        RECT 676.360 2.400 676.500 39.110 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 376.620 559.750 376.680 ;
        RECT 560.810 376.620 561.130 376.680 ;
        RECT 559.430 376.480 561.130 376.620 ;
        RECT 559.430 376.420 559.750 376.480 ;
        RECT 560.810 376.420 561.130 376.480 ;
        RECT 559.430 92.040 559.750 92.100 ;
        RECT 1173.070 92.040 1173.390 92.100 ;
        RECT 559.430 91.900 1173.390 92.040 ;
        RECT 559.430 91.840 559.750 91.900 ;
        RECT 1173.070 91.840 1173.390 91.900 ;
      LAYER via ;
        RECT 559.460 376.420 559.720 376.680 ;
        RECT 560.840 376.420 561.100 376.680 ;
        RECT 559.460 91.840 559.720 92.100 ;
        RECT 1173.100 91.840 1173.360 92.100 ;
      LAYER met2 ;
        RECT 561.190 400.250 561.470 404.000 ;
        RECT 560.900 400.110 561.470 400.250 ;
        RECT 560.900 376.710 561.040 400.110 ;
        RECT 561.190 400.000 561.470 400.110 ;
        RECT 559.460 376.390 559.720 376.710 ;
        RECT 560.840 376.390 561.100 376.710 ;
        RECT 559.520 92.130 559.660 376.390 ;
        RECT 559.460 91.810 559.720 92.130 ;
        RECT 1173.100 91.810 1173.360 92.130 ;
        RECT 1173.160 2.400 1173.300 91.810 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 92.380 567.110 92.440 ;
        RECT 1186.870 92.380 1187.190 92.440 ;
        RECT 566.790 92.240 1187.190 92.380 ;
        RECT 566.790 92.180 567.110 92.240 ;
        RECT 1186.870 92.180 1187.190 92.240 ;
      LAYER via ;
        RECT 566.820 92.180 567.080 92.440 ;
        RECT 1186.900 92.180 1187.160 92.440 ;
      LAYER met2 ;
        RECT 566.710 400.180 566.990 404.000 ;
        RECT 566.710 400.000 567.020 400.180 ;
        RECT 566.880 92.470 567.020 400.000 ;
        RECT 566.820 92.150 567.080 92.470 ;
        RECT 1186.900 92.150 1187.160 92.470 ;
        RECT 1186.960 82.870 1187.100 92.150 ;
        RECT 1186.960 82.730 1188.480 82.870 ;
        RECT 1188.340 1.770 1188.480 82.730 ;
        RECT 1190.430 1.770 1190.990 2.400 ;
        RECT 1188.340 1.630 1190.990 1.770 ;
        RECT 1190.430 -4.800 1190.990 1.630 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.250 92.720 567.570 92.780 ;
        RECT 1207.570 92.720 1207.890 92.780 ;
        RECT 567.250 92.580 1207.890 92.720 ;
        RECT 567.250 92.520 567.570 92.580 ;
        RECT 1207.570 92.520 1207.890 92.580 ;
      LAYER via ;
        RECT 567.280 92.520 567.540 92.780 ;
        RECT 1207.600 92.520 1207.860 92.780 ;
      LAYER met2 ;
        RECT 572.230 400.250 572.510 404.000 ;
        RECT 571.020 400.110 572.510 400.250 ;
        RECT 571.020 324.370 571.160 400.110 ;
        RECT 572.230 400.000 572.510 400.110 ;
        RECT 567.340 324.230 571.160 324.370 ;
        RECT 567.340 92.810 567.480 324.230 ;
        RECT 567.280 92.490 567.540 92.810 ;
        RECT 1207.600 92.490 1207.860 92.810 ;
        RECT 1207.660 82.870 1207.800 92.490 ;
        RECT 1207.660 82.730 1208.720 82.870 ;
        RECT 1208.580 2.400 1208.720 82.730 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.690 96.460 574.010 96.520 ;
        RECT 1221.370 96.460 1221.690 96.520 ;
        RECT 573.690 96.320 1221.690 96.460 ;
        RECT 573.690 96.260 574.010 96.320 ;
        RECT 1221.370 96.260 1221.690 96.320 ;
      LAYER via ;
        RECT 573.720 96.260 573.980 96.520 ;
        RECT 1221.400 96.260 1221.660 96.520 ;
      LAYER met2 ;
        RECT 577.750 400.250 578.030 404.000 ;
        RECT 576.540 400.110 578.030 400.250 ;
        RECT 576.540 324.370 576.680 400.110 ;
        RECT 577.750 400.000 578.030 400.110 ;
        RECT 573.780 324.230 576.680 324.370 ;
        RECT 573.780 96.550 573.920 324.230 ;
        RECT 573.720 96.230 573.980 96.550 ;
        RECT 1221.400 96.230 1221.660 96.550 ;
        RECT 1221.460 82.870 1221.600 96.230 ;
        RECT 1221.460 82.730 1226.200 82.870 ;
        RECT 1226.060 2.400 1226.200 82.730 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.050 96.120 581.370 96.180 ;
        RECT 1242.070 96.120 1242.390 96.180 ;
        RECT 581.050 95.980 1242.390 96.120 ;
        RECT 581.050 95.920 581.370 95.980 ;
        RECT 1242.070 95.920 1242.390 95.980 ;
      LAYER via ;
        RECT 581.080 95.920 581.340 96.180 ;
        RECT 1242.100 95.920 1242.360 96.180 ;
      LAYER met2 ;
        RECT 582.810 400.250 583.090 404.000 ;
        RECT 581.600 400.110 583.090 400.250 ;
        RECT 581.600 324.370 581.740 400.110 ;
        RECT 582.810 400.000 583.090 400.110 ;
        RECT 581.140 324.230 581.740 324.370 ;
        RECT 581.140 96.210 581.280 324.230 ;
        RECT 581.080 95.890 581.340 96.210 ;
        RECT 1242.100 95.890 1242.360 96.210 ;
        RECT 1242.160 1.770 1242.300 95.890 ;
        RECT 1243.790 1.770 1244.350 2.400 ;
        RECT 1242.160 1.630 1244.350 1.770 ;
        RECT 1243.790 -4.800 1244.350 1.630 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.950 95.780 588.270 95.840 ;
        RECT 1255.870 95.780 1256.190 95.840 ;
        RECT 587.950 95.640 1256.190 95.780 ;
        RECT 587.950 95.580 588.270 95.640 ;
        RECT 1255.870 95.580 1256.190 95.640 ;
        RECT 1255.870 20.980 1256.190 21.040 ;
        RECT 1261.850 20.980 1262.170 21.040 ;
        RECT 1255.870 20.840 1262.170 20.980 ;
        RECT 1255.870 20.780 1256.190 20.840 ;
        RECT 1261.850 20.780 1262.170 20.840 ;
      LAYER via ;
        RECT 587.980 95.580 588.240 95.840 ;
        RECT 1255.900 95.580 1256.160 95.840 ;
        RECT 1255.900 20.780 1256.160 21.040 ;
        RECT 1261.880 20.780 1262.140 21.040 ;
      LAYER met2 ;
        RECT 588.330 400.250 588.610 404.000 ;
        RECT 588.040 400.110 588.610 400.250 ;
        RECT 588.040 95.870 588.180 400.110 ;
        RECT 588.330 400.000 588.610 400.110 ;
        RECT 587.980 95.550 588.240 95.870 ;
        RECT 1255.900 95.550 1256.160 95.870 ;
        RECT 1255.960 21.070 1256.100 95.550 ;
        RECT 1255.900 20.750 1256.160 21.070 ;
        RECT 1261.880 20.750 1262.140 21.070 ;
        RECT 1261.940 2.400 1262.080 20.750 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 95.440 594.710 95.500 ;
        RECT 1276.570 95.440 1276.890 95.500 ;
        RECT 594.390 95.300 1276.890 95.440 ;
        RECT 594.390 95.240 594.710 95.300 ;
        RECT 1276.570 95.240 1276.890 95.300 ;
      LAYER via ;
        RECT 594.420 95.240 594.680 95.500 ;
        RECT 1276.600 95.240 1276.860 95.500 ;
      LAYER met2 ;
        RECT 593.850 400.180 594.130 404.000 ;
        RECT 593.850 400.000 594.160 400.180 ;
        RECT 594.020 386.650 594.160 400.000 ;
        RECT 594.020 386.510 594.620 386.650 ;
        RECT 594.480 95.530 594.620 386.510 ;
        RECT 594.420 95.210 594.680 95.530 ;
        RECT 1276.600 95.210 1276.860 95.530 ;
        RECT 1276.660 82.870 1276.800 95.210 ;
        RECT 1276.660 82.730 1279.560 82.870 ;
        RECT 1279.420 2.400 1279.560 82.730 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.850 386.140 595.170 386.200 ;
        RECT 598.070 386.140 598.390 386.200 ;
        RECT 594.850 386.000 598.390 386.140 ;
        RECT 594.850 385.940 595.170 386.000 ;
        RECT 598.070 385.940 598.390 386.000 ;
        RECT 594.850 95.100 595.170 95.160 ;
        RECT 1297.270 95.100 1297.590 95.160 ;
        RECT 594.850 94.960 1297.590 95.100 ;
        RECT 594.850 94.900 595.170 94.960 ;
        RECT 1297.270 94.900 1297.590 94.960 ;
      LAYER via ;
        RECT 594.880 385.940 595.140 386.200 ;
        RECT 598.100 385.940 598.360 386.200 ;
        RECT 594.880 94.900 595.140 95.160 ;
        RECT 1297.300 94.900 1297.560 95.160 ;
      LAYER met2 ;
        RECT 599.370 400.250 599.650 404.000 ;
        RECT 598.160 400.110 599.650 400.250 ;
        RECT 598.160 386.230 598.300 400.110 ;
        RECT 599.370 400.000 599.650 400.110 ;
        RECT 594.880 385.910 595.140 386.230 ;
        RECT 598.100 385.910 598.360 386.230 ;
        RECT 594.940 95.190 595.080 385.910 ;
        RECT 594.880 94.870 595.140 95.190 ;
        RECT 1297.300 94.870 1297.560 95.190 ;
        RECT 1297.360 2.400 1297.500 94.870 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 98.160 602.070 98.220 ;
        RECT 1311.070 98.160 1311.390 98.220 ;
        RECT 601.750 98.020 1311.390 98.160 ;
        RECT 601.750 97.960 602.070 98.020 ;
        RECT 1311.070 97.960 1311.390 98.020 ;
      LAYER via ;
        RECT 601.780 97.960 602.040 98.220 ;
        RECT 1311.100 97.960 1311.360 98.220 ;
      LAYER met2 ;
        RECT 604.890 400.250 605.170 404.000 ;
        RECT 603.680 400.110 605.170 400.250 ;
        RECT 603.680 324.370 603.820 400.110 ;
        RECT 604.890 400.000 605.170 400.110 ;
        RECT 601.840 324.230 603.820 324.370 ;
        RECT 601.840 98.250 601.980 324.230 ;
        RECT 601.780 97.930 602.040 98.250 ;
        RECT 1311.100 97.930 1311.360 98.250 ;
        RECT 1311.160 82.870 1311.300 97.930 ;
        RECT 1311.160 82.730 1312.680 82.870 ;
        RECT 1312.540 1.770 1312.680 82.730 ;
        RECT 1314.630 1.770 1315.190 2.400 ;
        RECT 1312.540 1.630 1315.190 1.770 ;
        RECT 1314.630 -4.800 1315.190 1.630 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 98.500 608.510 98.560 ;
        RECT 1331.770 98.500 1332.090 98.560 ;
        RECT 608.190 98.360 1332.090 98.500 ;
        RECT 608.190 98.300 608.510 98.360 ;
        RECT 1331.770 98.300 1332.090 98.360 ;
      LAYER via ;
        RECT 608.220 98.300 608.480 98.560 ;
        RECT 1331.800 98.300 1332.060 98.560 ;
      LAYER met2 ;
        RECT 610.410 400.250 610.690 404.000 ;
        RECT 609.200 400.110 610.690 400.250 ;
        RECT 609.200 324.370 609.340 400.110 ;
        RECT 610.410 400.000 610.690 400.110 ;
        RECT 608.280 324.230 609.340 324.370 ;
        RECT 608.280 98.590 608.420 324.230 ;
        RECT 608.220 98.270 608.480 98.590 ;
        RECT 1331.800 98.270 1332.060 98.590 ;
        RECT 1331.860 82.870 1332.000 98.270 ;
        RECT 1331.860 82.730 1332.920 82.870 ;
        RECT 1332.780 2.400 1332.920 82.730 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.550 38.320 408.870 38.380 ;
        RECT 694.210 38.320 694.530 38.380 ;
        RECT 408.550 38.180 694.530 38.320 ;
        RECT 408.550 38.120 408.870 38.180 ;
        RECT 694.210 38.120 694.530 38.180 ;
      LAYER via ;
        RECT 408.580 38.120 408.840 38.380 ;
        RECT 694.240 38.120 694.500 38.380 ;
      LAYER met2 ;
        RECT 413.530 400.250 413.810 404.000 ;
        RECT 412.320 400.110 413.810 400.250 ;
        RECT 412.320 398.210 412.460 400.110 ;
        RECT 413.530 400.000 413.810 400.110 ;
        RECT 410.020 398.070 412.460 398.210 ;
        RECT 410.020 351.970 410.160 398.070 ;
        RECT 408.640 351.830 410.160 351.970 ;
        RECT 408.640 38.410 408.780 351.830 ;
        RECT 408.580 38.090 408.840 38.410 ;
        RECT 694.240 38.090 694.500 38.410 ;
        RECT 694.300 2.400 694.440 38.090 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 98.840 615.410 98.900 ;
        RECT 1345.570 98.840 1345.890 98.900 ;
        RECT 615.090 98.700 1345.890 98.840 ;
        RECT 615.090 98.640 615.410 98.700 ;
        RECT 1345.570 98.640 1345.890 98.700 ;
      LAYER via ;
        RECT 615.120 98.640 615.380 98.900 ;
        RECT 1345.600 98.640 1345.860 98.900 ;
      LAYER met2 ;
        RECT 615.930 400.250 616.210 404.000 ;
        RECT 615.180 400.110 616.210 400.250 ;
        RECT 615.180 98.930 615.320 400.110 ;
        RECT 615.930 400.000 616.210 400.110 ;
        RECT 615.120 98.610 615.380 98.930 ;
        RECT 1345.600 98.610 1345.860 98.930 ;
        RECT 1345.660 82.870 1345.800 98.610 ;
        RECT 1345.660 82.730 1348.560 82.870 ;
        RECT 1348.420 17.410 1348.560 82.730 ;
        RECT 1348.420 17.270 1350.400 17.410 ;
        RECT 1350.260 2.400 1350.400 17.270 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.530 99.180 621.850 99.240 ;
        RECT 1366.270 99.180 1366.590 99.240 ;
        RECT 621.530 99.040 1366.590 99.180 ;
        RECT 621.530 98.980 621.850 99.040 ;
        RECT 1366.270 98.980 1366.590 99.040 ;
      LAYER via ;
        RECT 621.560 98.980 621.820 99.240 ;
        RECT 1366.300 98.980 1366.560 99.240 ;
      LAYER met2 ;
        RECT 621.450 400.180 621.730 404.000 ;
        RECT 621.450 400.000 621.760 400.180 ;
        RECT 621.620 99.270 621.760 400.000 ;
        RECT 621.560 98.950 621.820 99.270 ;
        RECT 1366.300 98.950 1366.560 99.270 ;
        RECT 1366.360 1.770 1366.500 98.950 ;
        RECT 1367.990 1.770 1368.550 2.400 ;
        RECT 1366.360 1.630 1368.550 1.770 ;
        RECT 1367.990 -4.800 1368.550 1.630 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 386.480 622.310 386.540 ;
        RECT 625.670 386.480 625.990 386.540 ;
        RECT 621.990 386.340 625.990 386.480 ;
        RECT 621.990 386.280 622.310 386.340 ;
        RECT 625.670 386.280 625.990 386.340 ;
        RECT 621.990 99.520 622.310 99.580 ;
        RECT 1380.070 99.520 1380.390 99.580 ;
        RECT 621.990 99.380 1380.390 99.520 ;
        RECT 621.990 99.320 622.310 99.380 ;
        RECT 1380.070 99.320 1380.390 99.380 ;
        RECT 1380.070 20.980 1380.390 21.040 ;
        RECT 1383.750 20.980 1384.070 21.040 ;
        RECT 1380.070 20.840 1384.070 20.980 ;
        RECT 1380.070 20.780 1380.390 20.840 ;
        RECT 1383.750 20.780 1384.070 20.840 ;
      LAYER via ;
        RECT 622.020 386.280 622.280 386.540 ;
        RECT 625.700 386.280 625.960 386.540 ;
        RECT 622.020 99.320 622.280 99.580 ;
        RECT 1380.100 99.320 1380.360 99.580 ;
        RECT 1380.100 20.780 1380.360 21.040 ;
        RECT 1383.780 20.780 1384.040 21.040 ;
      LAYER met2 ;
        RECT 626.970 400.250 627.250 404.000 ;
        RECT 625.760 400.110 627.250 400.250 ;
        RECT 625.760 386.570 625.900 400.110 ;
        RECT 626.970 400.000 627.250 400.110 ;
        RECT 622.020 386.250 622.280 386.570 ;
        RECT 625.700 386.250 625.960 386.570 ;
        RECT 622.080 99.610 622.220 386.250 ;
        RECT 622.020 99.290 622.280 99.610 ;
        RECT 1380.100 99.290 1380.360 99.610 ;
        RECT 1380.160 21.070 1380.300 99.290 ;
        RECT 1380.100 20.750 1380.360 21.070 ;
        RECT 1383.780 20.750 1384.040 21.070 ;
        RECT 1383.840 1.770 1383.980 20.750 ;
        RECT 1385.470 1.770 1386.030 2.400 ;
        RECT 1383.840 1.630 1386.030 1.770 ;
        RECT 1385.470 -4.800 1386.030 1.630 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.430 387.500 628.750 387.560 ;
        RECT 630.730 387.500 631.050 387.560 ;
        RECT 628.430 387.360 631.050 387.500 ;
        RECT 628.430 387.300 628.750 387.360 ;
        RECT 630.730 387.300 631.050 387.360 ;
        RECT 628.430 103.260 628.750 103.320 ;
        RECT 1400.770 103.260 1401.090 103.320 ;
        RECT 628.430 103.120 1401.090 103.260 ;
        RECT 628.430 103.060 628.750 103.120 ;
        RECT 1400.770 103.060 1401.090 103.120 ;
      LAYER via ;
        RECT 628.460 387.300 628.720 387.560 ;
        RECT 630.760 387.300 631.020 387.560 ;
        RECT 628.460 103.060 628.720 103.320 ;
        RECT 1400.800 103.060 1401.060 103.320 ;
      LAYER met2 ;
        RECT 632.030 400.250 632.310 404.000 ;
        RECT 630.820 400.110 632.310 400.250 ;
        RECT 630.820 387.590 630.960 400.110 ;
        RECT 632.030 400.000 632.310 400.110 ;
        RECT 628.460 387.270 628.720 387.590 ;
        RECT 630.760 387.270 631.020 387.590 ;
        RECT 628.520 103.350 628.660 387.270 ;
        RECT 628.460 103.030 628.720 103.350 ;
        RECT 1400.800 103.030 1401.060 103.350 ;
        RECT 1400.860 82.870 1401.000 103.030 ;
        RECT 1400.860 82.730 1403.760 82.870 ;
        RECT 1403.620 2.400 1403.760 82.730 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.790 102.920 636.110 102.980 ;
        RECT 1421.930 102.920 1422.250 102.980 ;
        RECT 635.790 102.780 1422.250 102.920 ;
        RECT 635.790 102.720 636.110 102.780 ;
        RECT 1421.930 102.720 1422.250 102.780 ;
      LAYER via ;
        RECT 635.820 102.720 636.080 102.980 ;
        RECT 1421.960 102.720 1422.220 102.980 ;
      LAYER met2 ;
        RECT 637.550 400.250 637.830 404.000 ;
        RECT 636.340 400.110 637.830 400.250 ;
        RECT 636.340 386.480 636.480 400.110 ;
        RECT 637.550 400.000 637.830 400.110 ;
        RECT 635.880 386.340 636.480 386.480 ;
        RECT 635.880 103.010 636.020 386.340 ;
        RECT 635.820 102.690 636.080 103.010 ;
        RECT 1421.960 102.690 1422.220 103.010 ;
        RECT 1422.020 17.410 1422.160 102.690 ;
        RECT 1421.560 17.270 1422.160 17.410 ;
        RECT 1421.560 2.400 1421.700 17.270 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.690 102.580 643.010 102.640 ;
        RECT 1435.270 102.580 1435.590 102.640 ;
        RECT 642.690 102.440 1435.590 102.580 ;
        RECT 642.690 102.380 643.010 102.440 ;
        RECT 1435.270 102.380 1435.590 102.440 ;
      LAYER via ;
        RECT 642.720 102.380 642.980 102.640 ;
        RECT 1435.300 102.380 1435.560 102.640 ;
      LAYER met2 ;
        RECT 643.070 400.250 643.350 404.000 ;
        RECT 642.780 400.110 643.350 400.250 ;
        RECT 642.780 102.670 642.920 400.110 ;
        RECT 643.070 400.000 643.350 400.110 ;
        RECT 642.720 102.350 642.980 102.670 ;
        RECT 1435.300 102.350 1435.560 102.670 ;
        RECT 1435.360 82.870 1435.500 102.350 ;
        RECT 1435.360 82.730 1436.880 82.870 ;
        RECT 1436.740 1.770 1436.880 82.730 ;
        RECT 1438.830 1.770 1439.390 2.400 ;
        RECT 1436.740 1.630 1439.390 1.770 ;
        RECT 1438.830 -4.800 1439.390 1.630 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.590 387.640 649.910 387.900 ;
        RECT 649.680 386.200 649.820 387.640 ;
        RECT 649.590 385.940 649.910 386.200 ;
        RECT 649.590 102.240 649.910 102.300 ;
        RECT 1455.970 102.240 1456.290 102.300 ;
        RECT 649.590 102.100 1456.290 102.240 ;
        RECT 649.590 102.040 649.910 102.100 ;
        RECT 1455.970 102.040 1456.290 102.100 ;
      LAYER via ;
        RECT 649.620 387.640 649.880 387.900 ;
        RECT 649.620 385.940 649.880 386.200 ;
        RECT 649.620 102.040 649.880 102.300 ;
        RECT 1456.000 102.040 1456.260 102.300 ;
      LAYER met2 ;
        RECT 648.590 400.250 648.870 404.000 ;
        RECT 648.590 400.110 649.820 400.250 ;
        RECT 648.590 400.000 648.870 400.110 ;
        RECT 649.680 387.930 649.820 400.110 ;
        RECT 649.620 387.610 649.880 387.930 ;
        RECT 649.620 385.910 649.880 386.230 ;
        RECT 649.680 102.330 649.820 385.910 ;
        RECT 649.620 102.010 649.880 102.330 ;
        RECT 1456.000 102.010 1456.260 102.330 ;
        RECT 1456.060 82.870 1456.200 102.010 ;
        RECT 1456.060 82.730 1457.120 82.870 ;
        RECT 1456.980 2.400 1457.120 82.730 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.050 101.900 650.370 101.960 ;
        RECT 1469.770 101.900 1470.090 101.960 ;
        RECT 650.050 101.760 1470.090 101.900 ;
        RECT 650.050 101.700 650.370 101.760 ;
        RECT 1469.770 101.700 1470.090 101.760 ;
      LAYER via ;
        RECT 650.080 101.700 650.340 101.960 ;
        RECT 1469.800 101.700 1470.060 101.960 ;
      LAYER met2 ;
        RECT 654.110 400.250 654.390 404.000 ;
        RECT 652.900 400.110 654.390 400.250 ;
        RECT 652.900 324.370 653.040 400.110 ;
        RECT 654.110 400.000 654.390 400.110 ;
        RECT 650.140 324.230 653.040 324.370 ;
        RECT 650.140 101.990 650.280 324.230 ;
        RECT 650.080 101.670 650.340 101.990 ;
        RECT 1469.800 101.670 1470.060 101.990 ;
        RECT 1469.860 82.870 1470.000 101.670 ;
        RECT 1469.860 82.730 1474.600 82.870 ;
        RECT 1474.460 2.400 1474.600 82.730 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.950 101.560 657.270 101.620 ;
        RECT 1490.470 101.560 1490.790 101.620 ;
        RECT 656.950 101.420 1490.790 101.560 ;
        RECT 656.950 101.360 657.270 101.420 ;
        RECT 1490.470 101.360 1490.790 101.420 ;
      LAYER via ;
        RECT 656.980 101.360 657.240 101.620 ;
        RECT 1490.500 101.360 1490.760 101.620 ;
      LAYER met2 ;
        RECT 659.630 400.250 659.910 404.000 ;
        RECT 658.420 400.110 659.910 400.250 ;
        RECT 658.420 324.370 658.560 400.110 ;
        RECT 659.630 400.000 659.910 400.110 ;
        RECT 657.040 324.230 658.560 324.370 ;
        RECT 657.040 101.650 657.180 324.230 ;
        RECT 656.980 101.330 657.240 101.650 ;
        RECT 1490.500 101.330 1490.760 101.650 ;
        RECT 1490.560 1.770 1490.700 101.330 ;
        RECT 1492.190 1.770 1492.750 2.400 ;
        RECT 1490.560 1.630 1492.750 1.770 ;
        RECT 1492.190 -4.800 1492.750 1.630 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.930 386.480 663.250 386.540 ;
        RECT 664.310 386.480 664.630 386.540 ;
        RECT 662.930 386.340 664.630 386.480 ;
        RECT 662.930 386.280 663.250 386.340 ;
        RECT 664.310 386.280 664.630 386.340 ;
        RECT 662.930 101.220 663.250 101.280 ;
        RECT 1504.270 101.220 1504.590 101.280 ;
        RECT 662.930 101.080 1504.590 101.220 ;
        RECT 662.930 101.020 663.250 101.080 ;
        RECT 1504.270 101.020 1504.590 101.080 ;
      LAYER via ;
        RECT 662.960 386.280 663.220 386.540 ;
        RECT 664.340 386.280 664.600 386.540 ;
        RECT 662.960 101.020 663.220 101.280 ;
        RECT 1504.300 101.020 1504.560 101.280 ;
      LAYER met2 ;
        RECT 665.150 400.250 665.430 404.000 ;
        RECT 664.400 400.110 665.430 400.250 ;
        RECT 664.400 386.570 664.540 400.110 ;
        RECT 665.150 400.000 665.430 400.110 ;
        RECT 662.960 386.250 663.220 386.570 ;
        RECT 664.340 386.250 664.600 386.570 ;
        RECT 663.020 101.310 663.160 386.250 ;
        RECT 662.960 100.990 663.220 101.310 ;
        RECT 1504.300 100.990 1504.560 101.310 ;
        RECT 1504.360 82.870 1504.500 100.990 ;
        RECT 1504.360 82.730 1507.720 82.870 ;
        RECT 1507.580 1.770 1507.720 82.730 ;
        RECT 1509.670 1.770 1510.230 2.400 ;
        RECT 1507.580 1.630 1510.230 1.770 ;
        RECT 1509.670 -4.800 1510.230 1.630 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.530 376.280 414.850 376.340 ;
        RECT 417.750 376.280 418.070 376.340 ;
        RECT 414.530 376.140 418.070 376.280 ;
        RECT 414.530 376.080 414.850 376.140 ;
        RECT 417.750 376.080 418.070 376.140 ;
        RECT 414.530 32.540 414.850 32.600 ;
        RECT 553.450 32.540 553.770 32.600 ;
        RECT 414.530 32.400 553.770 32.540 ;
        RECT 414.530 32.340 414.850 32.400 ;
        RECT 553.450 32.340 553.770 32.400 ;
        RECT 553.450 16.220 553.770 16.280 ;
        RECT 712.150 16.220 712.470 16.280 ;
        RECT 553.450 16.080 712.470 16.220 ;
        RECT 553.450 16.020 553.770 16.080 ;
        RECT 712.150 16.020 712.470 16.080 ;
      LAYER via ;
        RECT 414.560 376.080 414.820 376.340 ;
        RECT 417.780 376.080 418.040 376.340 ;
        RECT 414.560 32.340 414.820 32.600 ;
        RECT 553.480 32.340 553.740 32.600 ;
        RECT 553.480 16.020 553.740 16.280 ;
        RECT 712.180 16.020 712.440 16.280 ;
      LAYER met2 ;
        RECT 419.050 400.250 419.330 404.000 ;
        RECT 417.840 400.110 419.330 400.250 ;
        RECT 417.840 376.370 417.980 400.110 ;
        RECT 419.050 400.000 419.330 400.110 ;
        RECT 414.560 376.050 414.820 376.370 ;
        RECT 417.780 376.050 418.040 376.370 ;
        RECT 414.620 32.630 414.760 376.050 ;
        RECT 414.560 32.310 414.820 32.630 ;
        RECT 553.480 32.310 553.740 32.630 ;
        RECT 553.540 16.310 553.680 32.310 ;
        RECT 553.480 15.990 553.740 16.310 ;
        RECT 712.180 15.990 712.440 16.310 ;
        RECT 712.240 2.400 712.380 15.990 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.830 388.320 670.150 388.580 ;
        RECT 669.920 387.220 670.060 388.320 ;
        RECT 669.830 386.960 670.150 387.220 ;
        RECT 669.830 100.880 670.150 100.940 ;
        RECT 1524.970 100.880 1525.290 100.940 ;
        RECT 669.830 100.740 1525.290 100.880 ;
        RECT 669.830 100.680 670.150 100.740 ;
        RECT 1524.970 100.680 1525.290 100.740 ;
      LAYER via ;
        RECT 669.860 388.320 670.120 388.580 ;
        RECT 669.860 386.960 670.120 387.220 ;
        RECT 669.860 100.680 670.120 100.940 ;
        RECT 1525.000 100.680 1525.260 100.940 ;
      LAYER met2 ;
        RECT 670.670 400.250 670.950 404.000 ;
        RECT 669.920 400.110 670.950 400.250 ;
        RECT 669.920 388.610 670.060 400.110 ;
        RECT 670.670 400.000 670.950 400.110 ;
        RECT 669.860 388.290 670.120 388.610 ;
        RECT 669.860 386.930 670.120 387.250 ;
        RECT 669.920 100.970 670.060 386.930 ;
        RECT 669.860 100.650 670.120 100.970 ;
        RECT 1525.000 100.650 1525.260 100.970 ;
        RECT 1525.060 82.870 1525.200 100.650 ;
        RECT 1525.060 82.730 1527.960 82.870 ;
        RECT 1527.820 2.400 1527.960 82.730 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.290 386.480 670.610 386.540 ;
        RECT 674.890 386.480 675.210 386.540 ;
        RECT 670.290 386.340 675.210 386.480 ;
        RECT 670.290 386.280 670.610 386.340 ;
        RECT 674.890 386.280 675.210 386.340 ;
        RECT 670.290 100.540 670.610 100.600 ;
        RECT 1539.230 100.540 1539.550 100.600 ;
        RECT 670.290 100.400 1539.550 100.540 ;
        RECT 670.290 100.340 670.610 100.400 ;
        RECT 1539.230 100.340 1539.550 100.400 ;
        RECT 1539.230 20.980 1539.550 21.040 ;
        RECT 1545.210 20.980 1545.530 21.040 ;
        RECT 1539.230 20.840 1545.530 20.980 ;
        RECT 1539.230 20.780 1539.550 20.840 ;
        RECT 1545.210 20.780 1545.530 20.840 ;
      LAYER via ;
        RECT 670.320 386.280 670.580 386.540 ;
        RECT 674.920 386.280 675.180 386.540 ;
        RECT 670.320 100.340 670.580 100.600 ;
        RECT 1539.260 100.340 1539.520 100.600 ;
        RECT 1539.260 20.780 1539.520 21.040 ;
        RECT 1545.240 20.780 1545.500 21.040 ;
      LAYER met2 ;
        RECT 675.730 400.250 676.010 404.000 ;
        RECT 674.980 400.110 676.010 400.250 ;
        RECT 674.980 386.570 675.120 400.110 ;
        RECT 675.730 400.000 676.010 400.110 ;
        RECT 670.320 386.250 670.580 386.570 ;
        RECT 674.920 386.250 675.180 386.570 ;
        RECT 670.380 100.630 670.520 386.250 ;
        RECT 670.320 100.310 670.580 100.630 ;
        RECT 1539.260 100.310 1539.520 100.630 ;
        RECT 1539.320 21.070 1539.460 100.310 ;
        RECT 1539.260 20.750 1539.520 21.070 ;
        RECT 1545.240 20.750 1545.500 21.070 ;
        RECT 1545.300 2.400 1545.440 20.750 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.730 386.480 677.050 386.540 ;
        RECT 679.950 386.480 680.270 386.540 ;
        RECT 676.730 386.340 680.270 386.480 ;
        RECT 676.730 386.280 677.050 386.340 ;
        RECT 679.950 386.280 680.270 386.340 ;
        RECT 676.730 100.200 677.050 100.260 ;
        RECT 1559.470 100.200 1559.790 100.260 ;
        RECT 676.730 100.060 1559.790 100.200 ;
        RECT 676.730 100.000 677.050 100.060 ;
        RECT 1559.470 100.000 1559.790 100.060 ;
      LAYER via ;
        RECT 676.760 386.280 677.020 386.540 ;
        RECT 679.980 386.280 680.240 386.540 ;
        RECT 676.760 100.000 677.020 100.260 ;
        RECT 1559.500 100.000 1559.760 100.260 ;
      LAYER met2 ;
        RECT 681.250 400.250 681.530 404.000 ;
        RECT 680.040 400.110 681.530 400.250 ;
        RECT 680.040 386.570 680.180 400.110 ;
        RECT 681.250 400.000 681.530 400.110 ;
        RECT 676.760 386.250 677.020 386.570 ;
        RECT 679.980 386.250 680.240 386.570 ;
        RECT 676.820 100.290 676.960 386.250 ;
        RECT 676.760 99.970 677.020 100.290 ;
        RECT 1559.500 99.970 1559.760 100.290 ;
        RECT 1559.560 82.870 1559.700 99.970 ;
        RECT 1559.560 82.730 1561.080 82.870 ;
        RECT 1560.940 1.770 1561.080 82.730 ;
        RECT 1563.030 1.770 1563.590 2.400 ;
        RECT 1560.940 1.630 1563.590 1.770 ;
        RECT 1563.030 -4.800 1563.590 1.630 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.550 119.580 684.870 119.640 ;
        RECT 1580.170 119.580 1580.490 119.640 ;
        RECT 684.550 119.440 1580.490 119.580 ;
        RECT 684.550 119.380 684.870 119.440 ;
        RECT 1580.170 119.380 1580.490 119.440 ;
      LAYER via ;
        RECT 684.580 119.380 684.840 119.640 ;
        RECT 1580.200 119.380 1580.460 119.640 ;
      LAYER met2 ;
        RECT 686.770 400.250 687.050 404.000 ;
        RECT 685.560 400.110 687.050 400.250 ;
        RECT 685.560 324.370 685.700 400.110 ;
        RECT 686.770 400.000 687.050 400.110 ;
        RECT 684.640 324.230 685.700 324.370 ;
        RECT 684.640 119.670 684.780 324.230 ;
        RECT 684.580 119.350 684.840 119.670 ;
        RECT 1580.200 119.350 1580.460 119.670 ;
        RECT 1580.260 82.870 1580.400 119.350 ;
        RECT 1580.260 82.730 1581.320 82.870 ;
        RECT 1581.180 2.400 1581.320 82.730 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 691.450 119.920 691.770 119.980 ;
        RECT 1593.970 119.920 1594.290 119.980 ;
        RECT 691.450 119.780 1594.290 119.920 ;
        RECT 691.450 119.720 691.770 119.780 ;
        RECT 1593.970 119.720 1594.290 119.780 ;
      LAYER via ;
        RECT 691.480 119.720 691.740 119.980 ;
        RECT 1594.000 119.720 1594.260 119.980 ;
      LAYER met2 ;
        RECT 692.290 400.250 692.570 404.000 ;
        RECT 691.540 400.110 692.570 400.250 ;
        RECT 691.540 120.010 691.680 400.110 ;
        RECT 692.290 400.000 692.570 400.110 ;
        RECT 691.480 119.690 691.740 120.010 ;
        RECT 1594.000 119.690 1594.260 120.010 ;
        RECT 1594.060 82.870 1594.200 119.690 ;
        RECT 1594.060 82.730 1598.800 82.870 ;
        RECT 1598.660 2.400 1598.800 82.730 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 698.350 126.040 698.670 126.100 ;
        RECT 1614.670 126.040 1614.990 126.100 ;
        RECT 698.350 125.900 1614.990 126.040 ;
        RECT 698.350 125.840 698.670 125.900 ;
        RECT 1614.670 125.840 1614.990 125.900 ;
      LAYER via ;
        RECT 698.380 125.840 698.640 126.100 ;
        RECT 1614.700 125.840 1614.960 126.100 ;
      LAYER met2 ;
        RECT 697.810 400.250 698.090 404.000 ;
        RECT 697.810 400.110 699.500 400.250 ;
        RECT 697.810 400.000 698.090 400.110 ;
        RECT 699.360 324.370 699.500 400.110 ;
        RECT 698.440 324.230 699.500 324.370 ;
        RECT 698.440 126.130 698.580 324.230 ;
        RECT 698.380 125.810 698.640 126.130 ;
        RECT 1614.700 125.810 1614.960 126.130 ;
        RECT 1614.760 1.770 1614.900 125.810 ;
        RECT 1616.390 1.770 1616.950 2.400 ;
        RECT 1614.760 1.630 1616.950 1.770 ;
        RECT 1616.390 -4.800 1616.950 1.630 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.890 376.620 698.210 376.680 ;
        RECT 702.030 376.620 702.350 376.680 ;
        RECT 697.890 376.480 702.350 376.620 ;
        RECT 697.890 376.420 698.210 376.480 ;
        RECT 702.030 376.420 702.350 376.480 ;
        RECT 697.890 126.380 698.210 126.440 ;
        RECT 1628.470 126.380 1628.790 126.440 ;
        RECT 697.890 126.240 1628.790 126.380 ;
        RECT 697.890 126.180 698.210 126.240 ;
        RECT 1628.470 126.180 1628.790 126.240 ;
      LAYER via ;
        RECT 697.920 376.420 698.180 376.680 ;
        RECT 702.060 376.420 702.320 376.680 ;
        RECT 697.920 126.180 698.180 126.440 ;
        RECT 1628.500 126.180 1628.760 126.440 ;
      LAYER met2 ;
        RECT 703.330 400.250 703.610 404.000 ;
        RECT 702.120 400.110 703.610 400.250 ;
        RECT 702.120 376.710 702.260 400.110 ;
        RECT 703.330 400.000 703.610 400.110 ;
        RECT 697.920 376.390 698.180 376.710 ;
        RECT 702.060 376.390 702.320 376.710 ;
        RECT 697.980 126.470 698.120 376.390 ;
        RECT 697.920 126.150 698.180 126.470 ;
        RECT 1628.500 126.150 1628.760 126.470 ;
        RECT 1628.560 82.870 1628.700 126.150 ;
        RECT 1628.560 82.730 1631.920 82.870 ;
        RECT 1631.780 1.770 1631.920 82.730 ;
        RECT 1633.870 1.770 1634.430 2.400 ;
        RECT 1631.780 1.630 1634.430 1.770 ;
        RECT 1633.870 -4.800 1634.430 1.630 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.790 126.720 705.110 126.780 ;
        RECT 1649.170 126.720 1649.490 126.780 ;
        RECT 704.790 126.580 1649.490 126.720 ;
        RECT 704.790 126.520 705.110 126.580 ;
        RECT 1649.170 126.520 1649.490 126.580 ;
      LAYER via ;
        RECT 704.820 126.520 705.080 126.780 ;
        RECT 1649.200 126.520 1649.460 126.780 ;
      LAYER met2 ;
        RECT 708.850 400.250 709.130 404.000 ;
        RECT 707.640 400.110 709.130 400.250 ;
        RECT 707.640 351.970 707.780 400.110 ;
        RECT 708.850 400.000 709.130 400.110 ;
        RECT 704.880 351.830 707.780 351.970 ;
        RECT 704.880 126.810 705.020 351.830 ;
        RECT 704.820 126.490 705.080 126.810 ;
        RECT 1649.200 126.490 1649.460 126.810 ;
        RECT 1649.260 82.870 1649.400 126.490 ;
        RECT 1649.260 82.730 1652.160 82.870 ;
        RECT 1652.020 2.400 1652.160 82.730 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 712.150 127.060 712.470 127.120 ;
        RECT 1662.970 127.060 1663.290 127.120 ;
        RECT 712.150 126.920 1663.290 127.060 ;
        RECT 712.150 126.860 712.470 126.920 ;
        RECT 1662.970 126.860 1663.290 126.920 ;
        RECT 1662.970 15.200 1663.290 15.260 ;
        RECT 1669.410 15.200 1669.730 15.260 ;
        RECT 1662.970 15.060 1669.730 15.200 ;
        RECT 1662.970 15.000 1663.290 15.060 ;
        RECT 1669.410 15.000 1669.730 15.060 ;
      LAYER via ;
        RECT 712.180 126.860 712.440 127.120 ;
        RECT 1663.000 126.860 1663.260 127.120 ;
        RECT 1663.000 15.000 1663.260 15.260 ;
        RECT 1669.440 15.000 1669.700 15.260 ;
      LAYER met2 ;
        RECT 714.370 400.250 714.650 404.000 ;
        RECT 713.160 400.110 714.650 400.250 ;
        RECT 713.160 324.370 713.300 400.110 ;
        RECT 714.370 400.000 714.650 400.110 ;
        RECT 712.240 324.230 713.300 324.370 ;
        RECT 712.240 127.150 712.380 324.230 ;
        RECT 712.180 126.830 712.440 127.150 ;
        RECT 1663.000 126.830 1663.260 127.150 ;
        RECT 1663.060 15.290 1663.200 126.830 ;
        RECT 1663.000 14.970 1663.260 15.290 ;
        RECT 1669.440 14.970 1669.700 15.290 ;
        RECT 1669.500 2.400 1669.640 14.970 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 719.050 127.400 719.370 127.460 ;
        RECT 1683.670 127.400 1683.990 127.460 ;
        RECT 719.050 127.260 1683.990 127.400 ;
        RECT 719.050 127.200 719.370 127.260 ;
        RECT 1683.670 127.200 1683.990 127.260 ;
      LAYER via ;
        RECT 719.080 127.200 719.340 127.460 ;
        RECT 1683.700 127.200 1683.960 127.460 ;
      LAYER met2 ;
        RECT 719.890 400.250 720.170 404.000 ;
        RECT 719.140 400.110 720.170 400.250 ;
        RECT 719.140 127.490 719.280 400.110 ;
        RECT 719.890 400.000 720.170 400.110 ;
        RECT 719.080 127.170 719.340 127.490 ;
        RECT 1683.700 127.170 1683.960 127.490 ;
        RECT 1683.760 82.870 1683.900 127.170 ;
        RECT 1683.760 82.730 1685.280 82.870 ;
        RECT 1685.140 1.770 1685.280 82.730 ;
        RECT 1687.230 1.770 1687.790 2.400 ;
        RECT 1685.140 1.630 1687.790 1.770 ;
        RECT 1687.230 -4.800 1687.790 1.630 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.890 389.880 422.210 389.940 ;
        RECT 423.270 389.880 423.590 389.940 ;
        RECT 421.890 389.740 423.590 389.880 ;
        RECT 421.890 389.680 422.210 389.740 ;
        RECT 423.270 389.680 423.590 389.740 ;
        RECT 421.890 33.220 422.210 33.280 ;
        RECT 545.170 33.220 545.490 33.280 ;
        RECT 421.890 33.080 545.490 33.220 ;
        RECT 421.890 33.020 422.210 33.080 ;
        RECT 545.170 33.020 545.490 33.080 ;
        RECT 545.170 16.560 545.490 16.620 ;
        RECT 729.630 16.560 729.950 16.620 ;
        RECT 545.170 16.420 729.950 16.560 ;
        RECT 545.170 16.360 545.490 16.420 ;
        RECT 729.630 16.360 729.950 16.420 ;
      LAYER via ;
        RECT 421.920 389.680 422.180 389.940 ;
        RECT 423.300 389.680 423.560 389.940 ;
        RECT 421.920 33.020 422.180 33.280 ;
        RECT 545.200 33.020 545.460 33.280 ;
        RECT 545.200 16.360 545.460 16.620 ;
        RECT 729.660 16.360 729.920 16.620 ;
      LAYER met2 ;
        RECT 424.570 400.250 424.850 404.000 ;
        RECT 423.360 400.110 424.850 400.250 ;
        RECT 423.360 389.970 423.500 400.110 ;
        RECT 424.570 400.000 424.850 400.110 ;
        RECT 421.920 389.650 422.180 389.970 ;
        RECT 423.300 389.650 423.560 389.970 ;
        RECT 421.980 33.310 422.120 389.650 ;
        RECT 421.920 32.990 422.180 33.310 ;
        RECT 545.200 32.990 545.460 33.310 ;
        RECT 545.260 16.650 545.400 32.990 ;
        RECT 545.200 16.330 545.460 16.650 ;
        RECT 729.660 16.330 729.920 16.650 ;
        RECT 729.720 2.400 729.860 16.330 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.950 131.140 726.270 131.200 ;
        RECT 1704.370 131.140 1704.690 131.200 ;
        RECT 725.950 131.000 1704.690 131.140 ;
        RECT 725.950 130.940 726.270 131.000 ;
        RECT 1704.370 130.940 1704.690 131.000 ;
      LAYER via ;
        RECT 725.980 130.940 726.240 131.200 ;
        RECT 1704.400 130.940 1704.660 131.200 ;
      LAYER met2 ;
        RECT 724.950 400.250 725.230 404.000 ;
        RECT 724.950 400.110 726.640 400.250 ;
        RECT 724.950 400.000 725.230 400.110 ;
        RECT 726.500 351.970 726.640 400.110 ;
        RECT 726.500 351.830 727.100 351.970 ;
        RECT 726.960 324.370 727.100 351.830 ;
        RECT 726.040 324.230 727.100 324.370 ;
        RECT 726.040 131.230 726.180 324.230 ;
        RECT 725.980 130.910 726.240 131.230 ;
        RECT 1704.400 130.910 1704.660 131.230 ;
        RECT 1704.460 82.870 1704.600 130.910 ;
        RECT 1704.460 82.730 1705.060 82.870 ;
        RECT 1704.920 2.400 1705.060 82.730 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.490 376.280 725.810 376.340 ;
        RECT 729.170 376.280 729.490 376.340 ;
        RECT 725.490 376.140 729.490 376.280 ;
        RECT 725.490 376.080 725.810 376.140 ;
        RECT 729.170 376.080 729.490 376.140 ;
        RECT 725.490 130.800 725.810 130.860 ;
        RECT 1718.170 130.800 1718.490 130.860 ;
        RECT 725.490 130.660 1718.490 130.800 ;
        RECT 725.490 130.600 725.810 130.660 ;
        RECT 1718.170 130.600 1718.490 130.660 ;
      LAYER via ;
        RECT 725.520 376.080 725.780 376.340 ;
        RECT 729.200 376.080 729.460 376.340 ;
        RECT 725.520 130.600 725.780 130.860 ;
        RECT 1718.200 130.600 1718.460 130.860 ;
      LAYER met2 ;
        RECT 730.470 400.250 730.750 404.000 ;
        RECT 729.260 400.110 730.750 400.250 ;
        RECT 729.260 376.370 729.400 400.110 ;
        RECT 730.470 400.000 730.750 400.110 ;
        RECT 725.520 376.050 725.780 376.370 ;
        RECT 729.200 376.050 729.460 376.370 ;
        RECT 725.580 130.890 725.720 376.050 ;
        RECT 725.520 130.570 725.780 130.890 ;
        RECT 1718.200 130.570 1718.460 130.890 ;
        RECT 1718.260 82.870 1718.400 130.570 ;
        RECT 1718.260 82.730 1723.000 82.870 ;
        RECT 1722.860 2.400 1723.000 82.730 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.850 130.460 733.170 130.520 ;
        RECT 1738.870 130.460 1739.190 130.520 ;
        RECT 732.850 130.320 1739.190 130.460 ;
        RECT 732.850 130.260 733.170 130.320 ;
        RECT 1738.870 130.260 1739.190 130.320 ;
      LAYER via ;
        RECT 732.880 130.260 733.140 130.520 ;
        RECT 1738.900 130.260 1739.160 130.520 ;
      LAYER met2 ;
        RECT 735.990 400.250 736.270 404.000 ;
        RECT 734.780 400.110 736.270 400.250 ;
        RECT 734.780 324.370 734.920 400.110 ;
        RECT 735.990 400.000 736.270 400.110 ;
        RECT 732.940 324.230 734.920 324.370 ;
        RECT 732.940 130.550 733.080 324.230 ;
        RECT 732.880 130.230 733.140 130.550 ;
        RECT 1738.900 130.230 1739.160 130.550 ;
        RECT 1738.960 82.870 1739.100 130.230 ;
        RECT 1738.960 82.730 1740.480 82.870 ;
        RECT 1740.340 2.400 1740.480 82.730 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 739.290 130.120 739.610 130.180 ;
        RECT 1752.670 130.120 1752.990 130.180 ;
        RECT 739.290 129.980 1752.990 130.120 ;
        RECT 739.290 129.920 739.610 129.980 ;
        RECT 1752.670 129.920 1752.990 129.980 ;
      LAYER via ;
        RECT 739.320 129.920 739.580 130.180 ;
        RECT 1752.700 129.920 1752.960 130.180 ;
      LAYER met2 ;
        RECT 741.510 400.250 741.790 404.000 ;
        RECT 740.300 400.110 741.790 400.250 ;
        RECT 740.300 324.370 740.440 400.110 ;
        RECT 741.510 400.000 741.790 400.110 ;
        RECT 739.380 324.230 740.440 324.370 ;
        RECT 739.380 130.210 739.520 324.230 ;
        RECT 739.320 129.890 739.580 130.210 ;
        RECT 1752.700 129.890 1752.960 130.210 ;
        RECT 1752.760 82.870 1752.900 129.890 ;
        RECT 1752.760 82.730 1756.120 82.870 ;
        RECT 1755.980 1.770 1756.120 82.730 ;
        RECT 1758.070 1.770 1758.630 2.400 ;
        RECT 1755.980 1.630 1758.630 1.770 ;
        RECT 1758.070 -4.800 1758.630 1.630 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 746.650 129.780 746.970 129.840 ;
        RECT 1773.370 129.780 1773.690 129.840 ;
        RECT 746.650 129.640 1773.690 129.780 ;
        RECT 746.650 129.580 746.970 129.640 ;
        RECT 1773.370 129.580 1773.690 129.640 ;
      LAYER via ;
        RECT 746.680 129.580 746.940 129.840 ;
        RECT 1773.400 129.580 1773.660 129.840 ;
      LAYER met2 ;
        RECT 747.030 400.180 747.310 404.000 ;
        RECT 747.030 400.000 747.340 400.180 ;
        RECT 747.200 351.970 747.340 400.000 ;
        RECT 746.740 351.830 747.340 351.970 ;
        RECT 746.740 129.870 746.880 351.830 ;
        RECT 746.680 129.550 746.940 129.870 ;
        RECT 1773.400 129.550 1773.660 129.870 ;
        RECT 1773.460 82.870 1773.600 129.550 ;
        RECT 1773.460 82.730 1776.360 82.870 ;
        RECT 1776.220 2.400 1776.360 82.730 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 753.090 386.480 753.410 386.540 ;
        RECT 753.550 386.480 753.870 386.540 ;
        RECT 753.090 386.340 753.870 386.480 ;
        RECT 753.090 386.280 753.410 386.340 ;
        RECT 753.550 386.280 753.870 386.340 ;
        RECT 753.090 129.440 753.410 129.500 ;
        RECT 1787.170 129.440 1787.490 129.500 ;
        RECT 753.090 129.300 1787.490 129.440 ;
        RECT 753.090 129.240 753.410 129.300 ;
        RECT 1787.170 129.240 1787.490 129.300 ;
        RECT 1787.170 15.200 1787.490 15.260 ;
        RECT 1793.610 15.200 1793.930 15.260 ;
        RECT 1787.170 15.060 1793.930 15.200 ;
        RECT 1787.170 15.000 1787.490 15.060 ;
        RECT 1793.610 15.000 1793.930 15.060 ;
      LAYER via ;
        RECT 753.120 386.280 753.380 386.540 ;
        RECT 753.580 386.280 753.840 386.540 ;
        RECT 753.120 129.240 753.380 129.500 ;
        RECT 1787.200 129.240 1787.460 129.500 ;
        RECT 1787.200 15.000 1787.460 15.260 ;
        RECT 1793.640 15.000 1793.900 15.260 ;
      LAYER met2 ;
        RECT 752.550 400.250 752.830 404.000 ;
        RECT 752.550 400.110 753.780 400.250 ;
        RECT 752.550 400.000 752.830 400.110 ;
        RECT 753.640 386.570 753.780 400.110 ;
        RECT 753.120 386.250 753.380 386.570 ;
        RECT 753.580 386.250 753.840 386.570 ;
        RECT 753.180 129.530 753.320 386.250 ;
        RECT 753.120 129.210 753.380 129.530 ;
        RECT 1787.200 129.210 1787.460 129.530 ;
        RECT 1787.260 15.290 1787.400 129.210 ;
        RECT 1787.200 14.970 1787.460 15.290 ;
        RECT 1793.640 14.970 1793.900 15.290 ;
        RECT 1793.700 2.400 1793.840 14.970 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 758.150 392.600 758.470 392.660 ;
        RECT 1807.870 392.600 1808.190 392.660 ;
        RECT 758.150 392.460 1808.190 392.600 ;
        RECT 758.150 392.400 758.470 392.460 ;
        RECT 1807.870 392.400 1808.190 392.460 ;
      LAYER via ;
        RECT 758.180 392.400 758.440 392.660 ;
        RECT 1807.900 392.400 1808.160 392.660 ;
      LAYER met2 ;
        RECT 758.070 400.180 758.350 404.000 ;
        RECT 758.070 400.000 758.380 400.180 ;
        RECT 758.240 392.690 758.380 400.000 ;
        RECT 758.180 392.370 758.440 392.690 ;
        RECT 1807.900 392.370 1808.160 392.690 ;
        RECT 1807.960 82.870 1808.100 392.370 ;
        RECT 1807.960 82.730 1809.480 82.870 ;
        RECT 1809.340 1.770 1809.480 82.730 ;
        RECT 1811.430 1.770 1811.990 2.400 ;
        RECT 1809.340 1.630 1811.990 1.770 ;
        RECT 1811.430 -4.800 1811.990 1.630 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.450 129.100 760.770 129.160 ;
        RECT 1828.570 129.100 1828.890 129.160 ;
        RECT 760.450 128.960 1828.890 129.100 ;
        RECT 760.450 128.900 760.770 128.960 ;
        RECT 1828.570 128.900 1828.890 128.960 ;
      LAYER via ;
        RECT 760.480 128.900 760.740 129.160 ;
        RECT 1828.600 128.900 1828.860 129.160 ;
      LAYER met2 ;
        RECT 763.590 400.250 763.870 404.000 ;
        RECT 762.380 400.110 763.870 400.250 ;
        RECT 762.380 324.370 762.520 400.110 ;
        RECT 763.590 400.000 763.870 400.110 ;
        RECT 760.540 324.230 762.520 324.370 ;
        RECT 760.540 129.190 760.680 324.230 ;
        RECT 760.480 128.870 760.740 129.190 ;
        RECT 1828.600 128.870 1828.860 129.190 ;
        RECT 1828.660 82.870 1828.800 128.870 ;
        RECT 1828.660 82.730 1829.260 82.870 ;
        RECT 1829.120 2.400 1829.260 82.730 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 769.190 392.260 769.510 392.320 ;
        RECT 1842.370 392.260 1842.690 392.320 ;
        RECT 769.190 392.120 1842.690 392.260 ;
        RECT 769.190 392.060 769.510 392.120 ;
        RECT 1842.370 392.060 1842.690 392.120 ;
      LAYER via ;
        RECT 769.220 392.060 769.480 392.320 ;
        RECT 1842.400 392.060 1842.660 392.320 ;
      LAYER met2 ;
        RECT 769.110 400.180 769.390 404.000 ;
        RECT 769.110 400.000 769.420 400.180 ;
        RECT 769.280 392.350 769.420 400.000 ;
        RECT 769.220 392.030 769.480 392.350 ;
        RECT 1842.400 392.030 1842.660 392.350 ;
        RECT 1842.460 82.870 1842.600 392.030 ;
        RECT 1842.460 82.730 1847.200 82.870 ;
        RECT 1847.060 2.400 1847.200 82.730 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.790 128.760 774.110 128.820 ;
        RECT 1863.070 128.760 1863.390 128.820 ;
        RECT 773.790 128.620 1863.390 128.760 ;
        RECT 773.790 128.560 774.110 128.620 ;
        RECT 1863.070 128.560 1863.390 128.620 ;
      LAYER via ;
        RECT 773.820 128.560 774.080 128.820 ;
        RECT 1863.100 128.560 1863.360 128.820 ;
      LAYER met2 ;
        RECT 774.170 400.250 774.450 404.000 ;
        RECT 773.880 400.110 774.450 400.250 ;
        RECT 773.880 128.850 774.020 400.110 ;
        RECT 774.170 400.000 774.450 400.110 ;
        RECT 773.820 128.530 774.080 128.850 ;
        RECT 1863.100 128.530 1863.360 128.850 ;
        RECT 1863.160 82.870 1863.300 128.530 ;
        RECT 1863.160 82.730 1864.680 82.870 ;
        RECT 1864.540 2.400 1864.680 82.730 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.170 386.480 430.490 386.540 ;
        RECT 444.890 386.480 445.210 386.540 ;
        RECT 430.170 386.340 445.210 386.480 ;
        RECT 430.170 386.280 430.490 386.340 ;
        RECT 444.890 386.280 445.210 386.340 ;
        RECT 747.570 17.240 747.890 17.300 ;
        RECT 512.140 17.100 747.890 17.240 ;
        RECT 512.140 16.560 512.280 17.100 ;
        RECT 747.570 17.040 747.890 17.100 ;
        RECT 505.700 16.420 512.280 16.560 ;
        RECT 445.350 16.220 445.670 16.280 ;
        RECT 505.700 16.220 505.840 16.420 ;
        RECT 445.350 16.080 505.840 16.220 ;
        RECT 445.350 16.020 445.670 16.080 ;
      LAYER via ;
        RECT 430.200 386.280 430.460 386.540 ;
        RECT 444.920 386.280 445.180 386.540 ;
        RECT 747.600 17.040 747.860 17.300 ;
        RECT 445.380 16.020 445.640 16.280 ;
      LAYER met2 ;
        RECT 430.090 400.180 430.370 404.000 ;
        RECT 430.090 400.000 430.400 400.180 ;
        RECT 430.260 386.570 430.400 400.000 ;
        RECT 430.200 386.250 430.460 386.570 ;
        RECT 444.920 386.250 445.180 386.570 ;
        RECT 444.980 16.730 445.120 386.250 ;
        RECT 747.600 17.010 747.860 17.330 ;
        RECT 444.980 16.590 445.580 16.730 ;
        RECT 445.440 16.310 445.580 16.590 ;
        RECT 445.380 15.990 445.640 16.310 ;
        RECT 747.660 2.400 747.800 17.010 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.690 391.920 781.010 391.980 ;
        RECT 1876.870 391.920 1877.190 391.980 ;
        RECT 780.690 391.780 1877.190 391.920 ;
        RECT 780.690 391.720 781.010 391.780 ;
        RECT 1876.870 391.720 1877.190 391.780 ;
      LAYER via ;
        RECT 780.720 391.720 780.980 391.980 ;
        RECT 1876.900 391.720 1877.160 391.980 ;
      LAYER met2 ;
        RECT 779.690 400.250 779.970 404.000 ;
        RECT 779.690 400.110 780.920 400.250 ;
        RECT 779.690 400.000 779.970 400.110 ;
        RECT 780.780 392.010 780.920 400.110 ;
        RECT 780.720 391.690 780.980 392.010 ;
        RECT 1876.900 391.690 1877.160 392.010 ;
        RECT 1876.960 82.870 1877.100 391.690 ;
        RECT 1876.960 82.730 1880.320 82.870 ;
        RECT 1880.180 1.770 1880.320 82.730 ;
        RECT 1882.270 1.770 1882.830 2.400 ;
        RECT 1880.180 1.630 1882.830 1.770 ;
        RECT 1882.270 -4.800 1882.830 1.630 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.690 128.420 781.010 128.480 ;
        RECT 1897.570 128.420 1897.890 128.480 ;
        RECT 780.690 128.280 1897.890 128.420 ;
        RECT 780.690 128.220 781.010 128.280 ;
        RECT 1897.570 128.220 1897.890 128.280 ;
      LAYER via ;
        RECT 780.720 128.220 780.980 128.480 ;
        RECT 1897.600 128.220 1897.860 128.480 ;
      LAYER met2 ;
        RECT 785.210 400.250 785.490 404.000 ;
        RECT 784.000 400.110 785.490 400.250 ;
        RECT 784.000 399.570 784.140 400.110 ;
        RECT 785.210 400.000 785.490 400.110 ;
        RECT 782.620 399.430 784.140 399.570 ;
        RECT 782.620 324.370 782.760 399.430 ;
        RECT 780.780 324.230 782.760 324.370 ;
        RECT 780.780 128.510 780.920 324.230 ;
        RECT 780.720 128.190 780.980 128.510 ;
        RECT 1897.600 128.190 1897.860 128.510 ;
        RECT 1897.660 1.770 1897.800 128.190 ;
        RECT 1899.750 1.770 1900.310 2.400 ;
        RECT 1897.660 1.630 1900.310 1.770 ;
        RECT 1899.750 -4.800 1900.310 1.630 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 790.810 391.580 791.130 391.640 ;
        RECT 1911.370 391.580 1911.690 391.640 ;
        RECT 790.810 391.440 1911.690 391.580 ;
        RECT 790.810 391.380 791.130 391.440 ;
        RECT 1911.370 391.380 1911.690 391.440 ;
        RECT 1911.370 15.200 1911.690 15.260 ;
        RECT 1917.810 15.200 1918.130 15.260 ;
        RECT 1911.370 15.060 1918.130 15.200 ;
        RECT 1911.370 15.000 1911.690 15.060 ;
        RECT 1917.810 15.000 1918.130 15.060 ;
      LAYER via ;
        RECT 790.840 391.380 791.100 391.640 ;
        RECT 1911.400 391.380 1911.660 391.640 ;
        RECT 1911.400 15.000 1911.660 15.260 ;
        RECT 1917.840 15.000 1918.100 15.260 ;
      LAYER met2 ;
        RECT 790.730 400.180 791.010 404.000 ;
        RECT 790.730 400.000 791.040 400.180 ;
        RECT 790.900 391.670 791.040 400.000 ;
        RECT 790.840 391.350 791.100 391.670 ;
        RECT 1911.400 391.350 1911.660 391.670 ;
        RECT 1911.460 15.290 1911.600 391.350 ;
        RECT 1911.400 14.970 1911.660 15.290 ;
        RECT 1917.840 14.970 1918.100 15.290 ;
        RECT 1917.900 2.400 1918.040 14.970 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.950 128.080 795.270 128.140 ;
        RECT 1932.070 128.080 1932.390 128.140 ;
        RECT 794.950 127.940 1932.390 128.080 ;
        RECT 794.950 127.880 795.270 127.940 ;
        RECT 1932.070 127.880 1932.390 127.940 ;
      LAYER via ;
        RECT 794.980 127.880 795.240 128.140 ;
        RECT 1932.100 127.880 1932.360 128.140 ;
      LAYER met2 ;
        RECT 796.250 400.250 796.530 404.000 ;
        RECT 795.040 400.110 796.530 400.250 ;
        RECT 795.040 128.170 795.180 400.110 ;
        RECT 796.250 400.000 796.530 400.110 ;
        RECT 794.980 127.850 795.240 128.170 ;
        RECT 1932.100 127.850 1932.360 128.170 ;
        RECT 1932.160 82.870 1932.300 127.850 ;
        RECT 1932.160 82.730 1933.680 82.870 ;
        RECT 1933.540 1.770 1933.680 82.730 ;
        RECT 1935.630 1.770 1936.190 2.400 ;
        RECT 1933.540 1.630 1936.190 1.770 ;
        RECT 1935.630 -4.800 1936.190 1.630 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 801.850 391.240 802.170 391.300 ;
        RECT 1952.770 391.240 1953.090 391.300 ;
        RECT 801.850 391.100 1953.090 391.240 ;
        RECT 801.850 391.040 802.170 391.100 ;
        RECT 1952.770 391.040 1953.090 391.100 ;
      LAYER via ;
        RECT 801.880 391.040 802.140 391.300 ;
        RECT 1952.800 391.040 1953.060 391.300 ;
      LAYER met2 ;
        RECT 801.770 400.180 802.050 404.000 ;
        RECT 801.770 400.000 802.080 400.180 ;
        RECT 801.940 391.330 802.080 400.000 ;
        RECT 801.880 391.010 802.140 391.330 ;
        RECT 1952.800 391.010 1953.060 391.330 ;
        RECT 1952.860 82.870 1953.000 391.010 ;
        RECT 1952.860 82.730 1953.460 82.870 ;
        RECT 1953.320 2.400 1953.460 82.730 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.830 398.720 808.150 398.780 ;
        RECT 808.750 398.720 809.070 398.780 ;
        RECT 807.830 398.580 809.070 398.720 ;
        RECT 807.830 398.520 808.150 398.580 ;
        RECT 808.750 398.520 809.070 398.580 ;
        RECT 808.290 127.740 808.610 127.800 ;
        RECT 1966.570 127.740 1966.890 127.800 ;
        RECT 808.290 127.600 1966.890 127.740 ;
        RECT 808.290 127.540 808.610 127.600 ;
        RECT 1966.570 127.540 1966.890 127.600 ;
      LAYER via ;
        RECT 807.860 398.520 808.120 398.780 ;
        RECT 808.780 398.520 809.040 398.780 ;
        RECT 808.320 127.540 808.580 127.800 ;
        RECT 1966.600 127.540 1966.860 127.800 ;
      LAYER met2 ;
        RECT 807.290 400.250 807.570 404.000 ;
        RECT 807.290 400.110 808.060 400.250 ;
        RECT 807.290 400.000 807.570 400.110 ;
        RECT 807.920 398.810 808.060 400.110 ;
        RECT 807.860 398.490 808.120 398.810 ;
        RECT 808.780 398.490 809.040 398.810 ;
        RECT 808.840 351.970 808.980 398.490 ;
        RECT 808.380 351.830 808.980 351.970 ;
        RECT 808.380 127.830 808.520 351.830 ;
        RECT 808.320 127.510 808.580 127.830 ;
        RECT 1966.600 127.510 1966.860 127.830 ;
        RECT 1966.660 82.870 1966.800 127.510 ;
        RECT 1966.660 82.730 1971.400 82.870 ;
        RECT 1971.260 2.400 1971.400 82.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 812.890 390.900 813.210 390.960 ;
        RECT 1987.270 390.900 1987.590 390.960 ;
        RECT 812.890 390.760 1987.590 390.900 ;
        RECT 812.890 390.700 813.210 390.760 ;
        RECT 1987.270 390.700 1987.590 390.760 ;
      LAYER via ;
        RECT 812.920 390.700 813.180 390.960 ;
        RECT 1987.300 390.700 1987.560 390.960 ;
      LAYER met2 ;
        RECT 812.810 400.180 813.090 404.000 ;
        RECT 812.810 400.000 813.120 400.180 ;
        RECT 812.980 390.990 813.120 400.000 ;
        RECT 812.920 390.670 813.180 390.990 ;
        RECT 1987.300 390.670 1987.560 390.990 ;
        RECT 1987.360 82.870 1987.500 390.670 ;
        RECT 1987.360 82.730 1988.880 82.870 ;
        RECT 1988.740 2.400 1988.880 82.730 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.870 400.250 818.150 404.000 ;
        RECT 817.120 400.110 818.150 400.250 ;
        RECT 817.120 324.370 817.260 400.110 ;
        RECT 817.870 400.000 818.150 400.110 ;
        RECT 815.740 324.230 817.260 324.370 ;
        RECT 815.740 127.685 815.880 324.230 ;
        RECT 815.670 127.315 815.950 127.685 ;
        RECT 2001.090 127.315 2001.370 127.685 ;
        RECT 2001.160 82.870 2001.300 127.315 ;
        RECT 2001.160 82.730 2004.520 82.870 ;
        RECT 2004.380 1.770 2004.520 82.730 ;
        RECT 2006.470 1.770 2007.030 2.400 ;
        RECT 2004.380 1.630 2007.030 1.770 ;
        RECT 2006.470 -4.800 2007.030 1.630 ;
      LAYER via2 ;
        RECT 815.670 127.360 815.950 127.640 ;
        RECT 2001.090 127.360 2001.370 127.640 ;
      LAYER met3 ;
        RECT 815.645 127.650 815.975 127.665 ;
        RECT 2001.065 127.650 2001.395 127.665 ;
        RECT 815.645 127.350 2001.395 127.650 ;
        RECT 815.645 127.335 815.975 127.350 ;
        RECT 2001.065 127.335 2001.395 127.350 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 823.470 390.560 823.790 390.620 ;
        RECT 2021.770 390.560 2022.090 390.620 ;
        RECT 823.470 390.420 2022.090 390.560 ;
        RECT 823.470 390.360 823.790 390.420 ;
        RECT 2021.770 390.360 2022.090 390.420 ;
      LAYER via ;
        RECT 823.500 390.360 823.760 390.620 ;
        RECT 2021.800 390.360 2022.060 390.620 ;
      LAYER met2 ;
        RECT 823.390 400.180 823.670 404.000 ;
        RECT 823.390 400.000 823.700 400.180 ;
        RECT 823.560 390.650 823.700 400.000 ;
        RECT 823.500 390.330 823.760 390.650 ;
        RECT 2021.800 390.330 2022.060 390.650 ;
        RECT 2021.860 1.770 2022.000 390.330 ;
        RECT 2023.950 1.770 2024.510 2.400 ;
        RECT 2021.860 1.630 2024.510 1.770 ;
        RECT 2023.950 -4.800 2024.510 1.630 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.990 135.220 829.310 135.280 ;
        RECT 2035.570 135.220 2035.890 135.280 ;
        RECT 828.990 135.080 2035.890 135.220 ;
        RECT 828.990 135.020 829.310 135.080 ;
        RECT 2035.570 135.020 2035.890 135.080 ;
        RECT 2035.570 15.200 2035.890 15.260 ;
        RECT 2042.010 15.200 2042.330 15.260 ;
        RECT 2035.570 15.060 2042.330 15.200 ;
        RECT 2035.570 15.000 2035.890 15.060 ;
        RECT 2042.010 15.000 2042.330 15.060 ;
      LAYER via ;
        RECT 829.020 135.020 829.280 135.280 ;
        RECT 2035.600 135.020 2035.860 135.280 ;
        RECT 2035.600 15.000 2035.860 15.260 ;
        RECT 2042.040 15.000 2042.300 15.260 ;
      LAYER met2 ;
        RECT 828.910 400.250 829.190 404.000 ;
        RECT 828.910 400.110 830.140 400.250 ;
        RECT 828.910 400.000 829.190 400.110 ;
        RECT 830.000 324.370 830.140 400.110 ;
        RECT 829.080 324.230 830.140 324.370 ;
        RECT 829.080 135.310 829.220 324.230 ;
        RECT 829.020 134.990 829.280 135.310 ;
        RECT 2035.600 134.990 2035.860 135.310 ;
        RECT 2035.660 15.290 2035.800 134.990 ;
        RECT 2035.600 14.970 2035.860 15.290 ;
        RECT 2042.040 14.970 2042.300 15.290 ;
        RECT 2042.100 2.400 2042.240 14.970 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.690 33.560 436.010 33.620 ;
        RECT 552.990 33.560 553.310 33.620 ;
        RECT 435.690 33.420 553.310 33.560 ;
        RECT 435.690 33.360 436.010 33.420 ;
        RECT 552.990 33.360 553.310 33.420 ;
        RECT 552.990 19.960 553.310 20.020 ;
        RECT 765.050 19.960 765.370 20.020 ;
        RECT 552.990 19.820 765.370 19.960 ;
        RECT 552.990 19.760 553.310 19.820 ;
        RECT 765.050 19.760 765.370 19.820 ;
      LAYER via ;
        RECT 435.720 33.360 435.980 33.620 ;
        RECT 553.020 33.360 553.280 33.620 ;
        RECT 553.020 19.760 553.280 20.020 ;
        RECT 765.080 19.760 765.340 20.020 ;
      LAYER met2 ;
        RECT 435.610 400.250 435.890 404.000 ;
        RECT 434.860 400.110 435.890 400.250 ;
        RECT 434.860 386.470 435.000 400.110 ;
        RECT 435.610 400.000 435.890 400.110 ;
        RECT 434.860 386.330 435.460 386.470 ;
        RECT 435.320 375.770 435.460 386.330 ;
        RECT 435.320 375.630 435.920 375.770 ;
        RECT 435.780 33.650 435.920 375.630 ;
        RECT 435.720 33.330 435.980 33.650 ;
        RECT 553.020 33.330 553.280 33.650 ;
        RECT 553.080 20.050 553.220 33.330 ;
        RECT 553.020 19.730 553.280 20.050 ;
        RECT 765.080 19.730 765.340 20.050 ;
        RECT 765.140 2.400 765.280 19.730 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 834.510 390.220 834.830 390.280 ;
        RECT 2056.270 390.220 2056.590 390.280 ;
        RECT 834.510 390.080 2056.590 390.220 ;
        RECT 834.510 390.020 834.830 390.080 ;
        RECT 2056.270 390.020 2056.590 390.080 ;
      LAYER via ;
        RECT 834.540 390.020 834.800 390.280 ;
        RECT 2056.300 390.020 2056.560 390.280 ;
      LAYER met2 ;
        RECT 834.430 400.180 834.710 404.000 ;
        RECT 834.430 400.000 834.740 400.180 ;
        RECT 834.600 390.310 834.740 400.000 ;
        RECT 834.540 389.990 834.800 390.310 ;
        RECT 2056.300 389.990 2056.560 390.310 ;
        RECT 2056.360 82.870 2056.500 389.990 ;
        RECT 2056.360 82.730 2059.720 82.870 ;
        RECT 2059.580 2.400 2059.720 82.730 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.890 134.880 836.210 134.940 ;
        RECT 2076.970 134.880 2077.290 134.940 ;
        RECT 835.890 134.740 2077.290 134.880 ;
        RECT 835.890 134.680 836.210 134.740 ;
        RECT 2076.970 134.680 2077.290 134.740 ;
      LAYER via ;
        RECT 835.920 134.680 836.180 134.940 ;
        RECT 2077.000 134.680 2077.260 134.940 ;
      LAYER met2 ;
        RECT 839.950 400.250 840.230 404.000 ;
        RECT 838.740 400.110 840.230 400.250 ;
        RECT 838.740 324.370 838.880 400.110 ;
        RECT 839.950 400.000 840.230 400.110 ;
        RECT 835.980 324.230 838.880 324.370 ;
        RECT 835.980 134.970 836.120 324.230 ;
        RECT 835.920 134.650 836.180 134.970 ;
        RECT 2077.000 134.650 2077.260 134.970 ;
        RECT 2077.060 82.870 2077.200 134.650 ;
        RECT 2077.060 82.730 2077.660 82.870 ;
        RECT 2077.520 2.400 2077.660 82.730 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 845.550 389.880 845.870 389.940 ;
        RECT 2090.770 389.880 2091.090 389.940 ;
        RECT 845.550 389.740 2091.090 389.880 ;
        RECT 845.550 389.680 845.870 389.740 ;
        RECT 2090.770 389.680 2091.090 389.740 ;
      LAYER via ;
        RECT 845.580 389.680 845.840 389.940 ;
        RECT 2090.800 389.680 2091.060 389.940 ;
      LAYER met2 ;
        RECT 845.470 400.180 845.750 404.000 ;
        RECT 845.470 400.000 845.780 400.180 ;
        RECT 845.640 389.970 845.780 400.000 ;
        RECT 845.580 389.650 845.840 389.970 ;
        RECT 2090.800 389.650 2091.060 389.970 ;
        RECT 2090.860 82.870 2091.000 389.650 ;
        RECT 2090.860 82.730 2092.840 82.870 ;
        RECT 2092.700 1.770 2092.840 82.730 ;
        RECT 2094.790 1.770 2095.350 2.400 ;
        RECT 2092.700 1.630 2095.350 1.770 ;
        RECT 2094.790 -4.800 2095.350 1.630 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 850.150 134.540 850.470 134.600 ;
        RECT 2111.470 134.540 2111.790 134.600 ;
        RECT 850.150 134.400 2111.790 134.540 ;
        RECT 850.150 134.340 850.470 134.400 ;
        RECT 2111.470 134.340 2111.790 134.400 ;
      LAYER via ;
        RECT 850.180 134.340 850.440 134.600 ;
        RECT 2111.500 134.340 2111.760 134.600 ;
      LAYER met2 ;
        RECT 850.990 400.250 851.270 404.000 ;
        RECT 850.240 400.110 851.270 400.250 ;
        RECT 850.240 134.630 850.380 400.110 ;
        RECT 850.990 400.000 851.270 400.110 ;
        RECT 850.180 134.310 850.440 134.630 ;
        RECT 2111.500 134.310 2111.760 134.630 ;
        RECT 2111.560 82.870 2111.700 134.310 ;
        RECT 2111.560 82.730 2113.080 82.870 ;
        RECT 2112.940 2.400 2113.080 82.730 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 855.670 15.540 855.990 15.600 ;
        RECT 855.670 15.400 2063.170 15.540 ;
        RECT 855.670 15.340 855.990 15.400 ;
        RECT 2063.030 14.860 2063.170 15.400 ;
        RECT 2130.790 14.860 2131.110 14.920 ;
        RECT 2063.030 14.720 2131.110 14.860 ;
        RECT 2130.790 14.660 2131.110 14.720 ;
      LAYER via ;
        RECT 855.700 15.340 855.960 15.600 ;
        RECT 2130.820 14.660 2131.080 14.920 ;
      LAYER met2 ;
        RECT 856.510 400.250 856.790 404.000 ;
        RECT 855.760 400.110 856.790 400.250 ;
        RECT 855.760 15.630 855.900 400.110 ;
        RECT 856.510 400.000 856.790 400.110 ;
        RECT 855.700 15.310 855.960 15.630 ;
        RECT 2130.820 14.630 2131.080 14.950 ;
        RECT 2130.880 2.400 2131.020 14.630 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.130 386.140 856.450 386.200 ;
        RECT 860.730 386.140 861.050 386.200 ;
        RECT 856.130 386.000 861.050 386.140 ;
        RECT 856.130 385.940 856.450 386.000 ;
        RECT 860.730 385.940 861.050 386.000 ;
        RECT 856.130 15.880 856.450 15.940 ;
        RECT 856.130 15.740 2117.680 15.880 ;
        RECT 856.130 15.680 856.450 15.740 ;
        RECT 2117.540 15.200 2117.680 15.740 ;
        RECT 2148.270 15.200 2148.590 15.260 ;
        RECT 2117.540 15.060 2148.590 15.200 ;
        RECT 2148.270 15.000 2148.590 15.060 ;
      LAYER via ;
        RECT 856.160 385.940 856.420 386.200 ;
        RECT 860.760 385.940 861.020 386.200 ;
        RECT 856.160 15.680 856.420 15.940 ;
        RECT 2148.300 15.000 2148.560 15.260 ;
      LAYER met2 ;
        RECT 862.030 400.250 862.310 404.000 ;
        RECT 860.820 400.110 862.310 400.250 ;
        RECT 860.820 386.230 860.960 400.110 ;
        RECT 862.030 400.000 862.310 400.110 ;
        RECT 856.160 385.910 856.420 386.230 ;
        RECT 860.760 385.910 861.020 386.230 ;
        RECT 856.220 15.970 856.360 385.910 ;
        RECT 856.160 15.650 856.420 15.970 ;
        RECT 2148.300 14.970 2148.560 15.290 ;
        RECT 2148.360 2.400 2148.500 14.970 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 862.570 386.140 862.890 386.200 ;
        RECT 865.790 386.140 866.110 386.200 ;
        RECT 862.570 386.000 866.110 386.140 ;
        RECT 862.570 385.940 862.890 386.000 ;
        RECT 865.790 385.940 866.110 386.000 ;
        RECT 862.570 16.220 862.890 16.280 ;
        RECT 2166.210 16.220 2166.530 16.280 ;
        RECT 862.570 16.080 2166.530 16.220 ;
        RECT 862.570 16.020 862.890 16.080 ;
        RECT 2166.210 16.020 2166.530 16.080 ;
      LAYER via ;
        RECT 862.600 385.940 862.860 386.200 ;
        RECT 865.820 385.940 866.080 386.200 ;
        RECT 862.600 16.020 862.860 16.280 ;
        RECT 2166.240 16.020 2166.500 16.280 ;
      LAYER met2 ;
        RECT 867.090 400.250 867.370 404.000 ;
        RECT 865.880 400.110 867.370 400.250 ;
        RECT 865.880 386.230 866.020 400.110 ;
        RECT 867.090 400.000 867.370 400.110 ;
        RECT 862.600 385.910 862.860 386.230 ;
        RECT 865.820 385.910 866.080 386.230 ;
        RECT 862.660 16.310 862.800 385.910 ;
        RECT 862.600 15.990 862.860 16.310 ;
        RECT 2166.240 15.990 2166.500 16.310 ;
        RECT 2166.300 2.400 2166.440 15.990 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.470 386.480 869.790 386.540 ;
        RECT 871.310 386.480 871.630 386.540 ;
        RECT 869.470 386.340 871.630 386.480 ;
        RECT 869.470 386.280 869.790 386.340 ;
        RECT 871.310 386.280 871.630 386.340 ;
        RECT 869.470 16.560 869.790 16.620 ;
        RECT 2183.690 16.560 2184.010 16.620 ;
        RECT 869.470 16.420 2184.010 16.560 ;
        RECT 869.470 16.360 869.790 16.420 ;
        RECT 2183.690 16.360 2184.010 16.420 ;
      LAYER via ;
        RECT 869.500 386.280 869.760 386.540 ;
        RECT 871.340 386.280 871.600 386.540 ;
        RECT 869.500 16.360 869.760 16.620 ;
        RECT 2183.720 16.360 2183.980 16.620 ;
      LAYER met2 ;
        RECT 872.610 400.250 872.890 404.000 ;
        RECT 871.400 400.110 872.890 400.250 ;
        RECT 871.400 386.570 871.540 400.110 ;
        RECT 872.610 400.000 872.890 400.110 ;
        RECT 869.500 386.250 869.760 386.570 ;
        RECT 871.340 386.250 871.600 386.570 ;
        RECT 869.560 16.650 869.700 386.250 ;
        RECT 869.500 16.330 869.760 16.650 ;
        RECT 2183.720 16.330 2183.980 16.650 ;
        RECT 2183.780 2.400 2183.920 16.330 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.370 386.480 876.690 386.540 ;
        RECT 877.750 386.480 878.070 386.540 ;
        RECT 876.370 386.340 878.070 386.480 ;
        RECT 876.370 386.280 876.690 386.340 ;
        RECT 877.750 386.280 878.070 386.340 ;
        RECT 876.370 16.900 876.690 16.960 ;
        RECT 2201.170 16.900 2201.490 16.960 ;
        RECT 876.370 16.760 2201.490 16.900 ;
        RECT 876.370 16.700 876.690 16.760 ;
        RECT 2201.170 16.700 2201.490 16.760 ;
      LAYER via ;
        RECT 876.400 386.280 876.660 386.540 ;
        RECT 877.780 386.280 878.040 386.540 ;
        RECT 876.400 16.700 876.660 16.960 ;
        RECT 2201.200 16.700 2201.460 16.960 ;
      LAYER met2 ;
        RECT 878.130 400.250 878.410 404.000 ;
        RECT 877.840 400.110 878.410 400.250 ;
        RECT 877.840 386.570 877.980 400.110 ;
        RECT 878.130 400.000 878.410 400.110 ;
        RECT 876.400 386.250 876.660 386.570 ;
        RECT 877.780 386.250 878.040 386.570 ;
        RECT 876.460 16.990 876.600 386.250 ;
        RECT 876.400 16.670 876.660 16.990 ;
        RECT 2201.200 16.670 2201.460 16.990 ;
        RECT 2201.260 8.570 2201.400 16.670 ;
        RECT 2201.260 8.430 2201.860 8.570 ;
        RECT 2201.720 2.400 2201.860 8.430 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.270 20.640 883.590 20.700 ;
        RECT 2219.110 20.640 2219.430 20.700 ;
        RECT 883.270 20.500 2219.430 20.640 ;
        RECT 883.270 20.440 883.590 20.500 ;
        RECT 2219.110 20.440 2219.430 20.500 ;
      LAYER via ;
        RECT 883.300 20.440 883.560 20.700 ;
        RECT 2219.140 20.440 2219.400 20.700 ;
      LAYER met2 ;
        RECT 883.650 400.250 883.930 404.000 ;
        RECT 883.360 400.110 883.930 400.250 ;
        RECT 883.360 20.730 883.500 400.110 ;
        RECT 883.650 400.000 883.930 400.110 ;
        RECT 883.300 20.410 883.560 20.730 ;
        RECT 2219.140 20.410 2219.400 20.730 ;
        RECT 2219.200 2.400 2219.340 20.410 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 376.280 435.090 376.340 ;
        RECT 439.370 376.280 439.690 376.340 ;
        RECT 434.770 376.140 439.690 376.280 ;
        RECT 434.770 376.080 435.090 376.140 ;
        RECT 439.370 376.080 439.690 376.140 ;
      LAYER via ;
        RECT 434.800 376.080 435.060 376.340 ;
        RECT 439.400 376.080 439.660 376.340 ;
      LAYER met2 ;
        RECT 440.670 400.250 440.950 404.000 ;
        RECT 439.460 400.110 440.950 400.250 ;
        RECT 439.460 376.370 439.600 400.110 ;
        RECT 440.670 400.000 440.950 400.110 ;
        RECT 434.800 376.050 435.060 376.370 ;
        RECT 439.400 376.050 439.660 376.370 ;
        RECT 434.860 17.525 435.000 376.050 ;
        RECT 434.790 17.155 435.070 17.525 ;
        RECT 783.010 17.155 783.290 17.525 ;
        RECT 783.080 2.400 783.220 17.155 ;
        RECT 782.870 -4.800 783.430 2.400 ;
      LAYER via2 ;
        RECT 434.790 17.200 435.070 17.480 ;
        RECT 783.010 17.200 783.290 17.480 ;
      LAYER met3 ;
        RECT 434.765 17.490 435.095 17.505 ;
        RECT 782.985 17.490 783.315 17.505 ;
        RECT 434.765 17.190 783.315 17.490 ;
        RECT 434.765 17.175 435.095 17.190 ;
        RECT 782.985 17.175 783.315 17.190 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.730 386.480 884.050 386.540 ;
        RECT 887.870 386.480 888.190 386.540 ;
        RECT 883.730 386.340 888.190 386.480 ;
        RECT 883.730 386.280 884.050 386.340 ;
        RECT 887.870 386.280 888.190 386.340 ;
        RECT 883.730 20.300 884.050 20.360 ;
        RECT 2237.050 20.300 2237.370 20.360 ;
        RECT 883.730 20.160 2237.370 20.300 ;
        RECT 883.730 20.100 884.050 20.160 ;
        RECT 2237.050 20.100 2237.370 20.160 ;
      LAYER via ;
        RECT 883.760 386.280 884.020 386.540 ;
        RECT 887.900 386.280 888.160 386.540 ;
        RECT 883.760 20.100 884.020 20.360 ;
        RECT 2237.080 20.100 2237.340 20.360 ;
      LAYER met2 ;
        RECT 889.170 400.250 889.450 404.000 ;
        RECT 887.960 400.110 889.450 400.250 ;
        RECT 887.960 386.570 888.100 400.110 ;
        RECT 889.170 400.000 889.450 400.110 ;
        RECT 883.760 386.250 884.020 386.570 ;
        RECT 887.900 386.250 888.160 386.570 ;
        RECT 883.820 20.390 883.960 386.250 ;
        RECT 883.760 20.070 884.020 20.390 ;
        RECT 2237.080 20.070 2237.340 20.390 ;
        RECT 2237.140 2.400 2237.280 20.070 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.170 377.980 890.490 378.040 ;
        RECT 893.390 377.980 893.710 378.040 ;
        RECT 890.170 377.840 893.710 377.980 ;
        RECT 890.170 377.780 890.490 377.840 ;
        RECT 893.390 377.780 893.710 377.840 ;
        RECT 890.170 19.960 890.490 20.020 ;
        RECT 2254.530 19.960 2254.850 20.020 ;
        RECT 890.170 19.820 2254.850 19.960 ;
        RECT 890.170 19.760 890.490 19.820 ;
        RECT 2254.530 19.760 2254.850 19.820 ;
      LAYER via ;
        RECT 890.200 377.780 890.460 378.040 ;
        RECT 893.420 377.780 893.680 378.040 ;
        RECT 890.200 19.760 890.460 20.020 ;
        RECT 2254.560 19.760 2254.820 20.020 ;
      LAYER met2 ;
        RECT 894.690 400.250 894.970 404.000 ;
        RECT 893.480 400.110 894.970 400.250 ;
        RECT 893.480 378.070 893.620 400.110 ;
        RECT 894.690 400.000 894.970 400.110 ;
        RECT 890.200 377.750 890.460 378.070 ;
        RECT 893.420 377.750 893.680 378.070 ;
        RECT 890.260 20.050 890.400 377.750 ;
        RECT 890.200 19.730 890.460 20.050 ;
        RECT 2254.560 19.730 2254.820 20.050 ;
        RECT 2254.620 2.400 2254.760 19.730 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.070 384.440 897.390 384.500 ;
        RECT 898.910 384.440 899.230 384.500 ;
        RECT 897.070 384.300 899.230 384.440 ;
        RECT 897.070 384.240 897.390 384.300 ;
        RECT 898.910 384.240 899.230 384.300 ;
        RECT 897.070 19.620 897.390 19.680 ;
        RECT 2272.470 19.620 2272.790 19.680 ;
        RECT 897.070 19.480 2272.790 19.620 ;
        RECT 897.070 19.420 897.390 19.480 ;
        RECT 2272.470 19.420 2272.790 19.480 ;
      LAYER via ;
        RECT 897.100 384.240 897.360 384.500 ;
        RECT 898.940 384.240 899.200 384.500 ;
        RECT 897.100 19.420 897.360 19.680 ;
        RECT 2272.500 19.420 2272.760 19.680 ;
      LAYER met2 ;
        RECT 900.210 400.250 900.490 404.000 ;
        RECT 899.000 400.110 900.490 400.250 ;
        RECT 899.000 384.530 899.140 400.110 ;
        RECT 900.210 400.000 900.490 400.110 ;
        RECT 897.100 384.210 897.360 384.530 ;
        RECT 898.940 384.210 899.200 384.530 ;
        RECT 897.160 19.710 897.300 384.210 ;
        RECT 897.100 19.390 897.360 19.710 ;
        RECT 2272.500 19.390 2272.760 19.710 ;
        RECT 2272.560 2.400 2272.700 19.390 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 903.970 386.140 904.290 386.200 ;
        RECT 905.350 386.140 905.670 386.200 ;
        RECT 903.970 386.000 905.670 386.140 ;
        RECT 903.970 385.940 904.290 386.000 ;
        RECT 905.350 385.940 905.670 386.000 ;
        RECT 903.970 19.280 904.290 19.340 ;
        RECT 2290.410 19.280 2290.730 19.340 ;
        RECT 903.970 19.140 2290.730 19.280 ;
        RECT 903.970 19.080 904.290 19.140 ;
        RECT 2290.410 19.080 2290.730 19.140 ;
      LAYER via ;
        RECT 904.000 385.940 904.260 386.200 ;
        RECT 905.380 385.940 905.640 386.200 ;
        RECT 904.000 19.080 904.260 19.340 ;
        RECT 2290.440 19.080 2290.700 19.340 ;
      LAYER met2 ;
        RECT 905.730 400.250 906.010 404.000 ;
        RECT 905.440 400.110 906.010 400.250 ;
        RECT 905.440 386.230 905.580 400.110 ;
        RECT 905.730 400.000 906.010 400.110 ;
        RECT 904.000 385.910 904.260 386.230 ;
        RECT 905.380 385.910 905.640 386.230 ;
        RECT 904.060 19.370 904.200 385.910 ;
        RECT 904.000 19.050 904.260 19.370 ;
        RECT 2290.440 19.050 2290.700 19.370 ;
        RECT 2290.500 2.400 2290.640 19.050 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 910.870 18.940 911.190 19.000 ;
        RECT 2307.890 18.940 2308.210 19.000 ;
        RECT 910.870 18.800 2308.210 18.940 ;
        RECT 910.870 18.740 911.190 18.800 ;
        RECT 2307.890 18.740 2308.210 18.800 ;
      LAYER via ;
        RECT 910.900 18.740 911.160 19.000 ;
        RECT 2307.920 18.740 2308.180 19.000 ;
      LAYER met2 ;
        RECT 911.250 400.250 911.530 404.000 ;
        RECT 910.960 400.110 911.530 400.250 ;
        RECT 910.960 19.030 911.100 400.110 ;
        RECT 911.250 400.000 911.530 400.110 ;
        RECT 910.900 18.710 911.160 19.030 ;
        RECT 2307.920 18.710 2308.180 19.030 ;
        RECT 2307.980 2.400 2308.120 18.710 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.330 386.480 911.650 386.540 ;
        RECT 915.010 386.480 915.330 386.540 ;
        RECT 911.330 386.340 915.330 386.480 ;
        RECT 911.330 386.280 911.650 386.340 ;
        RECT 915.010 386.280 915.330 386.340 ;
        RECT 911.330 18.600 911.650 18.660 ;
        RECT 2325.830 18.600 2326.150 18.660 ;
        RECT 911.330 18.460 2326.150 18.600 ;
        RECT 911.330 18.400 911.650 18.460 ;
        RECT 2325.830 18.400 2326.150 18.460 ;
      LAYER via ;
        RECT 911.360 386.280 911.620 386.540 ;
        RECT 915.040 386.280 915.300 386.540 ;
        RECT 911.360 18.400 911.620 18.660 ;
        RECT 2325.860 18.400 2326.120 18.660 ;
      LAYER met2 ;
        RECT 916.310 400.250 916.590 404.000 ;
        RECT 915.100 400.110 916.590 400.250 ;
        RECT 915.100 386.570 915.240 400.110 ;
        RECT 916.310 400.000 916.590 400.110 ;
        RECT 911.360 386.250 911.620 386.570 ;
        RECT 915.040 386.250 915.300 386.570 ;
        RECT 911.420 18.690 911.560 386.250 ;
        RECT 911.360 18.370 911.620 18.690 ;
        RECT 2325.860 18.370 2326.120 18.690 ;
        RECT 2325.920 2.400 2326.060 18.370 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 917.770 386.140 918.090 386.200 ;
        RECT 920.530 386.140 920.850 386.200 ;
        RECT 917.770 386.000 920.850 386.140 ;
        RECT 917.770 385.940 918.090 386.000 ;
        RECT 920.530 385.940 920.850 386.000 ;
        RECT 917.770 18.260 918.090 18.320 ;
        RECT 2343.310 18.260 2343.630 18.320 ;
        RECT 917.770 18.120 2343.630 18.260 ;
        RECT 917.770 18.060 918.090 18.120 ;
        RECT 2343.310 18.060 2343.630 18.120 ;
      LAYER via ;
        RECT 917.800 385.940 918.060 386.200 ;
        RECT 920.560 385.940 920.820 386.200 ;
        RECT 917.800 18.060 918.060 18.320 ;
        RECT 2343.340 18.060 2343.600 18.320 ;
      LAYER met2 ;
        RECT 921.830 400.250 922.110 404.000 ;
        RECT 920.620 400.110 922.110 400.250 ;
        RECT 920.620 386.230 920.760 400.110 ;
        RECT 921.830 400.000 922.110 400.110 ;
        RECT 917.800 385.910 918.060 386.230 ;
        RECT 920.560 385.910 920.820 386.230 ;
        RECT 917.860 18.350 918.000 385.910 ;
        RECT 917.800 18.030 918.060 18.350 ;
        RECT 2343.340 18.030 2343.600 18.350 ;
        RECT 2343.400 2.400 2343.540 18.030 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 924.670 386.480 924.990 386.540 ;
        RECT 926.510 386.480 926.830 386.540 ;
        RECT 924.670 386.340 926.830 386.480 ;
        RECT 924.670 386.280 924.990 386.340 ;
        RECT 926.510 386.280 926.830 386.340 ;
        RECT 924.670 17.920 924.990 17.980 ;
        RECT 2361.250 17.920 2361.570 17.980 ;
        RECT 924.670 17.780 2361.570 17.920 ;
        RECT 924.670 17.720 924.990 17.780 ;
        RECT 2361.250 17.720 2361.570 17.780 ;
      LAYER via ;
        RECT 924.700 386.280 924.960 386.540 ;
        RECT 926.540 386.280 926.800 386.540 ;
        RECT 924.700 17.720 924.960 17.980 ;
        RECT 2361.280 17.720 2361.540 17.980 ;
      LAYER met2 ;
        RECT 927.350 400.250 927.630 404.000 ;
        RECT 926.600 400.110 927.630 400.250 ;
        RECT 926.600 386.570 926.740 400.110 ;
        RECT 927.350 400.000 927.630 400.110 ;
        RECT 924.700 386.250 924.960 386.570 ;
        RECT 926.540 386.250 926.800 386.570 ;
        RECT 924.760 18.010 924.900 386.250 ;
        RECT 924.700 17.690 924.960 18.010 ;
        RECT 2361.280 17.690 2361.540 18.010 ;
        RECT 2361.340 2.400 2361.480 17.690 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 17.580 931.890 17.640 ;
        RECT 931.570 17.440 2366.080 17.580 ;
        RECT 931.570 17.380 931.890 17.440 ;
        RECT 2365.940 17.240 2366.080 17.440 ;
        RECT 2378.730 17.240 2379.050 17.300 ;
        RECT 2365.940 17.100 2379.050 17.240 ;
        RECT 2378.730 17.040 2379.050 17.100 ;
      LAYER via ;
        RECT 931.600 17.380 931.860 17.640 ;
        RECT 2378.760 17.040 2379.020 17.300 ;
      LAYER met2 ;
        RECT 932.870 400.250 933.150 404.000 ;
        RECT 931.660 400.110 933.150 400.250 ;
        RECT 931.660 17.670 931.800 400.110 ;
        RECT 932.870 400.000 933.150 400.110 ;
        RECT 931.600 17.350 931.860 17.670 ;
        RECT 2378.760 17.010 2379.020 17.330 ;
        RECT 2378.820 2.400 2378.960 17.010 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.470 17.240 938.790 17.300 ;
        RECT 938.470 17.100 2352.970 17.240 ;
        RECT 938.470 17.040 938.790 17.100 ;
        RECT 2352.830 16.900 2352.970 17.100 ;
        RECT 2396.670 16.900 2396.990 16.960 ;
        RECT 2352.830 16.760 2396.990 16.900 ;
        RECT 2396.670 16.700 2396.990 16.760 ;
      LAYER via ;
        RECT 938.500 17.040 938.760 17.300 ;
        RECT 2396.700 16.700 2396.960 16.960 ;
      LAYER met2 ;
        RECT 938.390 400.180 938.670 404.000 ;
        RECT 938.390 400.000 938.700 400.180 ;
        RECT 938.560 17.330 938.700 400.000 ;
        RECT 938.500 17.010 938.760 17.330 ;
        RECT 2396.700 16.670 2396.960 16.990 ;
        RECT 2396.760 2.400 2396.900 16.670 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.270 386.480 446.590 386.540 ;
        RECT 451.790 386.480 452.110 386.540 ;
        RECT 446.270 386.340 452.110 386.480 ;
        RECT 446.270 386.280 446.590 386.340 ;
        RECT 451.790 386.280 452.110 386.340 ;
      LAYER via ;
        RECT 446.300 386.280 446.560 386.540 ;
        RECT 451.820 386.280 452.080 386.540 ;
      LAYER met2 ;
        RECT 446.190 400.180 446.470 404.000 ;
        RECT 446.190 400.000 446.500 400.180 ;
        RECT 446.360 386.570 446.500 400.000 ;
        RECT 446.300 386.250 446.560 386.570 ;
        RECT 451.820 386.250 452.080 386.570 ;
        RECT 451.880 82.870 452.020 386.250 ;
        RECT 451.880 82.730 452.480 82.870 ;
        RECT 452.340 16.845 452.480 82.730 ;
        RECT 452.270 16.475 452.550 16.845 ;
        RECT 800.490 16.475 800.770 16.845 ;
        RECT 800.560 2.400 800.700 16.475 ;
        RECT 800.350 -4.800 800.910 2.400 ;
      LAYER via2 ;
        RECT 452.270 16.520 452.550 16.800 ;
        RECT 800.490 16.520 800.770 16.800 ;
      LAYER met3 ;
        RECT 452.245 16.810 452.575 16.825 ;
        RECT 800.465 16.810 800.795 16.825 ;
        RECT 452.245 16.510 800.795 16.810 ;
        RECT 452.245 16.495 452.575 16.510 ;
        RECT 800.465 16.495 800.795 16.510 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 427.960 1117.730 428.020 ;
        RECT 2645.990 427.960 2646.310 428.020 ;
        RECT 1117.410 427.820 2646.310 427.960 ;
        RECT 1117.410 427.760 1117.730 427.820 ;
        RECT 2645.990 427.760 2646.310 427.820 ;
        RECT 2645.990 17.240 2646.310 17.300 ;
        RECT 2898.990 17.240 2899.310 17.300 ;
        RECT 2645.990 17.100 2899.310 17.240 ;
        RECT 2645.990 17.040 2646.310 17.100 ;
        RECT 2898.990 17.040 2899.310 17.100 ;
      LAYER via ;
        RECT 1117.440 427.760 1117.700 428.020 ;
        RECT 2646.020 427.760 2646.280 428.020 ;
        RECT 2646.020 17.040 2646.280 17.300 ;
        RECT 2899.020 17.040 2899.280 17.300 ;
      LAYER met2 ;
        RECT 1117.430 428.555 1117.710 428.925 ;
        RECT 1117.500 428.050 1117.640 428.555 ;
        RECT 1117.440 427.730 1117.700 428.050 ;
        RECT 2646.020 427.730 2646.280 428.050 ;
        RECT 2646.080 17.330 2646.220 427.730 ;
        RECT 2646.020 17.010 2646.280 17.330 ;
        RECT 2899.020 17.010 2899.280 17.330 ;
        RECT 2899.080 2.400 2899.220 17.010 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 1117.430 428.600 1117.710 428.880 ;
      LAYER met3 ;
        RECT 1096.000 429.960 1100.000 430.560 ;
        RECT 1098.790 428.890 1099.090 429.960 ;
        RECT 1117.405 428.890 1117.735 428.905 ;
        RECT 1098.790 428.590 1117.735 428.890 ;
        RECT 1117.405 428.575 1117.735 428.590 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 525.795 193.110 526.165 ;
        RECT 192.900 65.125 193.040 525.795 ;
        RECT 192.830 64.755 193.110 65.125 ;
        RECT 2904.990 64.755 2905.270 65.125 ;
        RECT 2905.060 2.400 2905.200 64.755 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 192.830 525.840 193.110 526.120 ;
        RECT 192.830 64.800 193.110 65.080 ;
        RECT 2904.990 64.800 2905.270 65.080 ;
      LAYER met3 ;
        RECT 200.000 528.560 204.000 529.160 ;
        RECT 192.805 526.130 193.135 526.145 ;
        RECT 200.870 526.130 201.170 528.560 ;
        RECT 192.805 525.830 201.170 526.130 ;
        RECT 192.805 525.815 193.135 525.830 ;
        RECT 192.805 65.090 193.135 65.105 ;
        RECT 2904.965 65.090 2905.295 65.105 ;
        RECT 192.805 64.790 2905.295 65.090 ;
        RECT 192.805 64.775 193.135 64.790 ;
        RECT 2904.965 64.775 2905.295 64.790 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 546.875 1114.950 547.245 ;
        RECT 1114.740 16.845 1114.880 546.875 ;
        RECT 1114.670 16.475 1114.950 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1114.670 546.920 1114.950 547.200 ;
        RECT 1114.670 16.520 1114.950 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
      LAYER met3 ;
        RECT 1096.000 549.640 1100.000 550.240 ;
        RECT 1098.790 547.210 1099.090 549.640 ;
        RECT 1114.645 547.210 1114.975 547.225 ;
        RECT 1098.790 546.910 1114.975 547.210 ;
        RECT 1114.645 546.895 1114.975 546.910 ;
        RECT 1114.645 16.810 1114.975 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 1114.645 16.510 2911.275 16.810 ;
        RECT 1114.645 16.495 1114.975 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1019.890 1007.660 1020.210 1007.720 ;
        RECT 1348.790 1007.660 1349.110 1007.720 ;
        RECT 1019.890 1007.520 1349.110 1007.660 ;
        RECT 1019.890 1007.460 1020.210 1007.520 ;
        RECT 1348.790 1007.460 1349.110 1007.520 ;
      LAYER via ;
        RECT 1019.920 1007.460 1020.180 1007.720 ;
        RECT 1348.820 1007.460 1349.080 1007.720 ;
      LAYER met2 ;
        RECT 1019.920 1007.430 1020.180 1007.750 ;
        RECT 1348.820 1007.430 1349.080 1007.750 ;
        RECT 1018.430 999.330 1018.710 1000.000 ;
        RECT 1019.980 999.330 1020.120 1007.430 ;
        RECT 1018.430 999.190 1020.120 999.330 ;
        RECT 1018.430 996.000 1018.710 999.190 ;
        RECT 1348.880 18.205 1349.020 1007.430 ;
        RECT 1348.810 17.835 1349.090 18.205 ;
        RECT 2916.950 17.155 2917.230 17.525 ;
        RECT 2917.020 2.400 2917.160 17.155 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
      LAYER via2 ;
        RECT 1348.810 17.880 1349.090 18.160 ;
        RECT 2916.950 17.200 2917.230 17.480 ;
      LAYER met3 ;
        RECT 1348.785 18.170 1349.115 18.185 ;
        RECT 1348.785 17.870 1387.050 18.170 ;
        RECT 1348.785 17.855 1349.115 17.870 ;
        RECT 1386.750 17.490 1387.050 17.870 ;
        RECT 2916.925 17.490 2917.255 17.505 ;
        RECT 1386.750 17.190 2917.255 17.490 ;
        RECT 2916.925 17.175 2917.255 17.190 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
        RECT 188.970 1010.000 192.070 3529.150 ;
        RECT 368.970 1010.000 372.070 3529.150 ;
        RECT 548.970 1010.000 552.070 3529.150 ;
        RECT 728.970 1010.000 732.070 3529.150 ;
        RECT 908.970 1010.000 912.070 3529.150 ;
        RECT 1088.970 1010.000 1092.070 3529.150 ;
        RECT 221.040 410.640 222.640 987.760 ;
        RECT 374.640 410.640 376.240 987.760 ;
        RECT 528.240 410.640 529.840 987.760 ;
        RECT 681.840 410.640 683.440 987.760 ;
        RECT 835.440 410.640 837.040 987.760 ;
        RECT 989.040 410.640 990.640 987.760 ;
        RECT 188.970 -9.470 192.070 390.000 ;
        RECT 368.970 -9.470 372.070 390.000 ;
        RECT 548.970 -9.470 552.070 390.000 ;
        RECT 728.970 -9.470 732.070 390.000 ;
        RECT 908.970 -9.470 912.070 390.000 ;
        RECT 1088.970 -9.470 1092.070 390.000 ;
        RECT 1268.970 -9.470 1272.070 3529.150 ;
        RECT 1448.970 -9.470 1452.070 3529.150 ;
        RECT 1628.970 -9.470 1632.070 3529.150 ;
        RECT 1808.970 -9.470 1812.070 3529.150 ;
        RECT 1988.970 -9.470 1992.070 3529.150 ;
        RECT 2168.970 -9.470 2172.070 3529.150 ;
        RECT 2348.970 -9.470 2352.070 3529.150 ;
        RECT 2528.970 -9.470 2532.070 3529.150 ;
        RECT 2708.970 -9.470 2712.070 3529.150 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER via4 ;
        RECT -9.870 3523.010 -8.690 3524.190 ;
        RECT -8.270 3523.010 -7.090 3524.190 ;
        RECT -9.870 3521.410 -8.690 3522.590 ;
        RECT -8.270 3521.410 -7.090 3522.590 ;
        RECT -9.870 3436.090 -8.690 3437.270 ;
        RECT -8.270 3436.090 -7.090 3437.270 ;
        RECT -9.870 3434.490 -8.690 3435.670 ;
        RECT -8.270 3434.490 -7.090 3435.670 ;
        RECT -9.870 3256.090 -8.690 3257.270 ;
        RECT -8.270 3256.090 -7.090 3257.270 ;
        RECT -9.870 3254.490 -8.690 3255.670 ;
        RECT -8.270 3254.490 -7.090 3255.670 ;
        RECT -9.870 3076.090 -8.690 3077.270 ;
        RECT -8.270 3076.090 -7.090 3077.270 ;
        RECT -9.870 3074.490 -8.690 3075.670 ;
        RECT -8.270 3074.490 -7.090 3075.670 ;
        RECT -9.870 2896.090 -8.690 2897.270 ;
        RECT -8.270 2896.090 -7.090 2897.270 ;
        RECT -9.870 2894.490 -8.690 2895.670 ;
        RECT -8.270 2894.490 -7.090 2895.670 ;
        RECT -9.870 2716.090 -8.690 2717.270 ;
        RECT -8.270 2716.090 -7.090 2717.270 ;
        RECT -9.870 2714.490 -8.690 2715.670 ;
        RECT -8.270 2714.490 -7.090 2715.670 ;
        RECT -9.870 2536.090 -8.690 2537.270 ;
        RECT -8.270 2536.090 -7.090 2537.270 ;
        RECT -9.870 2534.490 -8.690 2535.670 ;
        RECT -8.270 2534.490 -7.090 2535.670 ;
        RECT -9.870 2356.090 -8.690 2357.270 ;
        RECT -8.270 2356.090 -7.090 2357.270 ;
        RECT -9.870 2354.490 -8.690 2355.670 ;
        RECT -8.270 2354.490 -7.090 2355.670 ;
        RECT -9.870 2176.090 -8.690 2177.270 ;
        RECT -8.270 2176.090 -7.090 2177.270 ;
        RECT -9.870 2174.490 -8.690 2175.670 ;
        RECT -8.270 2174.490 -7.090 2175.670 ;
        RECT -9.870 1996.090 -8.690 1997.270 ;
        RECT -8.270 1996.090 -7.090 1997.270 ;
        RECT -9.870 1994.490 -8.690 1995.670 ;
        RECT -8.270 1994.490 -7.090 1995.670 ;
        RECT -9.870 1816.090 -8.690 1817.270 ;
        RECT -8.270 1816.090 -7.090 1817.270 ;
        RECT -9.870 1814.490 -8.690 1815.670 ;
        RECT -8.270 1814.490 -7.090 1815.670 ;
        RECT -9.870 1636.090 -8.690 1637.270 ;
        RECT -8.270 1636.090 -7.090 1637.270 ;
        RECT -9.870 1634.490 -8.690 1635.670 ;
        RECT -8.270 1634.490 -7.090 1635.670 ;
        RECT -9.870 1456.090 -8.690 1457.270 ;
        RECT -8.270 1456.090 -7.090 1457.270 ;
        RECT -9.870 1454.490 -8.690 1455.670 ;
        RECT -8.270 1454.490 -7.090 1455.670 ;
        RECT -9.870 1276.090 -8.690 1277.270 ;
        RECT -8.270 1276.090 -7.090 1277.270 ;
        RECT -9.870 1274.490 -8.690 1275.670 ;
        RECT -8.270 1274.490 -7.090 1275.670 ;
        RECT -9.870 1096.090 -8.690 1097.270 ;
        RECT -8.270 1096.090 -7.090 1097.270 ;
        RECT -9.870 1094.490 -8.690 1095.670 ;
        RECT -8.270 1094.490 -7.090 1095.670 ;
        RECT -9.870 916.090 -8.690 917.270 ;
        RECT -8.270 916.090 -7.090 917.270 ;
        RECT -9.870 914.490 -8.690 915.670 ;
        RECT -8.270 914.490 -7.090 915.670 ;
        RECT -9.870 736.090 -8.690 737.270 ;
        RECT -8.270 736.090 -7.090 737.270 ;
        RECT -9.870 734.490 -8.690 735.670 ;
        RECT -8.270 734.490 -7.090 735.670 ;
        RECT -9.870 556.090 -8.690 557.270 ;
        RECT -8.270 556.090 -7.090 557.270 ;
        RECT -9.870 554.490 -8.690 555.670 ;
        RECT -8.270 554.490 -7.090 555.670 ;
        RECT -9.870 376.090 -8.690 377.270 ;
        RECT -8.270 376.090 -7.090 377.270 ;
        RECT -9.870 374.490 -8.690 375.670 ;
        RECT -8.270 374.490 -7.090 375.670 ;
        RECT -9.870 196.090 -8.690 197.270 ;
        RECT -8.270 196.090 -7.090 197.270 ;
        RECT -9.870 194.490 -8.690 195.670 ;
        RECT -8.270 194.490 -7.090 195.670 ;
        RECT -9.870 16.090 -8.690 17.270 ;
        RECT -8.270 16.090 -7.090 17.270 ;
        RECT -9.870 14.490 -8.690 15.670 ;
        RECT -8.270 14.490 -7.090 15.670 ;
        RECT -9.870 -2.910 -8.690 -1.730 ;
        RECT -8.270 -2.910 -7.090 -1.730 ;
        RECT -9.870 -4.510 -8.690 -3.330 ;
        RECT -8.270 -4.510 -7.090 -3.330 ;
        RECT 9.130 3523.010 10.310 3524.190 ;
        RECT 10.730 3523.010 11.910 3524.190 ;
        RECT 9.130 3521.410 10.310 3522.590 ;
        RECT 10.730 3521.410 11.910 3522.590 ;
        RECT 9.130 3436.090 10.310 3437.270 ;
        RECT 10.730 3436.090 11.910 3437.270 ;
        RECT 9.130 3434.490 10.310 3435.670 ;
        RECT 10.730 3434.490 11.910 3435.670 ;
        RECT 9.130 3256.090 10.310 3257.270 ;
        RECT 10.730 3256.090 11.910 3257.270 ;
        RECT 9.130 3254.490 10.310 3255.670 ;
        RECT 10.730 3254.490 11.910 3255.670 ;
        RECT 9.130 3076.090 10.310 3077.270 ;
        RECT 10.730 3076.090 11.910 3077.270 ;
        RECT 9.130 3074.490 10.310 3075.670 ;
        RECT 10.730 3074.490 11.910 3075.670 ;
        RECT 9.130 2896.090 10.310 2897.270 ;
        RECT 10.730 2896.090 11.910 2897.270 ;
        RECT 9.130 2894.490 10.310 2895.670 ;
        RECT 10.730 2894.490 11.910 2895.670 ;
        RECT 9.130 2716.090 10.310 2717.270 ;
        RECT 10.730 2716.090 11.910 2717.270 ;
        RECT 9.130 2714.490 10.310 2715.670 ;
        RECT 10.730 2714.490 11.910 2715.670 ;
        RECT 9.130 2536.090 10.310 2537.270 ;
        RECT 10.730 2536.090 11.910 2537.270 ;
        RECT 9.130 2534.490 10.310 2535.670 ;
        RECT 10.730 2534.490 11.910 2535.670 ;
        RECT 9.130 2356.090 10.310 2357.270 ;
        RECT 10.730 2356.090 11.910 2357.270 ;
        RECT 9.130 2354.490 10.310 2355.670 ;
        RECT 10.730 2354.490 11.910 2355.670 ;
        RECT 9.130 2176.090 10.310 2177.270 ;
        RECT 10.730 2176.090 11.910 2177.270 ;
        RECT 9.130 2174.490 10.310 2175.670 ;
        RECT 10.730 2174.490 11.910 2175.670 ;
        RECT 9.130 1996.090 10.310 1997.270 ;
        RECT 10.730 1996.090 11.910 1997.270 ;
        RECT 9.130 1994.490 10.310 1995.670 ;
        RECT 10.730 1994.490 11.910 1995.670 ;
        RECT 9.130 1816.090 10.310 1817.270 ;
        RECT 10.730 1816.090 11.910 1817.270 ;
        RECT 9.130 1814.490 10.310 1815.670 ;
        RECT 10.730 1814.490 11.910 1815.670 ;
        RECT 9.130 1636.090 10.310 1637.270 ;
        RECT 10.730 1636.090 11.910 1637.270 ;
        RECT 9.130 1634.490 10.310 1635.670 ;
        RECT 10.730 1634.490 11.910 1635.670 ;
        RECT 9.130 1456.090 10.310 1457.270 ;
        RECT 10.730 1456.090 11.910 1457.270 ;
        RECT 9.130 1454.490 10.310 1455.670 ;
        RECT 10.730 1454.490 11.910 1455.670 ;
        RECT 9.130 1276.090 10.310 1277.270 ;
        RECT 10.730 1276.090 11.910 1277.270 ;
        RECT 9.130 1274.490 10.310 1275.670 ;
        RECT 10.730 1274.490 11.910 1275.670 ;
        RECT 9.130 1096.090 10.310 1097.270 ;
        RECT 10.730 1096.090 11.910 1097.270 ;
        RECT 9.130 1094.490 10.310 1095.670 ;
        RECT 10.730 1094.490 11.910 1095.670 ;
        RECT 189.130 3523.010 190.310 3524.190 ;
        RECT 190.730 3523.010 191.910 3524.190 ;
        RECT 189.130 3521.410 190.310 3522.590 ;
        RECT 190.730 3521.410 191.910 3522.590 ;
        RECT 189.130 3436.090 190.310 3437.270 ;
        RECT 190.730 3436.090 191.910 3437.270 ;
        RECT 189.130 3434.490 190.310 3435.670 ;
        RECT 190.730 3434.490 191.910 3435.670 ;
        RECT 189.130 3256.090 190.310 3257.270 ;
        RECT 190.730 3256.090 191.910 3257.270 ;
        RECT 189.130 3254.490 190.310 3255.670 ;
        RECT 190.730 3254.490 191.910 3255.670 ;
        RECT 189.130 3076.090 190.310 3077.270 ;
        RECT 190.730 3076.090 191.910 3077.270 ;
        RECT 189.130 3074.490 190.310 3075.670 ;
        RECT 190.730 3074.490 191.910 3075.670 ;
        RECT 189.130 2896.090 190.310 2897.270 ;
        RECT 190.730 2896.090 191.910 2897.270 ;
        RECT 189.130 2894.490 190.310 2895.670 ;
        RECT 190.730 2894.490 191.910 2895.670 ;
        RECT 189.130 2716.090 190.310 2717.270 ;
        RECT 190.730 2716.090 191.910 2717.270 ;
        RECT 189.130 2714.490 190.310 2715.670 ;
        RECT 190.730 2714.490 191.910 2715.670 ;
        RECT 189.130 2536.090 190.310 2537.270 ;
        RECT 190.730 2536.090 191.910 2537.270 ;
        RECT 189.130 2534.490 190.310 2535.670 ;
        RECT 190.730 2534.490 191.910 2535.670 ;
        RECT 189.130 2356.090 190.310 2357.270 ;
        RECT 190.730 2356.090 191.910 2357.270 ;
        RECT 189.130 2354.490 190.310 2355.670 ;
        RECT 190.730 2354.490 191.910 2355.670 ;
        RECT 189.130 2176.090 190.310 2177.270 ;
        RECT 190.730 2176.090 191.910 2177.270 ;
        RECT 189.130 2174.490 190.310 2175.670 ;
        RECT 190.730 2174.490 191.910 2175.670 ;
        RECT 189.130 1996.090 190.310 1997.270 ;
        RECT 190.730 1996.090 191.910 1997.270 ;
        RECT 189.130 1994.490 190.310 1995.670 ;
        RECT 190.730 1994.490 191.910 1995.670 ;
        RECT 189.130 1816.090 190.310 1817.270 ;
        RECT 190.730 1816.090 191.910 1817.270 ;
        RECT 189.130 1814.490 190.310 1815.670 ;
        RECT 190.730 1814.490 191.910 1815.670 ;
        RECT 189.130 1636.090 190.310 1637.270 ;
        RECT 190.730 1636.090 191.910 1637.270 ;
        RECT 189.130 1634.490 190.310 1635.670 ;
        RECT 190.730 1634.490 191.910 1635.670 ;
        RECT 189.130 1456.090 190.310 1457.270 ;
        RECT 190.730 1456.090 191.910 1457.270 ;
        RECT 189.130 1454.490 190.310 1455.670 ;
        RECT 190.730 1454.490 191.910 1455.670 ;
        RECT 189.130 1276.090 190.310 1277.270 ;
        RECT 190.730 1276.090 191.910 1277.270 ;
        RECT 189.130 1274.490 190.310 1275.670 ;
        RECT 190.730 1274.490 191.910 1275.670 ;
        RECT 189.130 1096.090 190.310 1097.270 ;
        RECT 190.730 1096.090 191.910 1097.270 ;
        RECT 189.130 1094.490 190.310 1095.670 ;
        RECT 190.730 1094.490 191.910 1095.670 ;
        RECT 369.130 3523.010 370.310 3524.190 ;
        RECT 370.730 3523.010 371.910 3524.190 ;
        RECT 369.130 3521.410 370.310 3522.590 ;
        RECT 370.730 3521.410 371.910 3522.590 ;
        RECT 369.130 3436.090 370.310 3437.270 ;
        RECT 370.730 3436.090 371.910 3437.270 ;
        RECT 369.130 3434.490 370.310 3435.670 ;
        RECT 370.730 3434.490 371.910 3435.670 ;
        RECT 369.130 3256.090 370.310 3257.270 ;
        RECT 370.730 3256.090 371.910 3257.270 ;
        RECT 369.130 3254.490 370.310 3255.670 ;
        RECT 370.730 3254.490 371.910 3255.670 ;
        RECT 369.130 3076.090 370.310 3077.270 ;
        RECT 370.730 3076.090 371.910 3077.270 ;
        RECT 369.130 3074.490 370.310 3075.670 ;
        RECT 370.730 3074.490 371.910 3075.670 ;
        RECT 369.130 2896.090 370.310 2897.270 ;
        RECT 370.730 2896.090 371.910 2897.270 ;
        RECT 369.130 2894.490 370.310 2895.670 ;
        RECT 370.730 2894.490 371.910 2895.670 ;
        RECT 369.130 2716.090 370.310 2717.270 ;
        RECT 370.730 2716.090 371.910 2717.270 ;
        RECT 369.130 2714.490 370.310 2715.670 ;
        RECT 370.730 2714.490 371.910 2715.670 ;
        RECT 369.130 2536.090 370.310 2537.270 ;
        RECT 370.730 2536.090 371.910 2537.270 ;
        RECT 369.130 2534.490 370.310 2535.670 ;
        RECT 370.730 2534.490 371.910 2535.670 ;
        RECT 369.130 2356.090 370.310 2357.270 ;
        RECT 370.730 2356.090 371.910 2357.270 ;
        RECT 369.130 2354.490 370.310 2355.670 ;
        RECT 370.730 2354.490 371.910 2355.670 ;
        RECT 369.130 2176.090 370.310 2177.270 ;
        RECT 370.730 2176.090 371.910 2177.270 ;
        RECT 369.130 2174.490 370.310 2175.670 ;
        RECT 370.730 2174.490 371.910 2175.670 ;
        RECT 369.130 1996.090 370.310 1997.270 ;
        RECT 370.730 1996.090 371.910 1997.270 ;
        RECT 369.130 1994.490 370.310 1995.670 ;
        RECT 370.730 1994.490 371.910 1995.670 ;
        RECT 369.130 1816.090 370.310 1817.270 ;
        RECT 370.730 1816.090 371.910 1817.270 ;
        RECT 369.130 1814.490 370.310 1815.670 ;
        RECT 370.730 1814.490 371.910 1815.670 ;
        RECT 369.130 1636.090 370.310 1637.270 ;
        RECT 370.730 1636.090 371.910 1637.270 ;
        RECT 369.130 1634.490 370.310 1635.670 ;
        RECT 370.730 1634.490 371.910 1635.670 ;
        RECT 369.130 1456.090 370.310 1457.270 ;
        RECT 370.730 1456.090 371.910 1457.270 ;
        RECT 369.130 1454.490 370.310 1455.670 ;
        RECT 370.730 1454.490 371.910 1455.670 ;
        RECT 369.130 1276.090 370.310 1277.270 ;
        RECT 370.730 1276.090 371.910 1277.270 ;
        RECT 369.130 1274.490 370.310 1275.670 ;
        RECT 370.730 1274.490 371.910 1275.670 ;
        RECT 369.130 1096.090 370.310 1097.270 ;
        RECT 370.730 1096.090 371.910 1097.270 ;
        RECT 369.130 1094.490 370.310 1095.670 ;
        RECT 370.730 1094.490 371.910 1095.670 ;
        RECT 549.130 3523.010 550.310 3524.190 ;
        RECT 550.730 3523.010 551.910 3524.190 ;
        RECT 549.130 3521.410 550.310 3522.590 ;
        RECT 550.730 3521.410 551.910 3522.590 ;
        RECT 549.130 3436.090 550.310 3437.270 ;
        RECT 550.730 3436.090 551.910 3437.270 ;
        RECT 549.130 3434.490 550.310 3435.670 ;
        RECT 550.730 3434.490 551.910 3435.670 ;
        RECT 549.130 3256.090 550.310 3257.270 ;
        RECT 550.730 3256.090 551.910 3257.270 ;
        RECT 549.130 3254.490 550.310 3255.670 ;
        RECT 550.730 3254.490 551.910 3255.670 ;
        RECT 549.130 3076.090 550.310 3077.270 ;
        RECT 550.730 3076.090 551.910 3077.270 ;
        RECT 549.130 3074.490 550.310 3075.670 ;
        RECT 550.730 3074.490 551.910 3075.670 ;
        RECT 549.130 2896.090 550.310 2897.270 ;
        RECT 550.730 2896.090 551.910 2897.270 ;
        RECT 549.130 2894.490 550.310 2895.670 ;
        RECT 550.730 2894.490 551.910 2895.670 ;
        RECT 549.130 2716.090 550.310 2717.270 ;
        RECT 550.730 2716.090 551.910 2717.270 ;
        RECT 549.130 2714.490 550.310 2715.670 ;
        RECT 550.730 2714.490 551.910 2715.670 ;
        RECT 549.130 2536.090 550.310 2537.270 ;
        RECT 550.730 2536.090 551.910 2537.270 ;
        RECT 549.130 2534.490 550.310 2535.670 ;
        RECT 550.730 2534.490 551.910 2535.670 ;
        RECT 549.130 2356.090 550.310 2357.270 ;
        RECT 550.730 2356.090 551.910 2357.270 ;
        RECT 549.130 2354.490 550.310 2355.670 ;
        RECT 550.730 2354.490 551.910 2355.670 ;
        RECT 549.130 2176.090 550.310 2177.270 ;
        RECT 550.730 2176.090 551.910 2177.270 ;
        RECT 549.130 2174.490 550.310 2175.670 ;
        RECT 550.730 2174.490 551.910 2175.670 ;
        RECT 549.130 1996.090 550.310 1997.270 ;
        RECT 550.730 1996.090 551.910 1997.270 ;
        RECT 549.130 1994.490 550.310 1995.670 ;
        RECT 550.730 1994.490 551.910 1995.670 ;
        RECT 549.130 1816.090 550.310 1817.270 ;
        RECT 550.730 1816.090 551.910 1817.270 ;
        RECT 549.130 1814.490 550.310 1815.670 ;
        RECT 550.730 1814.490 551.910 1815.670 ;
        RECT 549.130 1636.090 550.310 1637.270 ;
        RECT 550.730 1636.090 551.910 1637.270 ;
        RECT 549.130 1634.490 550.310 1635.670 ;
        RECT 550.730 1634.490 551.910 1635.670 ;
        RECT 549.130 1456.090 550.310 1457.270 ;
        RECT 550.730 1456.090 551.910 1457.270 ;
        RECT 549.130 1454.490 550.310 1455.670 ;
        RECT 550.730 1454.490 551.910 1455.670 ;
        RECT 549.130 1276.090 550.310 1277.270 ;
        RECT 550.730 1276.090 551.910 1277.270 ;
        RECT 549.130 1274.490 550.310 1275.670 ;
        RECT 550.730 1274.490 551.910 1275.670 ;
        RECT 549.130 1096.090 550.310 1097.270 ;
        RECT 550.730 1096.090 551.910 1097.270 ;
        RECT 549.130 1094.490 550.310 1095.670 ;
        RECT 550.730 1094.490 551.910 1095.670 ;
        RECT 729.130 3523.010 730.310 3524.190 ;
        RECT 730.730 3523.010 731.910 3524.190 ;
        RECT 729.130 3521.410 730.310 3522.590 ;
        RECT 730.730 3521.410 731.910 3522.590 ;
        RECT 729.130 3436.090 730.310 3437.270 ;
        RECT 730.730 3436.090 731.910 3437.270 ;
        RECT 729.130 3434.490 730.310 3435.670 ;
        RECT 730.730 3434.490 731.910 3435.670 ;
        RECT 729.130 3256.090 730.310 3257.270 ;
        RECT 730.730 3256.090 731.910 3257.270 ;
        RECT 729.130 3254.490 730.310 3255.670 ;
        RECT 730.730 3254.490 731.910 3255.670 ;
        RECT 729.130 3076.090 730.310 3077.270 ;
        RECT 730.730 3076.090 731.910 3077.270 ;
        RECT 729.130 3074.490 730.310 3075.670 ;
        RECT 730.730 3074.490 731.910 3075.670 ;
        RECT 729.130 2896.090 730.310 2897.270 ;
        RECT 730.730 2896.090 731.910 2897.270 ;
        RECT 729.130 2894.490 730.310 2895.670 ;
        RECT 730.730 2894.490 731.910 2895.670 ;
        RECT 729.130 2716.090 730.310 2717.270 ;
        RECT 730.730 2716.090 731.910 2717.270 ;
        RECT 729.130 2714.490 730.310 2715.670 ;
        RECT 730.730 2714.490 731.910 2715.670 ;
        RECT 729.130 2536.090 730.310 2537.270 ;
        RECT 730.730 2536.090 731.910 2537.270 ;
        RECT 729.130 2534.490 730.310 2535.670 ;
        RECT 730.730 2534.490 731.910 2535.670 ;
        RECT 729.130 2356.090 730.310 2357.270 ;
        RECT 730.730 2356.090 731.910 2357.270 ;
        RECT 729.130 2354.490 730.310 2355.670 ;
        RECT 730.730 2354.490 731.910 2355.670 ;
        RECT 729.130 2176.090 730.310 2177.270 ;
        RECT 730.730 2176.090 731.910 2177.270 ;
        RECT 729.130 2174.490 730.310 2175.670 ;
        RECT 730.730 2174.490 731.910 2175.670 ;
        RECT 729.130 1996.090 730.310 1997.270 ;
        RECT 730.730 1996.090 731.910 1997.270 ;
        RECT 729.130 1994.490 730.310 1995.670 ;
        RECT 730.730 1994.490 731.910 1995.670 ;
        RECT 729.130 1816.090 730.310 1817.270 ;
        RECT 730.730 1816.090 731.910 1817.270 ;
        RECT 729.130 1814.490 730.310 1815.670 ;
        RECT 730.730 1814.490 731.910 1815.670 ;
        RECT 729.130 1636.090 730.310 1637.270 ;
        RECT 730.730 1636.090 731.910 1637.270 ;
        RECT 729.130 1634.490 730.310 1635.670 ;
        RECT 730.730 1634.490 731.910 1635.670 ;
        RECT 729.130 1456.090 730.310 1457.270 ;
        RECT 730.730 1456.090 731.910 1457.270 ;
        RECT 729.130 1454.490 730.310 1455.670 ;
        RECT 730.730 1454.490 731.910 1455.670 ;
        RECT 729.130 1276.090 730.310 1277.270 ;
        RECT 730.730 1276.090 731.910 1277.270 ;
        RECT 729.130 1274.490 730.310 1275.670 ;
        RECT 730.730 1274.490 731.910 1275.670 ;
        RECT 729.130 1096.090 730.310 1097.270 ;
        RECT 730.730 1096.090 731.910 1097.270 ;
        RECT 729.130 1094.490 730.310 1095.670 ;
        RECT 730.730 1094.490 731.910 1095.670 ;
        RECT 909.130 3523.010 910.310 3524.190 ;
        RECT 910.730 3523.010 911.910 3524.190 ;
        RECT 909.130 3521.410 910.310 3522.590 ;
        RECT 910.730 3521.410 911.910 3522.590 ;
        RECT 909.130 3436.090 910.310 3437.270 ;
        RECT 910.730 3436.090 911.910 3437.270 ;
        RECT 909.130 3434.490 910.310 3435.670 ;
        RECT 910.730 3434.490 911.910 3435.670 ;
        RECT 909.130 3256.090 910.310 3257.270 ;
        RECT 910.730 3256.090 911.910 3257.270 ;
        RECT 909.130 3254.490 910.310 3255.670 ;
        RECT 910.730 3254.490 911.910 3255.670 ;
        RECT 909.130 3076.090 910.310 3077.270 ;
        RECT 910.730 3076.090 911.910 3077.270 ;
        RECT 909.130 3074.490 910.310 3075.670 ;
        RECT 910.730 3074.490 911.910 3075.670 ;
        RECT 909.130 2896.090 910.310 2897.270 ;
        RECT 910.730 2896.090 911.910 2897.270 ;
        RECT 909.130 2894.490 910.310 2895.670 ;
        RECT 910.730 2894.490 911.910 2895.670 ;
        RECT 909.130 2716.090 910.310 2717.270 ;
        RECT 910.730 2716.090 911.910 2717.270 ;
        RECT 909.130 2714.490 910.310 2715.670 ;
        RECT 910.730 2714.490 911.910 2715.670 ;
        RECT 909.130 2536.090 910.310 2537.270 ;
        RECT 910.730 2536.090 911.910 2537.270 ;
        RECT 909.130 2534.490 910.310 2535.670 ;
        RECT 910.730 2534.490 911.910 2535.670 ;
        RECT 909.130 2356.090 910.310 2357.270 ;
        RECT 910.730 2356.090 911.910 2357.270 ;
        RECT 909.130 2354.490 910.310 2355.670 ;
        RECT 910.730 2354.490 911.910 2355.670 ;
        RECT 909.130 2176.090 910.310 2177.270 ;
        RECT 910.730 2176.090 911.910 2177.270 ;
        RECT 909.130 2174.490 910.310 2175.670 ;
        RECT 910.730 2174.490 911.910 2175.670 ;
        RECT 909.130 1996.090 910.310 1997.270 ;
        RECT 910.730 1996.090 911.910 1997.270 ;
        RECT 909.130 1994.490 910.310 1995.670 ;
        RECT 910.730 1994.490 911.910 1995.670 ;
        RECT 909.130 1816.090 910.310 1817.270 ;
        RECT 910.730 1816.090 911.910 1817.270 ;
        RECT 909.130 1814.490 910.310 1815.670 ;
        RECT 910.730 1814.490 911.910 1815.670 ;
        RECT 909.130 1636.090 910.310 1637.270 ;
        RECT 910.730 1636.090 911.910 1637.270 ;
        RECT 909.130 1634.490 910.310 1635.670 ;
        RECT 910.730 1634.490 911.910 1635.670 ;
        RECT 909.130 1456.090 910.310 1457.270 ;
        RECT 910.730 1456.090 911.910 1457.270 ;
        RECT 909.130 1454.490 910.310 1455.670 ;
        RECT 910.730 1454.490 911.910 1455.670 ;
        RECT 909.130 1276.090 910.310 1277.270 ;
        RECT 910.730 1276.090 911.910 1277.270 ;
        RECT 909.130 1274.490 910.310 1275.670 ;
        RECT 910.730 1274.490 911.910 1275.670 ;
        RECT 909.130 1096.090 910.310 1097.270 ;
        RECT 910.730 1096.090 911.910 1097.270 ;
        RECT 909.130 1094.490 910.310 1095.670 ;
        RECT 910.730 1094.490 911.910 1095.670 ;
        RECT 1089.130 3523.010 1090.310 3524.190 ;
        RECT 1090.730 3523.010 1091.910 3524.190 ;
        RECT 1089.130 3521.410 1090.310 3522.590 ;
        RECT 1090.730 3521.410 1091.910 3522.590 ;
        RECT 1089.130 3436.090 1090.310 3437.270 ;
        RECT 1090.730 3436.090 1091.910 3437.270 ;
        RECT 1089.130 3434.490 1090.310 3435.670 ;
        RECT 1090.730 3434.490 1091.910 3435.670 ;
        RECT 1089.130 3256.090 1090.310 3257.270 ;
        RECT 1090.730 3256.090 1091.910 3257.270 ;
        RECT 1089.130 3254.490 1090.310 3255.670 ;
        RECT 1090.730 3254.490 1091.910 3255.670 ;
        RECT 1089.130 3076.090 1090.310 3077.270 ;
        RECT 1090.730 3076.090 1091.910 3077.270 ;
        RECT 1089.130 3074.490 1090.310 3075.670 ;
        RECT 1090.730 3074.490 1091.910 3075.670 ;
        RECT 1089.130 2896.090 1090.310 2897.270 ;
        RECT 1090.730 2896.090 1091.910 2897.270 ;
        RECT 1089.130 2894.490 1090.310 2895.670 ;
        RECT 1090.730 2894.490 1091.910 2895.670 ;
        RECT 1089.130 2716.090 1090.310 2717.270 ;
        RECT 1090.730 2716.090 1091.910 2717.270 ;
        RECT 1089.130 2714.490 1090.310 2715.670 ;
        RECT 1090.730 2714.490 1091.910 2715.670 ;
        RECT 1089.130 2536.090 1090.310 2537.270 ;
        RECT 1090.730 2536.090 1091.910 2537.270 ;
        RECT 1089.130 2534.490 1090.310 2535.670 ;
        RECT 1090.730 2534.490 1091.910 2535.670 ;
        RECT 1089.130 2356.090 1090.310 2357.270 ;
        RECT 1090.730 2356.090 1091.910 2357.270 ;
        RECT 1089.130 2354.490 1090.310 2355.670 ;
        RECT 1090.730 2354.490 1091.910 2355.670 ;
        RECT 1089.130 2176.090 1090.310 2177.270 ;
        RECT 1090.730 2176.090 1091.910 2177.270 ;
        RECT 1089.130 2174.490 1090.310 2175.670 ;
        RECT 1090.730 2174.490 1091.910 2175.670 ;
        RECT 1089.130 1996.090 1090.310 1997.270 ;
        RECT 1090.730 1996.090 1091.910 1997.270 ;
        RECT 1089.130 1994.490 1090.310 1995.670 ;
        RECT 1090.730 1994.490 1091.910 1995.670 ;
        RECT 1089.130 1816.090 1090.310 1817.270 ;
        RECT 1090.730 1816.090 1091.910 1817.270 ;
        RECT 1089.130 1814.490 1090.310 1815.670 ;
        RECT 1090.730 1814.490 1091.910 1815.670 ;
        RECT 1089.130 1636.090 1090.310 1637.270 ;
        RECT 1090.730 1636.090 1091.910 1637.270 ;
        RECT 1089.130 1634.490 1090.310 1635.670 ;
        RECT 1090.730 1634.490 1091.910 1635.670 ;
        RECT 1089.130 1456.090 1090.310 1457.270 ;
        RECT 1090.730 1456.090 1091.910 1457.270 ;
        RECT 1089.130 1454.490 1090.310 1455.670 ;
        RECT 1090.730 1454.490 1091.910 1455.670 ;
        RECT 1089.130 1276.090 1090.310 1277.270 ;
        RECT 1090.730 1276.090 1091.910 1277.270 ;
        RECT 1089.130 1274.490 1090.310 1275.670 ;
        RECT 1090.730 1274.490 1091.910 1275.670 ;
        RECT 1089.130 1096.090 1090.310 1097.270 ;
        RECT 1090.730 1096.090 1091.910 1097.270 ;
        RECT 1089.130 1094.490 1090.310 1095.670 ;
        RECT 1090.730 1094.490 1091.910 1095.670 ;
        RECT 1269.130 3523.010 1270.310 3524.190 ;
        RECT 1270.730 3523.010 1271.910 3524.190 ;
        RECT 1269.130 3521.410 1270.310 3522.590 ;
        RECT 1270.730 3521.410 1271.910 3522.590 ;
        RECT 1269.130 3436.090 1270.310 3437.270 ;
        RECT 1270.730 3436.090 1271.910 3437.270 ;
        RECT 1269.130 3434.490 1270.310 3435.670 ;
        RECT 1270.730 3434.490 1271.910 3435.670 ;
        RECT 1269.130 3256.090 1270.310 3257.270 ;
        RECT 1270.730 3256.090 1271.910 3257.270 ;
        RECT 1269.130 3254.490 1270.310 3255.670 ;
        RECT 1270.730 3254.490 1271.910 3255.670 ;
        RECT 1269.130 3076.090 1270.310 3077.270 ;
        RECT 1270.730 3076.090 1271.910 3077.270 ;
        RECT 1269.130 3074.490 1270.310 3075.670 ;
        RECT 1270.730 3074.490 1271.910 3075.670 ;
        RECT 1269.130 2896.090 1270.310 2897.270 ;
        RECT 1270.730 2896.090 1271.910 2897.270 ;
        RECT 1269.130 2894.490 1270.310 2895.670 ;
        RECT 1270.730 2894.490 1271.910 2895.670 ;
        RECT 1269.130 2716.090 1270.310 2717.270 ;
        RECT 1270.730 2716.090 1271.910 2717.270 ;
        RECT 1269.130 2714.490 1270.310 2715.670 ;
        RECT 1270.730 2714.490 1271.910 2715.670 ;
        RECT 1269.130 2536.090 1270.310 2537.270 ;
        RECT 1270.730 2536.090 1271.910 2537.270 ;
        RECT 1269.130 2534.490 1270.310 2535.670 ;
        RECT 1270.730 2534.490 1271.910 2535.670 ;
        RECT 1269.130 2356.090 1270.310 2357.270 ;
        RECT 1270.730 2356.090 1271.910 2357.270 ;
        RECT 1269.130 2354.490 1270.310 2355.670 ;
        RECT 1270.730 2354.490 1271.910 2355.670 ;
        RECT 1269.130 2176.090 1270.310 2177.270 ;
        RECT 1270.730 2176.090 1271.910 2177.270 ;
        RECT 1269.130 2174.490 1270.310 2175.670 ;
        RECT 1270.730 2174.490 1271.910 2175.670 ;
        RECT 1269.130 1996.090 1270.310 1997.270 ;
        RECT 1270.730 1996.090 1271.910 1997.270 ;
        RECT 1269.130 1994.490 1270.310 1995.670 ;
        RECT 1270.730 1994.490 1271.910 1995.670 ;
        RECT 1269.130 1816.090 1270.310 1817.270 ;
        RECT 1270.730 1816.090 1271.910 1817.270 ;
        RECT 1269.130 1814.490 1270.310 1815.670 ;
        RECT 1270.730 1814.490 1271.910 1815.670 ;
        RECT 1269.130 1636.090 1270.310 1637.270 ;
        RECT 1270.730 1636.090 1271.910 1637.270 ;
        RECT 1269.130 1634.490 1270.310 1635.670 ;
        RECT 1270.730 1634.490 1271.910 1635.670 ;
        RECT 1269.130 1456.090 1270.310 1457.270 ;
        RECT 1270.730 1456.090 1271.910 1457.270 ;
        RECT 1269.130 1454.490 1270.310 1455.670 ;
        RECT 1270.730 1454.490 1271.910 1455.670 ;
        RECT 1269.130 1276.090 1270.310 1277.270 ;
        RECT 1270.730 1276.090 1271.910 1277.270 ;
        RECT 1269.130 1274.490 1270.310 1275.670 ;
        RECT 1270.730 1274.490 1271.910 1275.670 ;
        RECT 1269.130 1096.090 1270.310 1097.270 ;
        RECT 1270.730 1096.090 1271.910 1097.270 ;
        RECT 1269.130 1094.490 1270.310 1095.670 ;
        RECT 1270.730 1094.490 1271.910 1095.670 ;
        RECT 9.130 916.090 10.310 917.270 ;
        RECT 10.730 916.090 11.910 917.270 ;
        RECT 9.130 914.490 10.310 915.670 ;
        RECT 10.730 914.490 11.910 915.670 ;
        RECT 9.130 736.090 10.310 737.270 ;
        RECT 10.730 736.090 11.910 737.270 ;
        RECT 9.130 734.490 10.310 735.670 ;
        RECT 10.730 734.490 11.910 735.670 ;
        RECT 9.130 556.090 10.310 557.270 ;
        RECT 10.730 556.090 11.910 557.270 ;
        RECT 9.130 554.490 10.310 555.670 ;
        RECT 10.730 554.490 11.910 555.670 ;
        RECT 221.250 916.090 222.430 917.270 ;
        RECT 221.250 914.490 222.430 915.670 ;
        RECT 221.250 736.090 222.430 737.270 ;
        RECT 221.250 734.490 222.430 735.670 ;
        RECT 221.250 556.090 222.430 557.270 ;
        RECT 221.250 554.490 222.430 555.670 ;
        RECT 374.850 916.090 376.030 917.270 ;
        RECT 374.850 914.490 376.030 915.670 ;
        RECT 374.850 736.090 376.030 737.270 ;
        RECT 374.850 734.490 376.030 735.670 ;
        RECT 374.850 556.090 376.030 557.270 ;
        RECT 374.850 554.490 376.030 555.670 ;
        RECT 528.450 916.090 529.630 917.270 ;
        RECT 528.450 914.490 529.630 915.670 ;
        RECT 528.450 736.090 529.630 737.270 ;
        RECT 528.450 734.490 529.630 735.670 ;
        RECT 528.450 556.090 529.630 557.270 ;
        RECT 528.450 554.490 529.630 555.670 ;
        RECT 682.050 916.090 683.230 917.270 ;
        RECT 682.050 914.490 683.230 915.670 ;
        RECT 682.050 736.090 683.230 737.270 ;
        RECT 682.050 734.490 683.230 735.670 ;
        RECT 682.050 556.090 683.230 557.270 ;
        RECT 682.050 554.490 683.230 555.670 ;
        RECT 835.650 916.090 836.830 917.270 ;
        RECT 835.650 914.490 836.830 915.670 ;
        RECT 835.650 736.090 836.830 737.270 ;
        RECT 835.650 734.490 836.830 735.670 ;
        RECT 835.650 556.090 836.830 557.270 ;
        RECT 835.650 554.490 836.830 555.670 ;
        RECT 989.250 916.090 990.430 917.270 ;
        RECT 989.250 914.490 990.430 915.670 ;
        RECT 989.250 736.090 990.430 737.270 ;
        RECT 989.250 734.490 990.430 735.670 ;
        RECT 989.250 556.090 990.430 557.270 ;
        RECT 989.250 554.490 990.430 555.670 ;
        RECT 1269.130 916.090 1270.310 917.270 ;
        RECT 1270.730 916.090 1271.910 917.270 ;
        RECT 1269.130 914.490 1270.310 915.670 ;
        RECT 1270.730 914.490 1271.910 915.670 ;
        RECT 1269.130 736.090 1270.310 737.270 ;
        RECT 1270.730 736.090 1271.910 737.270 ;
        RECT 1269.130 734.490 1270.310 735.670 ;
        RECT 1270.730 734.490 1271.910 735.670 ;
        RECT 1269.130 556.090 1270.310 557.270 ;
        RECT 1270.730 556.090 1271.910 557.270 ;
        RECT 1269.130 554.490 1270.310 555.670 ;
        RECT 1270.730 554.490 1271.910 555.670 ;
        RECT 9.130 376.090 10.310 377.270 ;
        RECT 10.730 376.090 11.910 377.270 ;
        RECT 9.130 374.490 10.310 375.670 ;
        RECT 10.730 374.490 11.910 375.670 ;
        RECT 9.130 196.090 10.310 197.270 ;
        RECT 10.730 196.090 11.910 197.270 ;
        RECT 9.130 194.490 10.310 195.670 ;
        RECT 10.730 194.490 11.910 195.670 ;
        RECT 9.130 16.090 10.310 17.270 ;
        RECT 10.730 16.090 11.910 17.270 ;
        RECT 9.130 14.490 10.310 15.670 ;
        RECT 10.730 14.490 11.910 15.670 ;
        RECT 9.130 -2.910 10.310 -1.730 ;
        RECT 10.730 -2.910 11.910 -1.730 ;
        RECT 9.130 -4.510 10.310 -3.330 ;
        RECT 10.730 -4.510 11.910 -3.330 ;
        RECT 189.130 376.090 190.310 377.270 ;
        RECT 190.730 376.090 191.910 377.270 ;
        RECT 189.130 374.490 190.310 375.670 ;
        RECT 190.730 374.490 191.910 375.670 ;
        RECT 189.130 196.090 190.310 197.270 ;
        RECT 190.730 196.090 191.910 197.270 ;
        RECT 189.130 194.490 190.310 195.670 ;
        RECT 190.730 194.490 191.910 195.670 ;
        RECT 189.130 16.090 190.310 17.270 ;
        RECT 190.730 16.090 191.910 17.270 ;
        RECT 189.130 14.490 190.310 15.670 ;
        RECT 190.730 14.490 191.910 15.670 ;
        RECT 189.130 -2.910 190.310 -1.730 ;
        RECT 190.730 -2.910 191.910 -1.730 ;
        RECT 189.130 -4.510 190.310 -3.330 ;
        RECT 190.730 -4.510 191.910 -3.330 ;
        RECT 369.130 376.090 370.310 377.270 ;
        RECT 370.730 376.090 371.910 377.270 ;
        RECT 369.130 374.490 370.310 375.670 ;
        RECT 370.730 374.490 371.910 375.670 ;
        RECT 369.130 196.090 370.310 197.270 ;
        RECT 370.730 196.090 371.910 197.270 ;
        RECT 369.130 194.490 370.310 195.670 ;
        RECT 370.730 194.490 371.910 195.670 ;
        RECT 369.130 16.090 370.310 17.270 ;
        RECT 370.730 16.090 371.910 17.270 ;
        RECT 369.130 14.490 370.310 15.670 ;
        RECT 370.730 14.490 371.910 15.670 ;
        RECT 369.130 -2.910 370.310 -1.730 ;
        RECT 370.730 -2.910 371.910 -1.730 ;
        RECT 369.130 -4.510 370.310 -3.330 ;
        RECT 370.730 -4.510 371.910 -3.330 ;
        RECT 549.130 376.090 550.310 377.270 ;
        RECT 550.730 376.090 551.910 377.270 ;
        RECT 549.130 374.490 550.310 375.670 ;
        RECT 550.730 374.490 551.910 375.670 ;
        RECT 549.130 196.090 550.310 197.270 ;
        RECT 550.730 196.090 551.910 197.270 ;
        RECT 549.130 194.490 550.310 195.670 ;
        RECT 550.730 194.490 551.910 195.670 ;
        RECT 549.130 16.090 550.310 17.270 ;
        RECT 550.730 16.090 551.910 17.270 ;
        RECT 549.130 14.490 550.310 15.670 ;
        RECT 550.730 14.490 551.910 15.670 ;
        RECT 549.130 -2.910 550.310 -1.730 ;
        RECT 550.730 -2.910 551.910 -1.730 ;
        RECT 549.130 -4.510 550.310 -3.330 ;
        RECT 550.730 -4.510 551.910 -3.330 ;
        RECT 729.130 376.090 730.310 377.270 ;
        RECT 730.730 376.090 731.910 377.270 ;
        RECT 729.130 374.490 730.310 375.670 ;
        RECT 730.730 374.490 731.910 375.670 ;
        RECT 729.130 196.090 730.310 197.270 ;
        RECT 730.730 196.090 731.910 197.270 ;
        RECT 729.130 194.490 730.310 195.670 ;
        RECT 730.730 194.490 731.910 195.670 ;
        RECT 729.130 16.090 730.310 17.270 ;
        RECT 730.730 16.090 731.910 17.270 ;
        RECT 729.130 14.490 730.310 15.670 ;
        RECT 730.730 14.490 731.910 15.670 ;
        RECT 729.130 -2.910 730.310 -1.730 ;
        RECT 730.730 -2.910 731.910 -1.730 ;
        RECT 729.130 -4.510 730.310 -3.330 ;
        RECT 730.730 -4.510 731.910 -3.330 ;
        RECT 909.130 376.090 910.310 377.270 ;
        RECT 910.730 376.090 911.910 377.270 ;
        RECT 909.130 374.490 910.310 375.670 ;
        RECT 910.730 374.490 911.910 375.670 ;
        RECT 909.130 196.090 910.310 197.270 ;
        RECT 910.730 196.090 911.910 197.270 ;
        RECT 909.130 194.490 910.310 195.670 ;
        RECT 910.730 194.490 911.910 195.670 ;
        RECT 909.130 16.090 910.310 17.270 ;
        RECT 910.730 16.090 911.910 17.270 ;
        RECT 909.130 14.490 910.310 15.670 ;
        RECT 910.730 14.490 911.910 15.670 ;
        RECT 909.130 -2.910 910.310 -1.730 ;
        RECT 910.730 -2.910 911.910 -1.730 ;
        RECT 909.130 -4.510 910.310 -3.330 ;
        RECT 910.730 -4.510 911.910 -3.330 ;
        RECT 1089.130 376.090 1090.310 377.270 ;
        RECT 1090.730 376.090 1091.910 377.270 ;
        RECT 1089.130 374.490 1090.310 375.670 ;
        RECT 1090.730 374.490 1091.910 375.670 ;
        RECT 1089.130 196.090 1090.310 197.270 ;
        RECT 1090.730 196.090 1091.910 197.270 ;
        RECT 1089.130 194.490 1090.310 195.670 ;
        RECT 1090.730 194.490 1091.910 195.670 ;
        RECT 1089.130 16.090 1090.310 17.270 ;
        RECT 1090.730 16.090 1091.910 17.270 ;
        RECT 1089.130 14.490 1090.310 15.670 ;
        RECT 1090.730 14.490 1091.910 15.670 ;
        RECT 1089.130 -2.910 1090.310 -1.730 ;
        RECT 1090.730 -2.910 1091.910 -1.730 ;
        RECT 1089.130 -4.510 1090.310 -3.330 ;
        RECT 1090.730 -4.510 1091.910 -3.330 ;
        RECT 1269.130 376.090 1270.310 377.270 ;
        RECT 1270.730 376.090 1271.910 377.270 ;
        RECT 1269.130 374.490 1270.310 375.670 ;
        RECT 1270.730 374.490 1271.910 375.670 ;
        RECT 1269.130 196.090 1270.310 197.270 ;
        RECT 1270.730 196.090 1271.910 197.270 ;
        RECT 1269.130 194.490 1270.310 195.670 ;
        RECT 1270.730 194.490 1271.910 195.670 ;
        RECT 1269.130 16.090 1270.310 17.270 ;
        RECT 1270.730 16.090 1271.910 17.270 ;
        RECT 1269.130 14.490 1270.310 15.670 ;
        RECT 1270.730 14.490 1271.910 15.670 ;
        RECT 1269.130 -2.910 1270.310 -1.730 ;
        RECT 1270.730 -2.910 1271.910 -1.730 ;
        RECT 1269.130 -4.510 1270.310 -3.330 ;
        RECT 1270.730 -4.510 1271.910 -3.330 ;
        RECT 1449.130 3523.010 1450.310 3524.190 ;
        RECT 1450.730 3523.010 1451.910 3524.190 ;
        RECT 1449.130 3521.410 1450.310 3522.590 ;
        RECT 1450.730 3521.410 1451.910 3522.590 ;
        RECT 1449.130 3436.090 1450.310 3437.270 ;
        RECT 1450.730 3436.090 1451.910 3437.270 ;
        RECT 1449.130 3434.490 1450.310 3435.670 ;
        RECT 1450.730 3434.490 1451.910 3435.670 ;
        RECT 1449.130 3256.090 1450.310 3257.270 ;
        RECT 1450.730 3256.090 1451.910 3257.270 ;
        RECT 1449.130 3254.490 1450.310 3255.670 ;
        RECT 1450.730 3254.490 1451.910 3255.670 ;
        RECT 1449.130 3076.090 1450.310 3077.270 ;
        RECT 1450.730 3076.090 1451.910 3077.270 ;
        RECT 1449.130 3074.490 1450.310 3075.670 ;
        RECT 1450.730 3074.490 1451.910 3075.670 ;
        RECT 1449.130 2896.090 1450.310 2897.270 ;
        RECT 1450.730 2896.090 1451.910 2897.270 ;
        RECT 1449.130 2894.490 1450.310 2895.670 ;
        RECT 1450.730 2894.490 1451.910 2895.670 ;
        RECT 1449.130 2716.090 1450.310 2717.270 ;
        RECT 1450.730 2716.090 1451.910 2717.270 ;
        RECT 1449.130 2714.490 1450.310 2715.670 ;
        RECT 1450.730 2714.490 1451.910 2715.670 ;
        RECT 1449.130 2536.090 1450.310 2537.270 ;
        RECT 1450.730 2536.090 1451.910 2537.270 ;
        RECT 1449.130 2534.490 1450.310 2535.670 ;
        RECT 1450.730 2534.490 1451.910 2535.670 ;
        RECT 1449.130 2356.090 1450.310 2357.270 ;
        RECT 1450.730 2356.090 1451.910 2357.270 ;
        RECT 1449.130 2354.490 1450.310 2355.670 ;
        RECT 1450.730 2354.490 1451.910 2355.670 ;
        RECT 1449.130 2176.090 1450.310 2177.270 ;
        RECT 1450.730 2176.090 1451.910 2177.270 ;
        RECT 1449.130 2174.490 1450.310 2175.670 ;
        RECT 1450.730 2174.490 1451.910 2175.670 ;
        RECT 1449.130 1996.090 1450.310 1997.270 ;
        RECT 1450.730 1996.090 1451.910 1997.270 ;
        RECT 1449.130 1994.490 1450.310 1995.670 ;
        RECT 1450.730 1994.490 1451.910 1995.670 ;
        RECT 1449.130 1816.090 1450.310 1817.270 ;
        RECT 1450.730 1816.090 1451.910 1817.270 ;
        RECT 1449.130 1814.490 1450.310 1815.670 ;
        RECT 1450.730 1814.490 1451.910 1815.670 ;
        RECT 1449.130 1636.090 1450.310 1637.270 ;
        RECT 1450.730 1636.090 1451.910 1637.270 ;
        RECT 1449.130 1634.490 1450.310 1635.670 ;
        RECT 1450.730 1634.490 1451.910 1635.670 ;
        RECT 1449.130 1456.090 1450.310 1457.270 ;
        RECT 1450.730 1456.090 1451.910 1457.270 ;
        RECT 1449.130 1454.490 1450.310 1455.670 ;
        RECT 1450.730 1454.490 1451.910 1455.670 ;
        RECT 1449.130 1276.090 1450.310 1277.270 ;
        RECT 1450.730 1276.090 1451.910 1277.270 ;
        RECT 1449.130 1274.490 1450.310 1275.670 ;
        RECT 1450.730 1274.490 1451.910 1275.670 ;
        RECT 1449.130 1096.090 1450.310 1097.270 ;
        RECT 1450.730 1096.090 1451.910 1097.270 ;
        RECT 1449.130 1094.490 1450.310 1095.670 ;
        RECT 1450.730 1094.490 1451.910 1095.670 ;
        RECT 1449.130 916.090 1450.310 917.270 ;
        RECT 1450.730 916.090 1451.910 917.270 ;
        RECT 1449.130 914.490 1450.310 915.670 ;
        RECT 1450.730 914.490 1451.910 915.670 ;
        RECT 1449.130 736.090 1450.310 737.270 ;
        RECT 1450.730 736.090 1451.910 737.270 ;
        RECT 1449.130 734.490 1450.310 735.670 ;
        RECT 1450.730 734.490 1451.910 735.670 ;
        RECT 1449.130 556.090 1450.310 557.270 ;
        RECT 1450.730 556.090 1451.910 557.270 ;
        RECT 1449.130 554.490 1450.310 555.670 ;
        RECT 1450.730 554.490 1451.910 555.670 ;
        RECT 1449.130 376.090 1450.310 377.270 ;
        RECT 1450.730 376.090 1451.910 377.270 ;
        RECT 1449.130 374.490 1450.310 375.670 ;
        RECT 1450.730 374.490 1451.910 375.670 ;
        RECT 1449.130 196.090 1450.310 197.270 ;
        RECT 1450.730 196.090 1451.910 197.270 ;
        RECT 1449.130 194.490 1450.310 195.670 ;
        RECT 1450.730 194.490 1451.910 195.670 ;
        RECT 1449.130 16.090 1450.310 17.270 ;
        RECT 1450.730 16.090 1451.910 17.270 ;
        RECT 1449.130 14.490 1450.310 15.670 ;
        RECT 1450.730 14.490 1451.910 15.670 ;
        RECT 1449.130 -2.910 1450.310 -1.730 ;
        RECT 1450.730 -2.910 1451.910 -1.730 ;
        RECT 1449.130 -4.510 1450.310 -3.330 ;
        RECT 1450.730 -4.510 1451.910 -3.330 ;
        RECT 1629.130 3523.010 1630.310 3524.190 ;
        RECT 1630.730 3523.010 1631.910 3524.190 ;
        RECT 1629.130 3521.410 1630.310 3522.590 ;
        RECT 1630.730 3521.410 1631.910 3522.590 ;
        RECT 1629.130 3436.090 1630.310 3437.270 ;
        RECT 1630.730 3436.090 1631.910 3437.270 ;
        RECT 1629.130 3434.490 1630.310 3435.670 ;
        RECT 1630.730 3434.490 1631.910 3435.670 ;
        RECT 1629.130 3256.090 1630.310 3257.270 ;
        RECT 1630.730 3256.090 1631.910 3257.270 ;
        RECT 1629.130 3254.490 1630.310 3255.670 ;
        RECT 1630.730 3254.490 1631.910 3255.670 ;
        RECT 1629.130 3076.090 1630.310 3077.270 ;
        RECT 1630.730 3076.090 1631.910 3077.270 ;
        RECT 1629.130 3074.490 1630.310 3075.670 ;
        RECT 1630.730 3074.490 1631.910 3075.670 ;
        RECT 1629.130 2896.090 1630.310 2897.270 ;
        RECT 1630.730 2896.090 1631.910 2897.270 ;
        RECT 1629.130 2894.490 1630.310 2895.670 ;
        RECT 1630.730 2894.490 1631.910 2895.670 ;
        RECT 1629.130 2716.090 1630.310 2717.270 ;
        RECT 1630.730 2716.090 1631.910 2717.270 ;
        RECT 1629.130 2714.490 1630.310 2715.670 ;
        RECT 1630.730 2714.490 1631.910 2715.670 ;
        RECT 1629.130 2536.090 1630.310 2537.270 ;
        RECT 1630.730 2536.090 1631.910 2537.270 ;
        RECT 1629.130 2534.490 1630.310 2535.670 ;
        RECT 1630.730 2534.490 1631.910 2535.670 ;
        RECT 1629.130 2356.090 1630.310 2357.270 ;
        RECT 1630.730 2356.090 1631.910 2357.270 ;
        RECT 1629.130 2354.490 1630.310 2355.670 ;
        RECT 1630.730 2354.490 1631.910 2355.670 ;
        RECT 1629.130 2176.090 1630.310 2177.270 ;
        RECT 1630.730 2176.090 1631.910 2177.270 ;
        RECT 1629.130 2174.490 1630.310 2175.670 ;
        RECT 1630.730 2174.490 1631.910 2175.670 ;
        RECT 1629.130 1996.090 1630.310 1997.270 ;
        RECT 1630.730 1996.090 1631.910 1997.270 ;
        RECT 1629.130 1994.490 1630.310 1995.670 ;
        RECT 1630.730 1994.490 1631.910 1995.670 ;
        RECT 1629.130 1816.090 1630.310 1817.270 ;
        RECT 1630.730 1816.090 1631.910 1817.270 ;
        RECT 1629.130 1814.490 1630.310 1815.670 ;
        RECT 1630.730 1814.490 1631.910 1815.670 ;
        RECT 1629.130 1636.090 1630.310 1637.270 ;
        RECT 1630.730 1636.090 1631.910 1637.270 ;
        RECT 1629.130 1634.490 1630.310 1635.670 ;
        RECT 1630.730 1634.490 1631.910 1635.670 ;
        RECT 1629.130 1456.090 1630.310 1457.270 ;
        RECT 1630.730 1456.090 1631.910 1457.270 ;
        RECT 1629.130 1454.490 1630.310 1455.670 ;
        RECT 1630.730 1454.490 1631.910 1455.670 ;
        RECT 1629.130 1276.090 1630.310 1277.270 ;
        RECT 1630.730 1276.090 1631.910 1277.270 ;
        RECT 1629.130 1274.490 1630.310 1275.670 ;
        RECT 1630.730 1274.490 1631.910 1275.670 ;
        RECT 1629.130 1096.090 1630.310 1097.270 ;
        RECT 1630.730 1096.090 1631.910 1097.270 ;
        RECT 1629.130 1094.490 1630.310 1095.670 ;
        RECT 1630.730 1094.490 1631.910 1095.670 ;
        RECT 1629.130 916.090 1630.310 917.270 ;
        RECT 1630.730 916.090 1631.910 917.270 ;
        RECT 1629.130 914.490 1630.310 915.670 ;
        RECT 1630.730 914.490 1631.910 915.670 ;
        RECT 1629.130 736.090 1630.310 737.270 ;
        RECT 1630.730 736.090 1631.910 737.270 ;
        RECT 1629.130 734.490 1630.310 735.670 ;
        RECT 1630.730 734.490 1631.910 735.670 ;
        RECT 1629.130 556.090 1630.310 557.270 ;
        RECT 1630.730 556.090 1631.910 557.270 ;
        RECT 1629.130 554.490 1630.310 555.670 ;
        RECT 1630.730 554.490 1631.910 555.670 ;
        RECT 1629.130 376.090 1630.310 377.270 ;
        RECT 1630.730 376.090 1631.910 377.270 ;
        RECT 1629.130 374.490 1630.310 375.670 ;
        RECT 1630.730 374.490 1631.910 375.670 ;
        RECT 1629.130 196.090 1630.310 197.270 ;
        RECT 1630.730 196.090 1631.910 197.270 ;
        RECT 1629.130 194.490 1630.310 195.670 ;
        RECT 1630.730 194.490 1631.910 195.670 ;
        RECT 1629.130 16.090 1630.310 17.270 ;
        RECT 1630.730 16.090 1631.910 17.270 ;
        RECT 1629.130 14.490 1630.310 15.670 ;
        RECT 1630.730 14.490 1631.910 15.670 ;
        RECT 1629.130 -2.910 1630.310 -1.730 ;
        RECT 1630.730 -2.910 1631.910 -1.730 ;
        RECT 1629.130 -4.510 1630.310 -3.330 ;
        RECT 1630.730 -4.510 1631.910 -3.330 ;
        RECT 1809.130 3523.010 1810.310 3524.190 ;
        RECT 1810.730 3523.010 1811.910 3524.190 ;
        RECT 1809.130 3521.410 1810.310 3522.590 ;
        RECT 1810.730 3521.410 1811.910 3522.590 ;
        RECT 1809.130 3436.090 1810.310 3437.270 ;
        RECT 1810.730 3436.090 1811.910 3437.270 ;
        RECT 1809.130 3434.490 1810.310 3435.670 ;
        RECT 1810.730 3434.490 1811.910 3435.670 ;
        RECT 1809.130 3256.090 1810.310 3257.270 ;
        RECT 1810.730 3256.090 1811.910 3257.270 ;
        RECT 1809.130 3254.490 1810.310 3255.670 ;
        RECT 1810.730 3254.490 1811.910 3255.670 ;
        RECT 1809.130 3076.090 1810.310 3077.270 ;
        RECT 1810.730 3076.090 1811.910 3077.270 ;
        RECT 1809.130 3074.490 1810.310 3075.670 ;
        RECT 1810.730 3074.490 1811.910 3075.670 ;
        RECT 1809.130 2896.090 1810.310 2897.270 ;
        RECT 1810.730 2896.090 1811.910 2897.270 ;
        RECT 1809.130 2894.490 1810.310 2895.670 ;
        RECT 1810.730 2894.490 1811.910 2895.670 ;
        RECT 1809.130 2716.090 1810.310 2717.270 ;
        RECT 1810.730 2716.090 1811.910 2717.270 ;
        RECT 1809.130 2714.490 1810.310 2715.670 ;
        RECT 1810.730 2714.490 1811.910 2715.670 ;
        RECT 1809.130 2536.090 1810.310 2537.270 ;
        RECT 1810.730 2536.090 1811.910 2537.270 ;
        RECT 1809.130 2534.490 1810.310 2535.670 ;
        RECT 1810.730 2534.490 1811.910 2535.670 ;
        RECT 1809.130 2356.090 1810.310 2357.270 ;
        RECT 1810.730 2356.090 1811.910 2357.270 ;
        RECT 1809.130 2354.490 1810.310 2355.670 ;
        RECT 1810.730 2354.490 1811.910 2355.670 ;
        RECT 1809.130 2176.090 1810.310 2177.270 ;
        RECT 1810.730 2176.090 1811.910 2177.270 ;
        RECT 1809.130 2174.490 1810.310 2175.670 ;
        RECT 1810.730 2174.490 1811.910 2175.670 ;
        RECT 1809.130 1996.090 1810.310 1997.270 ;
        RECT 1810.730 1996.090 1811.910 1997.270 ;
        RECT 1809.130 1994.490 1810.310 1995.670 ;
        RECT 1810.730 1994.490 1811.910 1995.670 ;
        RECT 1809.130 1816.090 1810.310 1817.270 ;
        RECT 1810.730 1816.090 1811.910 1817.270 ;
        RECT 1809.130 1814.490 1810.310 1815.670 ;
        RECT 1810.730 1814.490 1811.910 1815.670 ;
        RECT 1809.130 1636.090 1810.310 1637.270 ;
        RECT 1810.730 1636.090 1811.910 1637.270 ;
        RECT 1809.130 1634.490 1810.310 1635.670 ;
        RECT 1810.730 1634.490 1811.910 1635.670 ;
        RECT 1809.130 1456.090 1810.310 1457.270 ;
        RECT 1810.730 1456.090 1811.910 1457.270 ;
        RECT 1809.130 1454.490 1810.310 1455.670 ;
        RECT 1810.730 1454.490 1811.910 1455.670 ;
        RECT 1809.130 1276.090 1810.310 1277.270 ;
        RECT 1810.730 1276.090 1811.910 1277.270 ;
        RECT 1809.130 1274.490 1810.310 1275.670 ;
        RECT 1810.730 1274.490 1811.910 1275.670 ;
        RECT 1809.130 1096.090 1810.310 1097.270 ;
        RECT 1810.730 1096.090 1811.910 1097.270 ;
        RECT 1809.130 1094.490 1810.310 1095.670 ;
        RECT 1810.730 1094.490 1811.910 1095.670 ;
        RECT 1809.130 916.090 1810.310 917.270 ;
        RECT 1810.730 916.090 1811.910 917.270 ;
        RECT 1809.130 914.490 1810.310 915.670 ;
        RECT 1810.730 914.490 1811.910 915.670 ;
        RECT 1809.130 736.090 1810.310 737.270 ;
        RECT 1810.730 736.090 1811.910 737.270 ;
        RECT 1809.130 734.490 1810.310 735.670 ;
        RECT 1810.730 734.490 1811.910 735.670 ;
        RECT 1809.130 556.090 1810.310 557.270 ;
        RECT 1810.730 556.090 1811.910 557.270 ;
        RECT 1809.130 554.490 1810.310 555.670 ;
        RECT 1810.730 554.490 1811.910 555.670 ;
        RECT 1809.130 376.090 1810.310 377.270 ;
        RECT 1810.730 376.090 1811.910 377.270 ;
        RECT 1809.130 374.490 1810.310 375.670 ;
        RECT 1810.730 374.490 1811.910 375.670 ;
        RECT 1809.130 196.090 1810.310 197.270 ;
        RECT 1810.730 196.090 1811.910 197.270 ;
        RECT 1809.130 194.490 1810.310 195.670 ;
        RECT 1810.730 194.490 1811.910 195.670 ;
        RECT 1809.130 16.090 1810.310 17.270 ;
        RECT 1810.730 16.090 1811.910 17.270 ;
        RECT 1809.130 14.490 1810.310 15.670 ;
        RECT 1810.730 14.490 1811.910 15.670 ;
        RECT 1809.130 -2.910 1810.310 -1.730 ;
        RECT 1810.730 -2.910 1811.910 -1.730 ;
        RECT 1809.130 -4.510 1810.310 -3.330 ;
        RECT 1810.730 -4.510 1811.910 -3.330 ;
        RECT 1989.130 3523.010 1990.310 3524.190 ;
        RECT 1990.730 3523.010 1991.910 3524.190 ;
        RECT 1989.130 3521.410 1990.310 3522.590 ;
        RECT 1990.730 3521.410 1991.910 3522.590 ;
        RECT 1989.130 3436.090 1990.310 3437.270 ;
        RECT 1990.730 3436.090 1991.910 3437.270 ;
        RECT 1989.130 3434.490 1990.310 3435.670 ;
        RECT 1990.730 3434.490 1991.910 3435.670 ;
        RECT 1989.130 3256.090 1990.310 3257.270 ;
        RECT 1990.730 3256.090 1991.910 3257.270 ;
        RECT 1989.130 3254.490 1990.310 3255.670 ;
        RECT 1990.730 3254.490 1991.910 3255.670 ;
        RECT 1989.130 3076.090 1990.310 3077.270 ;
        RECT 1990.730 3076.090 1991.910 3077.270 ;
        RECT 1989.130 3074.490 1990.310 3075.670 ;
        RECT 1990.730 3074.490 1991.910 3075.670 ;
        RECT 1989.130 2896.090 1990.310 2897.270 ;
        RECT 1990.730 2896.090 1991.910 2897.270 ;
        RECT 1989.130 2894.490 1990.310 2895.670 ;
        RECT 1990.730 2894.490 1991.910 2895.670 ;
        RECT 1989.130 2716.090 1990.310 2717.270 ;
        RECT 1990.730 2716.090 1991.910 2717.270 ;
        RECT 1989.130 2714.490 1990.310 2715.670 ;
        RECT 1990.730 2714.490 1991.910 2715.670 ;
        RECT 1989.130 2536.090 1990.310 2537.270 ;
        RECT 1990.730 2536.090 1991.910 2537.270 ;
        RECT 1989.130 2534.490 1990.310 2535.670 ;
        RECT 1990.730 2534.490 1991.910 2535.670 ;
        RECT 1989.130 2356.090 1990.310 2357.270 ;
        RECT 1990.730 2356.090 1991.910 2357.270 ;
        RECT 1989.130 2354.490 1990.310 2355.670 ;
        RECT 1990.730 2354.490 1991.910 2355.670 ;
        RECT 1989.130 2176.090 1990.310 2177.270 ;
        RECT 1990.730 2176.090 1991.910 2177.270 ;
        RECT 1989.130 2174.490 1990.310 2175.670 ;
        RECT 1990.730 2174.490 1991.910 2175.670 ;
        RECT 1989.130 1996.090 1990.310 1997.270 ;
        RECT 1990.730 1996.090 1991.910 1997.270 ;
        RECT 1989.130 1994.490 1990.310 1995.670 ;
        RECT 1990.730 1994.490 1991.910 1995.670 ;
        RECT 1989.130 1816.090 1990.310 1817.270 ;
        RECT 1990.730 1816.090 1991.910 1817.270 ;
        RECT 1989.130 1814.490 1990.310 1815.670 ;
        RECT 1990.730 1814.490 1991.910 1815.670 ;
        RECT 1989.130 1636.090 1990.310 1637.270 ;
        RECT 1990.730 1636.090 1991.910 1637.270 ;
        RECT 1989.130 1634.490 1990.310 1635.670 ;
        RECT 1990.730 1634.490 1991.910 1635.670 ;
        RECT 1989.130 1456.090 1990.310 1457.270 ;
        RECT 1990.730 1456.090 1991.910 1457.270 ;
        RECT 1989.130 1454.490 1990.310 1455.670 ;
        RECT 1990.730 1454.490 1991.910 1455.670 ;
        RECT 1989.130 1276.090 1990.310 1277.270 ;
        RECT 1990.730 1276.090 1991.910 1277.270 ;
        RECT 1989.130 1274.490 1990.310 1275.670 ;
        RECT 1990.730 1274.490 1991.910 1275.670 ;
        RECT 1989.130 1096.090 1990.310 1097.270 ;
        RECT 1990.730 1096.090 1991.910 1097.270 ;
        RECT 1989.130 1094.490 1990.310 1095.670 ;
        RECT 1990.730 1094.490 1991.910 1095.670 ;
        RECT 1989.130 916.090 1990.310 917.270 ;
        RECT 1990.730 916.090 1991.910 917.270 ;
        RECT 1989.130 914.490 1990.310 915.670 ;
        RECT 1990.730 914.490 1991.910 915.670 ;
        RECT 1989.130 736.090 1990.310 737.270 ;
        RECT 1990.730 736.090 1991.910 737.270 ;
        RECT 1989.130 734.490 1990.310 735.670 ;
        RECT 1990.730 734.490 1991.910 735.670 ;
        RECT 1989.130 556.090 1990.310 557.270 ;
        RECT 1990.730 556.090 1991.910 557.270 ;
        RECT 1989.130 554.490 1990.310 555.670 ;
        RECT 1990.730 554.490 1991.910 555.670 ;
        RECT 1989.130 376.090 1990.310 377.270 ;
        RECT 1990.730 376.090 1991.910 377.270 ;
        RECT 1989.130 374.490 1990.310 375.670 ;
        RECT 1990.730 374.490 1991.910 375.670 ;
        RECT 1989.130 196.090 1990.310 197.270 ;
        RECT 1990.730 196.090 1991.910 197.270 ;
        RECT 1989.130 194.490 1990.310 195.670 ;
        RECT 1990.730 194.490 1991.910 195.670 ;
        RECT 1989.130 16.090 1990.310 17.270 ;
        RECT 1990.730 16.090 1991.910 17.270 ;
        RECT 1989.130 14.490 1990.310 15.670 ;
        RECT 1990.730 14.490 1991.910 15.670 ;
        RECT 1989.130 -2.910 1990.310 -1.730 ;
        RECT 1990.730 -2.910 1991.910 -1.730 ;
        RECT 1989.130 -4.510 1990.310 -3.330 ;
        RECT 1990.730 -4.510 1991.910 -3.330 ;
        RECT 2169.130 3523.010 2170.310 3524.190 ;
        RECT 2170.730 3523.010 2171.910 3524.190 ;
        RECT 2169.130 3521.410 2170.310 3522.590 ;
        RECT 2170.730 3521.410 2171.910 3522.590 ;
        RECT 2169.130 3436.090 2170.310 3437.270 ;
        RECT 2170.730 3436.090 2171.910 3437.270 ;
        RECT 2169.130 3434.490 2170.310 3435.670 ;
        RECT 2170.730 3434.490 2171.910 3435.670 ;
        RECT 2169.130 3256.090 2170.310 3257.270 ;
        RECT 2170.730 3256.090 2171.910 3257.270 ;
        RECT 2169.130 3254.490 2170.310 3255.670 ;
        RECT 2170.730 3254.490 2171.910 3255.670 ;
        RECT 2169.130 3076.090 2170.310 3077.270 ;
        RECT 2170.730 3076.090 2171.910 3077.270 ;
        RECT 2169.130 3074.490 2170.310 3075.670 ;
        RECT 2170.730 3074.490 2171.910 3075.670 ;
        RECT 2169.130 2896.090 2170.310 2897.270 ;
        RECT 2170.730 2896.090 2171.910 2897.270 ;
        RECT 2169.130 2894.490 2170.310 2895.670 ;
        RECT 2170.730 2894.490 2171.910 2895.670 ;
        RECT 2169.130 2716.090 2170.310 2717.270 ;
        RECT 2170.730 2716.090 2171.910 2717.270 ;
        RECT 2169.130 2714.490 2170.310 2715.670 ;
        RECT 2170.730 2714.490 2171.910 2715.670 ;
        RECT 2169.130 2536.090 2170.310 2537.270 ;
        RECT 2170.730 2536.090 2171.910 2537.270 ;
        RECT 2169.130 2534.490 2170.310 2535.670 ;
        RECT 2170.730 2534.490 2171.910 2535.670 ;
        RECT 2169.130 2356.090 2170.310 2357.270 ;
        RECT 2170.730 2356.090 2171.910 2357.270 ;
        RECT 2169.130 2354.490 2170.310 2355.670 ;
        RECT 2170.730 2354.490 2171.910 2355.670 ;
        RECT 2169.130 2176.090 2170.310 2177.270 ;
        RECT 2170.730 2176.090 2171.910 2177.270 ;
        RECT 2169.130 2174.490 2170.310 2175.670 ;
        RECT 2170.730 2174.490 2171.910 2175.670 ;
        RECT 2169.130 1996.090 2170.310 1997.270 ;
        RECT 2170.730 1996.090 2171.910 1997.270 ;
        RECT 2169.130 1994.490 2170.310 1995.670 ;
        RECT 2170.730 1994.490 2171.910 1995.670 ;
        RECT 2169.130 1816.090 2170.310 1817.270 ;
        RECT 2170.730 1816.090 2171.910 1817.270 ;
        RECT 2169.130 1814.490 2170.310 1815.670 ;
        RECT 2170.730 1814.490 2171.910 1815.670 ;
        RECT 2169.130 1636.090 2170.310 1637.270 ;
        RECT 2170.730 1636.090 2171.910 1637.270 ;
        RECT 2169.130 1634.490 2170.310 1635.670 ;
        RECT 2170.730 1634.490 2171.910 1635.670 ;
        RECT 2169.130 1456.090 2170.310 1457.270 ;
        RECT 2170.730 1456.090 2171.910 1457.270 ;
        RECT 2169.130 1454.490 2170.310 1455.670 ;
        RECT 2170.730 1454.490 2171.910 1455.670 ;
        RECT 2169.130 1276.090 2170.310 1277.270 ;
        RECT 2170.730 1276.090 2171.910 1277.270 ;
        RECT 2169.130 1274.490 2170.310 1275.670 ;
        RECT 2170.730 1274.490 2171.910 1275.670 ;
        RECT 2169.130 1096.090 2170.310 1097.270 ;
        RECT 2170.730 1096.090 2171.910 1097.270 ;
        RECT 2169.130 1094.490 2170.310 1095.670 ;
        RECT 2170.730 1094.490 2171.910 1095.670 ;
        RECT 2169.130 916.090 2170.310 917.270 ;
        RECT 2170.730 916.090 2171.910 917.270 ;
        RECT 2169.130 914.490 2170.310 915.670 ;
        RECT 2170.730 914.490 2171.910 915.670 ;
        RECT 2169.130 736.090 2170.310 737.270 ;
        RECT 2170.730 736.090 2171.910 737.270 ;
        RECT 2169.130 734.490 2170.310 735.670 ;
        RECT 2170.730 734.490 2171.910 735.670 ;
        RECT 2169.130 556.090 2170.310 557.270 ;
        RECT 2170.730 556.090 2171.910 557.270 ;
        RECT 2169.130 554.490 2170.310 555.670 ;
        RECT 2170.730 554.490 2171.910 555.670 ;
        RECT 2169.130 376.090 2170.310 377.270 ;
        RECT 2170.730 376.090 2171.910 377.270 ;
        RECT 2169.130 374.490 2170.310 375.670 ;
        RECT 2170.730 374.490 2171.910 375.670 ;
        RECT 2169.130 196.090 2170.310 197.270 ;
        RECT 2170.730 196.090 2171.910 197.270 ;
        RECT 2169.130 194.490 2170.310 195.670 ;
        RECT 2170.730 194.490 2171.910 195.670 ;
        RECT 2169.130 16.090 2170.310 17.270 ;
        RECT 2170.730 16.090 2171.910 17.270 ;
        RECT 2169.130 14.490 2170.310 15.670 ;
        RECT 2170.730 14.490 2171.910 15.670 ;
        RECT 2169.130 -2.910 2170.310 -1.730 ;
        RECT 2170.730 -2.910 2171.910 -1.730 ;
        RECT 2169.130 -4.510 2170.310 -3.330 ;
        RECT 2170.730 -4.510 2171.910 -3.330 ;
        RECT 2349.130 3523.010 2350.310 3524.190 ;
        RECT 2350.730 3523.010 2351.910 3524.190 ;
        RECT 2349.130 3521.410 2350.310 3522.590 ;
        RECT 2350.730 3521.410 2351.910 3522.590 ;
        RECT 2349.130 3436.090 2350.310 3437.270 ;
        RECT 2350.730 3436.090 2351.910 3437.270 ;
        RECT 2349.130 3434.490 2350.310 3435.670 ;
        RECT 2350.730 3434.490 2351.910 3435.670 ;
        RECT 2349.130 3256.090 2350.310 3257.270 ;
        RECT 2350.730 3256.090 2351.910 3257.270 ;
        RECT 2349.130 3254.490 2350.310 3255.670 ;
        RECT 2350.730 3254.490 2351.910 3255.670 ;
        RECT 2349.130 3076.090 2350.310 3077.270 ;
        RECT 2350.730 3076.090 2351.910 3077.270 ;
        RECT 2349.130 3074.490 2350.310 3075.670 ;
        RECT 2350.730 3074.490 2351.910 3075.670 ;
        RECT 2349.130 2896.090 2350.310 2897.270 ;
        RECT 2350.730 2896.090 2351.910 2897.270 ;
        RECT 2349.130 2894.490 2350.310 2895.670 ;
        RECT 2350.730 2894.490 2351.910 2895.670 ;
        RECT 2349.130 2716.090 2350.310 2717.270 ;
        RECT 2350.730 2716.090 2351.910 2717.270 ;
        RECT 2349.130 2714.490 2350.310 2715.670 ;
        RECT 2350.730 2714.490 2351.910 2715.670 ;
        RECT 2349.130 2536.090 2350.310 2537.270 ;
        RECT 2350.730 2536.090 2351.910 2537.270 ;
        RECT 2349.130 2534.490 2350.310 2535.670 ;
        RECT 2350.730 2534.490 2351.910 2535.670 ;
        RECT 2349.130 2356.090 2350.310 2357.270 ;
        RECT 2350.730 2356.090 2351.910 2357.270 ;
        RECT 2349.130 2354.490 2350.310 2355.670 ;
        RECT 2350.730 2354.490 2351.910 2355.670 ;
        RECT 2349.130 2176.090 2350.310 2177.270 ;
        RECT 2350.730 2176.090 2351.910 2177.270 ;
        RECT 2349.130 2174.490 2350.310 2175.670 ;
        RECT 2350.730 2174.490 2351.910 2175.670 ;
        RECT 2349.130 1996.090 2350.310 1997.270 ;
        RECT 2350.730 1996.090 2351.910 1997.270 ;
        RECT 2349.130 1994.490 2350.310 1995.670 ;
        RECT 2350.730 1994.490 2351.910 1995.670 ;
        RECT 2349.130 1816.090 2350.310 1817.270 ;
        RECT 2350.730 1816.090 2351.910 1817.270 ;
        RECT 2349.130 1814.490 2350.310 1815.670 ;
        RECT 2350.730 1814.490 2351.910 1815.670 ;
        RECT 2349.130 1636.090 2350.310 1637.270 ;
        RECT 2350.730 1636.090 2351.910 1637.270 ;
        RECT 2349.130 1634.490 2350.310 1635.670 ;
        RECT 2350.730 1634.490 2351.910 1635.670 ;
        RECT 2349.130 1456.090 2350.310 1457.270 ;
        RECT 2350.730 1456.090 2351.910 1457.270 ;
        RECT 2349.130 1454.490 2350.310 1455.670 ;
        RECT 2350.730 1454.490 2351.910 1455.670 ;
        RECT 2349.130 1276.090 2350.310 1277.270 ;
        RECT 2350.730 1276.090 2351.910 1277.270 ;
        RECT 2349.130 1274.490 2350.310 1275.670 ;
        RECT 2350.730 1274.490 2351.910 1275.670 ;
        RECT 2349.130 1096.090 2350.310 1097.270 ;
        RECT 2350.730 1096.090 2351.910 1097.270 ;
        RECT 2349.130 1094.490 2350.310 1095.670 ;
        RECT 2350.730 1094.490 2351.910 1095.670 ;
        RECT 2349.130 916.090 2350.310 917.270 ;
        RECT 2350.730 916.090 2351.910 917.270 ;
        RECT 2349.130 914.490 2350.310 915.670 ;
        RECT 2350.730 914.490 2351.910 915.670 ;
        RECT 2349.130 736.090 2350.310 737.270 ;
        RECT 2350.730 736.090 2351.910 737.270 ;
        RECT 2349.130 734.490 2350.310 735.670 ;
        RECT 2350.730 734.490 2351.910 735.670 ;
        RECT 2349.130 556.090 2350.310 557.270 ;
        RECT 2350.730 556.090 2351.910 557.270 ;
        RECT 2349.130 554.490 2350.310 555.670 ;
        RECT 2350.730 554.490 2351.910 555.670 ;
        RECT 2349.130 376.090 2350.310 377.270 ;
        RECT 2350.730 376.090 2351.910 377.270 ;
        RECT 2349.130 374.490 2350.310 375.670 ;
        RECT 2350.730 374.490 2351.910 375.670 ;
        RECT 2349.130 196.090 2350.310 197.270 ;
        RECT 2350.730 196.090 2351.910 197.270 ;
        RECT 2349.130 194.490 2350.310 195.670 ;
        RECT 2350.730 194.490 2351.910 195.670 ;
        RECT 2349.130 16.090 2350.310 17.270 ;
        RECT 2350.730 16.090 2351.910 17.270 ;
        RECT 2349.130 14.490 2350.310 15.670 ;
        RECT 2350.730 14.490 2351.910 15.670 ;
        RECT 2349.130 -2.910 2350.310 -1.730 ;
        RECT 2350.730 -2.910 2351.910 -1.730 ;
        RECT 2349.130 -4.510 2350.310 -3.330 ;
        RECT 2350.730 -4.510 2351.910 -3.330 ;
        RECT 2529.130 3523.010 2530.310 3524.190 ;
        RECT 2530.730 3523.010 2531.910 3524.190 ;
        RECT 2529.130 3521.410 2530.310 3522.590 ;
        RECT 2530.730 3521.410 2531.910 3522.590 ;
        RECT 2529.130 3436.090 2530.310 3437.270 ;
        RECT 2530.730 3436.090 2531.910 3437.270 ;
        RECT 2529.130 3434.490 2530.310 3435.670 ;
        RECT 2530.730 3434.490 2531.910 3435.670 ;
        RECT 2529.130 3256.090 2530.310 3257.270 ;
        RECT 2530.730 3256.090 2531.910 3257.270 ;
        RECT 2529.130 3254.490 2530.310 3255.670 ;
        RECT 2530.730 3254.490 2531.910 3255.670 ;
        RECT 2529.130 3076.090 2530.310 3077.270 ;
        RECT 2530.730 3076.090 2531.910 3077.270 ;
        RECT 2529.130 3074.490 2530.310 3075.670 ;
        RECT 2530.730 3074.490 2531.910 3075.670 ;
        RECT 2529.130 2896.090 2530.310 2897.270 ;
        RECT 2530.730 2896.090 2531.910 2897.270 ;
        RECT 2529.130 2894.490 2530.310 2895.670 ;
        RECT 2530.730 2894.490 2531.910 2895.670 ;
        RECT 2529.130 2716.090 2530.310 2717.270 ;
        RECT 2530.730 2716.090 2531.910 2717.270 ;
        RECT 2529.130 2714.490 2530.310 2715.670 ;
        RECT 2530.730 2714.490 2531.910 2715.670 ;
        RECT 2529.130 2536.090 2530.310 2537.270 ;
        RECT 2530.730 2536.090 2531.910 2537.270 ;
        RECT 2529.130 2534.490 2530.310 2535.670 ;
        RECT 2530.730 2534.490 2531.910 2535.670 ;
        RECT 2529.130 2356.090 2530.310 2357.270 ;
        RECT 2530.730 2356.090 2531.910 2357.270 ;
        RECT 2529.130 2354.490 2530.310 2355.670 ;
        RECT 2530.730 2354.490 2531.910 2355.670 ;
        RECT 2529.130 2176.090 2530.310 2177.270 ;
        RECT 2530.730 2176.090 2531.910 2177.270 ;
        RECT 2529.130 2174.490 2530.310 2175.670 ;
        RECT 2530.730 2174.490 2531.910 2175.670 ;
        RECT 2529.130 1996.090 2530.310 1997.270 ;
        RECT 2530.730 1996.090 2531.910 1997.270 ;
        RECT 2529.130 1994.490 2530.310 1995.670 ;
        RECT 2530.730 1994.490 2531.910 1995.670 ;
        RECT 2529.130 1816.090 2530.310 1817.270 ;
        RECT 2530.730 1816.090 2531.910 1817.270 ;
        RECT 2529.130 1814.490 2530.310 1815.670 ;
        RECT 2530.730 1814.490 2531.910 1815.670 ;
        RECT 2529.130 1636.090 2530.310 1637.270 ;
        RECT 2530.730 1636.090 2531.910 1637.270 ;
        RECT 2529.130 1634.490 2530.310 1635.670 ;
        RECT 2530.730 1634.490 2531.910 1635.670 ;
        RECT 2529.130 1456.090 2530.310 1457.270 ;
        RECT 2530.730 1456.090 2531.910 1457.270 ;
        RECT 2529.130 1454.490 2530.310 1455.670 ;
        RECT 2530.730 1454.490 2531.910 1455.670 ;
        RECT 2529.130 1276.090 2530.310 1277.270 ;
        RECT 2530.730 1276.090 2531.910 1277.270 ;
        RECT 2529.130 1274.490 2530.310 1275.670 ;
        RECT 2530.730 1274.490 2531.910 1275.670 ;
        RECT 2529.130 1096.090 2530.310 1097.270 ;
        RECT 2530.730 1096.090 2531.910 1097.270 ;
        RECT 2529.130 1094.490 2530.310 1095.670 ;
        RECT 2530.730 1094.490 2531.910 1095.670 ;
        RECT 2529.130 916.090 2530.310 917.270 ;
        RECT 2530.730 916.090 2531.910 917.270 ;
        RECT 2529.130 914.490 2530.310 915.670 ;
        RECT 2530.730 914.490 2531.910 915.670 ;
        RECT 2529.130 736.090 2530.310 737.270 ;
        RECT 2530.730 736.090 2531.910 737.270 ;
        RECT 2529.130 734.490 2530.310 735.670 ;
        RECT 2530.730 734.490 2531.910 735.670 ;
        RECT 2529.130 556.090 2530.310 557.270 ;
        RECT 2530.730 556.090 2531.910 557.270 ;
        RECT 2529.130 554.490 2530.310 555.670 ;
        RECT 2530.730 554.490 2531.910 555.670 ;
        RECT 2529.130 376.090 2530.310 377.270 ;
        RECT 2530.730 376.090 2531.910 377.270 ;
        RECT 2529.130 374.490 2530.310 375.670 ;
        RECT 2530.730 374.490 2531.910 375.670 ;
        RECT 2529.130 196.090 2530.310 197.270 ;
        RECT 2530.730 196.090 2531.910 197.270 ;
        RECT 2529.130 194.490 2530.310 195.670 ;
        RECT 2530.730 194.490 2531.910 195.670 ;
        RECT 2529.130 16.090 2530.310 17.270 ;
        RECT 2530.730 16.090 2531.910 17.270 ;
        RECT 2529.130 14.490 2530.310 15.670 ;
        RECT 2530.730 14.490 2531.910 15.670 ;
        RECT 2529.130 -2.910 2530.310 -1.730 ;
        RECT 2530.730 -2.910 2531.910 -1.730 ;
        RECT 2529.130 -4.510 2530.310 -3.330 ;
        RECT 2530.730 -4.510 2531.910 -3.330 ;
        RECT 2709.130 3523.010 2710.310 3524.190 ;
        RECT 2710.730 3523.010 2711.910 3524.190 ;
        RECT 2709.130 3521.410 2710.310 3522.590 ;
        RECT 2710.730 3521.410 2711.910 3522.590 ;
        RECT 2709.130 3436.090 2710.310 3437.270 ;
        RECT 2710.730 3436.090 2711.910 3437.270 ;
        RECT 2709.130 3434.490 2710.310 3435.670 ;
        RECT 2710.730 3434.490 2711.910 3435.670 ;
        RECT 2709.130 3256.090 2710.310 3257.270 ;
        RECT 2710.730 3256.090 2711.910 3257.270 ;
        RECT 2709.130 3254.490 2710.310 3255.670 ;
        RECT 2710.730 3254.490 2711.910 3255.670 ;
        RECT 2709.130 3076.090 2710.310 3077.270 ;
        RECT 2710.730 3076.090 2711.910 3077.270 ;
        RECT 2709.130 3074.490 2710.310 3075.670 ;
        RECT 2710.730 3074.490 2711.910 3075.670 ;
        RECT 2709.130 2896.090 2710.310 2897.270 ;
        RECT 2710.730 2896.090 2711.910 2897.270 ;
        RECT 2709.130 2894.490 2710.310 2895.670 ;
        RECT 2710.730 2894.490 2711.910 2895.670 ;
        RECT 2709.130 2716.090 2710.310 2717.270 ;
        RECT 2710.730 2716.090 2711.910 2717.270 ;
        RECT 2709.130 2714.490 2710.310 2715.670 ;
        RECT 2710.730 2714.490 2711.910 2715.670 ;
        RECT 2709.130 2536.090 2710.310 2537.270 ;
        RECT 2710.730 2536.090 2711.910 2537.270 ;
        RECT 2709.130 2534.490 2710.310 2535.670 ;
        RECT 2710.730 2534.490 2711.910 2535.670 ;
        RECT 2709.130 2356.090 2710.310 2357.270 ;
        RECT 2710.730 2356.090 2711.910 2357.270 ;
        RECT 2709.130 2354.490 2710.310 2355.670 ;
        RECT 2710.730 2354.490 2711.910 2355.670 ;
        RECT 2709.130 2176.090 2710.310 2177.270 ;
        RECT 2710.730 2176.090 2711.910 2177.270 ;
        RECT 2709.130 2174.490 2710.310 2175.670 ;
        RECT 2710.730 2174.490 2711.910 2175.670 ;
        RECT 2709.130 1996.090 2710.310 1997.270 ;
        RECT 2710.730 1996.090 2711.910 1997.270 ;
        RECT 2709.130 1994.490 2710.310 1995.670 ;
        RECT 2710.730 1994.490 2711.910 1995.670 ;
        RECT 2709.130 1816.090 2710.310 1817.270 ;
        RECT 2710.730 1816.090 2711.910 1817.270 ;
        RECT 2709.130 1814.490 2710.310 1815.670 ;
        RECT 2710.730 1814.490 2711.910 1815.670 ;
        RECT 2709.130 1636.090 2710.310 1637.270 ;
        RECT 2710.730 1636.090 2711.910 1637.270 ;
        RECT 2709.130 1634.490 2710.310 1635.670 ;
        RECT 2710.730 1634.490 2711.910 1635.670 ;
        RECT 2709.130 1456.090 2710.310 1457.270 ;
        RECT 2710.730 1456.090 2711.910 1457.270 ;
        RECT 2709.130 1454.490 2710.310 1455.670 ;
        RECT 2710.730 1454.490 2711.910 1455.670 ;
        RECT 2709.130 1276.090 2710.310 1277.270 ;
        RECT 2710.730 1276.090 2711.910 1277.270 ;
        RECT 2709.130 1274.490 2710.310 1275.670 ;
        RECT 2710.730 1274.490 2711.910 1275.670 ;
        RECT 2709.130 1096.090 2710.310 1097.270 ;
        RECT 2710.730 1096.090 2711.910 1097.270 ;
        RECT 2709.130 1094.490 2710.310 1095.670 ;
        RECT 2710.730 1094.490 2711.910 1095.670 ;
        RECT 2709.130 916.090 2710.310 917.270 ;
        RECT 2710.730 916.090 2711.910 917.270 ;
        RECT 2709.130 914.490 2710.310 915.670 ;
        RECT 2710.730 914.490 2711.910 915.670 ;
        RECT 2709.130 736.090 2710.310 737.270 ;
        RECT 2710.730 736.090 2711.910 737.270 ;
        RECT 2709.130 734.490 2710.310 735.670 ;
        RECT 2710.730 734.490 2711.910 735.670 ;
        RECT 2709.130 556.090 2710.310 557.270 ;
        RECT 2710.730 556.090 2711.910 557.270 ;
        RECT 2709.130 554.490 2710.310 555.670 ;
        RECT 2710.730 554.490 2711.910 555.670 ;
        RECT 2709.130 376.090 2710.310 377.270 ;
        RECT 2710.730 376.090 2711.910 377.270 ;
        RECT 2709.130 374.490 2710.310 375.670 ;
        RECT 2710.730 374.490 2711.910 375.670 ;
        RECT 2709.130 196.090 2710.310 197.270 ;
        RECT 2710.730 196.090 2711.910 197.270 ;
        RECT 2709.130 194.490 2710.310 195.670 ;
        RECT 2710.730 194.490 2711.910 195.670 ;
        RECT 2709.130 16.090 2710.310 17.270 ;
        RECT 2710.730 16.090 2711.910 17.270 ;
        RECT 2709.130 14.490 2710.310 15.670 ;
        RECT 2710.730 14.490 2711.910 15.670 ;
        RECT 2709.130 -2.910 2710.310 -1.730 ;
        RECT 2710.730 -2.910 2711.910 -1.730 ;
        RECT 2709.130 -4.510 2710.310 -3.330 ;
        RECT 2710.730 -4.510 2711.910 -3.330 ;
        RECT 2889.130 3523.010 2890.310 3524.190 ;
        RECT 2890.730 3523.010 2891.910 3524.190 ;
        RECT 2889.130 3521.410 2890.310 3522.590 ;
        RECT 2890.730 3521.410 2891.910 3522.590 ;
        RECT 2889.130 3436.090 2890.310 3437.270 ;
        RECT 2890.730 3436.090 2891.910 3437.270 ;
        RECT 2889.130 3434.490 2890.310 3435.670 ;
        RECT 2890.730 3434.490 2891.910 3435.670 ;
        RECT 2889.130 3256.090 2890.310 3257.270 ;
        RECT 2890.730 3256.090 2891.910 3257.270 ;
        RECT 2889.130 3254.490 2890.310 3255.670 ;
        RECT 2890.730 3254.490 2891.910 3255.670 ;
        RECT 2889.130 3076.090 2890.310 3077.270 ;
        RECT 2890.730 3076.090 2891.910 3077.270 ;
        RECT 2889.130 3074.490 2890.310 3075.670 ;
        RECT 2890.730 3074.490 2891.910 3075.670 ;
        RECT 2889.130 2896.090 2890.310 2897.270 ;
        RECT 2890.730 2896.090 2891.910 2897.270 ;
        RECT 2889.130 2894.490 2890.310 2895.670 ;
        RECT 2890.730 2894.490 2891.910 2895.670 ;
        RECT 2889.130 2716.090 2890.310 2717.270 ;
        RECT 2890.730 2716.090 2891.910 2717.270 ;
        RECT 2889.130 2714.490 2890.310 2715.670 ;
        RECT 2890.730 2714.490 2891.910 2715.670 ;
        RECT 2889.130 2536.090 2890.310 2537.270 ;
        RECT 2890.730 2536.090 2891.910 2537.270 ;
        RECT 2889.130 2534.490 2890.310 2535.670 ;
        RECT 2890.730 2534.490 2891.910 2535.670 ;
        RECT 2889.130 2356.090 2890.310 2357.270 ;
        RECT 2890.730 2356.090 2891.910 2357.270 ;
        RECT 2889.130 2354.490 2890.310 2355.670 ;
        RECT 2890.730 2354.490 2891.910 2355.670 ;
        RECT 2889.130 2176.090 2890.310 2177.270 ;
        RECT 2890.730 2176.090 2891.910 2177.270 ;
        RECT 2889.130 2174.490 2890.310 2175.670 ;
        RECT 2890.730 2174.490 2891.910 2175.670 ;
        RECT 2889.130 1996.090 2890.310 1997.270 ;
        RECT 2890.730 1996.090 2891.910 1997.270 ;
        RECT 2889.130 1994.490 2890.310 1995.670 ;
        RECT 2890.730 1994.490 2891.910 1995.670 ;
        RECT 2889.130 1816.090 2890.310 1817.270 ;
        RECT 2890.730 1816.090 2891.910 1817.270 ;
        RECT 2889.130 1814.490 2890.310 1815.670 ;
        RECT 2890.730 1814.490 2891.910 1815.670 ;
        RECT 2889.130 1636.090 2890.310 1637.270 ;
        RECT 2890.730 1636.090 2891.910 1637.270 ;
        RECT 2889.130 1634.490 2890.310 1635.670 ;
        RECT 2890.730 1634.490 2891.910 1635.670 ;
        RECT 2889.130 1456.090 2890.310 1457.270 ;
        RECT 2890.730 1456.090 2891.910 1457.270 ;
        RECT 2889.130 1454.490 2890.310 1455.670 ;
        RECT 2890.730 1454.490 2891.910 1455.670 ;
        RECT 2889.130 1276.090 2890.310 1277.270 ;
        RECT 2890.730 1276.090 2891.910 1277.270 ;
        RECT 2889.130 1274.490 2890.310 1275.670 ;
        RECT 2890.730 1274.490 2891.910 1275.670 ;
        RECT 2889.130 1096.090 2890.310 1097.270 ;
        RECT 2890.730 1096.090 2891.910 1097.270 ;
        RECT 2889.130 1094.490 2890.310 1095.670 ;
        RECT 2890.730 1094.490 2891.910 1095.670 ;
        RECT 2889.130 916.090 2890.310 917.270 ;
        RECT 2890.730 916.090 2891.910 917.270 ;
        RECT 2889.130 914.490 2890.310 915.670 ;
        RECT 2890.730 914.490 2891.910 915.670 ;
        RECT 2889.130 736.090 2890.310 737.270 ;
        RECT 2890.730 736.090 2891.910 737.270 ;
        RECT 2889.130 734.490 2890.310 735.670 ;
        RECT 2890.730 734.490 2891.910 735.670 ;
        RECT 2889.130 556.090 2890.310 557.270 ;
        RECT 2890.730 556.090 2891.910 557.270 ;
        RECT 2889.130 554.490 2890.310 555.670 ;
        RECT 2890.730 554.490 2891.910 555.670 ;
        RECT 2889.130 376.090 2890.310 377.270 ;
        RECT 2890.730 376.090 2891.910 377.270 ;
        RECT 2889.130 374.490 2890.310 375.670 ;
        RECT 2890.730 374.490 2891.910 375.670 ;
        RECT 2889.130 196.090 2890.310 197.270 ;
        RECT 2890.730 196.090 2891.910 197.270 ;
        RECT 2889.130 194.490 2890.310 195.670 ;
        RECT 2890.730 194.490 2891.910 195.670 ;
        RECT 2889.130 16.090 2890.310 17.270 ;
        RECT 2890.730 16.090 2891.910 17.270 ;
        RECT 2889.130 14.490 2890.310 15.670 ;
        RECT 2890.730 14.490 2891.910 15.670 ;
        RECT 2889.130 -2.910 2890.310 -1.730 ;
        RECT 2890.730 -2.910 2891.910 -1.730 ;
        RECT 2889.130 -4.510 2890.310 -3.330 ;
        RECT 2890.730 -4.510 2891.910 -3.330 ;
        RECT 2926.710 3523.010 2927.890 3524.190 ;
        RECT 2928.310 3523.010 2929.490 3524.190 ;
        RECT 2926.710 3521.410 2927.890 3522.590 ;
        RECT 2928.310 3521.410 2929.490 3522.590 ;
        RECT 2926.710 3436.090 2927.890 3437.270 ;
        RECT 2928.310 3436.090 2929.490 3437.270 ;
        RECT 2926.710 3434.490 2927.890 3435.670 ;
        RECT 2928.310 3434.490 2929.490 3435.670 ;
        RECT 2926.710 3256.090 2927.890 3257.270 ;
        RECT 2928.310 3256.090 2929.490 3257.270 ;
        RECT 2926.710 3254.490 2927.890 3255.670 ;
        RECT 2928.310 3254.490 2929.490 3255.670 ;
        RECT 2926.710 3076.090 2927.890 3077.270 ;
        RECT 2928.310 3076.090 2929.490 3077.270 ;
        RECT 2926.710 3074.490 2927.890 3075.670 ;
        RECT 2928.310 3074.490 2929.490 3075.670 ;
        RECT 2926.710 2896.090 2927.890 2897.270 ;
        RECT 2928.310 2896.090 2929.490 2897.270 ;
        RECT 2926.710 2894.490 2927.890 2895.670 ;
        RECT 2928.310 2894.490 2929.490 2895.670 ;
        RECT 2926.710 2716.090 2927.890 2717.270 ;
        RECT 2928.310 2716.090 2929.490 2717.270 ;
        RECT 2926.710 2714.490 2927.890 2715.670 ;
        RECT 2928.310 2714.490 2929.490 2715.670 ;
        RECT 2926.710 2536.090 2927.890 2537.270 ;
        RECT 2928.310 2536.090 2929.490 2537.270 ;
        RECT 2926.710 2534.490 2927.890 2535.670 ;
        RECT 2928.310 2534.490 2929.490 2535.670 ;
        RECT 2926.710 2356.090 2927.890 2357.270 ;
        RECT 2928.310 2356.090 2929.490 2357.270 ;
        RECT 2926.710 2354.490 2927.890 2355.670 ;
        RECT 2928.310 2354.490 2929.490 2355.670 ;
        RECT 2926.710 2176.090 2927.890 2177.270 ;
        RECT 2928.310 2176.090 2929.490 2177.270 ;
        RECT 2926.710 2174.490 2927.890 2175.670 ;
        RECT 2928.310 2174.490 2929.490 2175.670 ;
        RECT 2926.710 1996.090 2927.890 1997.270 ;
        RECT 2928.310 1996.090 2929.490 1997.270 ;
        RECT 2926.710 1994.490 2927.890 1995.670 ;
        RECT 2928.310 1994.490 2929.490 1995.670 ;
        RECT 2926.710 1816.090 2927.890 1817.270 ;
        RECT 2928.310 1816.090 2929.490 1817.270 ;
        RECT 2926.710 1814.490 2927.890 1815.670 ;
        RECT 2928.310 1814.490 2929.490 1815.670 ;
        RECT 2926.710 1636.090 2927.890 1637.270 ;
        RECT 2928.310 1636.090 2929.490 1637.270 ;
        RECT 2926.710 1634.490 2927.890 1635.670 ;
        RECT 2928.310 1634.490 2929.490 1635.670 ;
        RECT 2926.710 1456.090 2927.890 1457.270 ;
        RECT 2928.310 1456.090 2929.490 1457.270 ;
        RECT 2926.710 1454.490 2927.890 1455.670 ;
        RECT 2928.310 1454.490 2929.490 1455.670 ;
        RECT 2926.710 1276.090 2927.890 1277.270 ;
        RECT 2928.310 1276.090 2929.490 1277.270 ;
        RECT 2926.710 1274.490 2927.890 1275.670 ;
        RECT 2928.310 1274.490 2929.490 1275.670 ;
        RECT 2926.710 1096.090 2927.890 1097.270 ;
        RECT 2928.310 1096.090 2929.490 1097.270 ;
        RECT 2926.710 1094.490 2927.890 1095.670 ;
        RECT 2928.310 1094.490 2929.490 1095.670 ;
        RECT 2926.710 916.090 2927.890 917.270 ;
        RECT 2928.310 916.090 2929.490 917.270 ;
        RECT 2926.710 914.490 2927.890 915.670 ;
        RECT 2928.310 914.490 2929.490 915.670 ;
        RECT 2926.710 736.090 2927.890 737.270 ;
        RECT 2928.310 736.090 2929.490 737.270 ;
        RECT 2926.710 734.490 2927.890 735.670 ;
        RECT 2928.310 734.490 2929.490 735.670 ;
        RECT 2926.710 556.090 2927.890 557.270 ;
        RECT 2928.310 556.090 2929.490 557.270 ;
        RECT 2926.710 554.490 2927.890 555.670 ;
        RECT 2928.310 554.490 2929.490 555.670 ;
        RECT 2926.710 376.090 2927.890 377.270 ;
        RECT 2928.310 376.090 2929.490 377.270 ;
        RECT 2926.710 374.490 2927.890 375.670 ;
        RECT 2928.310 374.490 2929.490 375.670 ;
        RECT 2926.710 196.090 2927.890 197.270 ;
        RECT 2928.310 196.090 2929.490 197.270 ;
        RECT 2926.710 194.490 2927.890 195.670 ;
        RECT 2928.310 194.490 2929.490 195.670 ;
        RECT 2926.710 16.090 2927.890 17.270 ;
        RECT 2928.310 16.090 2929.490 17.270 ;
        RECT 2926.710 14.490 2927.890 15.670 ;
        RECT 2928.310 14.490 2929.490 15.670 ;
        RECT 2926.710 -2.910 2927.890 -1.730 ;
        RECT 2928.310 -2.910 2929.490 -1.730 ;
        RECT 2926.710 -4.510 2927.890 -3.330 ;
        RECT 2928.310 -4.510 2929.490 -3.330 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
        RECT -14.830 914.330 2934.450 917.430 ;
        RECT -14.830 734.330 2934.450 737.430 ;
        RECT -14.830 554.330 2934.450 557.430 ;
        RECT -14.830 374.330 2934.450 377.430 ;
        RECT -14.830 194.330 2934.450 197.430 ;
        RECT -14.830 14.330 2934.450 17.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
        RECT 207.570 1010.000 210.670 3538.750 ;
        RECT 387.570 1010.000 390.670 3538.750 ;
        RECT 567.570 1010.000 570.670 3538.750 ;
        RECT 747.570 1010.000 750.670 3538.750 ;
        RECT 927.570 1010.000 930.670 3538.750 ;
        RECT 1107.570 1010.000 1110.670 3538.750 ;
        RECT 207.570 -19.070 210.670 390.000 ;
        RECT 387.570 -19.070 390.670 390.000 ;
        RECT 567.570 -19.070 570.670 390.000 ;
        RECT 747.570 -19.070 750.670 390.000 ;
        RECT 927.570 -19.070 930.670 390.000 ;
        RECT 1107.570 -19.070 1110.670 390.000 ;
        RECT 1287.570 -19.070 1290.670 3538.750 ;
        RECT 1467.570 -19.070 1470.670 3538.750 ;
        RECT 1647.570 -19.070 1650.670 3538.750 ;
        RECT 1827.570 -19.070 1830.670 3538.750 ;
        RECT 2007.570 -19.070 2010.670 3538.750 ;
        RECT 2187.570 -19.070 2190.670 3538.750 ;
        RECT 2367.570 -19.070 2370.670 3538.750 ;
        RECT 2547.570 -19.070 2550.670 3538.750 ;
        RECT 2727.570 -19.070 2730.670 3538.750 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER via4 ;
        RECT -19.470 3532.610 -18.290 3533.790 ;
        RECT -17.870 3532.610 -16.690 3533.790 ;
        RECT -19.470 3531.010 -18.290 3532.190 ;
        RECT -17.870 3531.010 -16.690 3532.190 ;
        RECT -19.470 3454.690 -18.290 3455.870 ;
        RECT -17.870 3454.690 -16.690 3455.870 ;
        RECT -19.470 3453.090 -18.290 3454.270 ;
        RECT -17.870 3453.090 -16.690 3454.270 ;
        RECT -19.470 3274.690 -18.290 3275.870 ;
        RECT -17.870 3274.690 -16.690 3275.870 ;
        RECT -19.470 3273.090 -18.290 3274.270 ;
        RECT -17.870 3273.090 -16.690 3274.270 ;
        RECT -19.470 3094.690 -18.290 3095.870 ;
        RECT -17.870 3094.690 -16.690 3095.870 ;
        RECT -19.470 3093.090 -18.290 3094.270 ;
        RECT -17.870 3093.090 -16.690 3094.270 ;
        RECT -19.470 2914.690 -18.290 2915.870 ;
        RECT -17.870 2914.690 -16.690 2915.870 ;
        RECT -19.470 2913.090 -18.290 2914.270 ;
        RECT -17.870 2913.090 -16.690 2914.270 ;
        RECT -19.470 2734.690 -18.290 2735.870 ;
        RECT -17.870 2734.690 -16.690 2735.870 ;
        RECT -19.470 2733.090 -18.290 2734.270 ;
        RECT -17.870 2733.090 -16.690 2734.270 ;
        RECT -19.470 2554.690 -18.290 2555.870 ;
        RECT -17.870 2554.690 -16.690 2555.870 ;
        RECT -19.470 2553.090 -18.290 2554.270 ;
        RECT -17.870 2553.090 -16.690 2554.270 ;
        RECT -19.470 2374.690 -18.290 2375.870 ;
        RECT -17.870 2374.690 -16.690 2375.870 ;
        RECT -19.470 2373.090 -18.290 2374.270 ;
        RECT -17.870 2373.090 -16.690 2374.270 ;
        RECT -19.470 2194.690 -18.290 2195.870 ;
        RECT -17.870 2194.690 -16.690 2195.870 ;
        RECT -19.470 2193.090 -18.290 2194.270 ;
        RECT -17.870 2193.090 -16.690 2194.270 ;
        RECT -19.470 2014.690 -18.290 2015.870 ;
        RECT -17.870 2014.690 -16.690 2015.870 ;
        RECT -19.470 2013.090 -18.290 2014.270 ;
        RECT -17.870 2013.090 -16.690 2014.270 ;
        RECT -19.470 1834.690 -18.290 1835.870 ;
        RECT -17.870 1834.690 -16.690 1835.870 ;
        RECT -19.470 1833.090 -18.290 1834.270 ;
        RECT -17.870 1833.090 -16.690 1834.270 ;
        RECT -19.470 1654.690 -18.290 1655.870 ;
        RECT -17.870 1654.690 -16.690 1655.870 ;
        RECT -19.470 1653.090 -18.290 1654.270 ;
        RECT -17.870 1653.090 -16.690 1654.270 ;
        RECT -19.470 1474.690 -18.290 1475.870 ;
        RECT -17.870 1474.690 -16.690 1475.870 ;
        RECT -19.470 1473.090 -18.290 1474.270 ;
        RECT -17.870 1473.090 -16.690 1474.270 ;
        RECT -19.470 1294.690 -18.290 1295.870 ;
        RECT -17.870 1294.690 -16.690 1295.870 ;
        RECT -19.470 1293.090 -18.290 1294.270 ;
        RECT -17.870 1293.090 -16.690 1294.270 ;
        RECT -19.470 1114.690 -18.290 1115.870 ;
        RECT -17.870 1114.690 -16.690 1115.870 ;
        RECT -19.470 1113.090 -18.290 1114.270 ;
        RECT -17.870 1113.090 -16.690 1114.270 ;
        RECT -19.470 934.690 -18.290 935.870 ;
        RECT -17.870 934.690 -16.690 935.870 ;
        RECT -19.470 933.090 -18.290 934.270 ;
        RECT -17.870 933.090 -16.690 934.270 ;
        RECT -19.470 754.690 -18.290 755.870 ;
        RECT -17.870 754.690 -16.690 755.870 ;
        RECT -19.470 753.090 -18.290 754.270 ;
        RECT -17.870 753.090 -16.690 754.270 ;
        RECT -19.470 574.690 -18.290 575.870 ;
        RECT -17.870 574.690 -16.690 575.870 ;
        RECT -19.470 573.090 -18.290 574.270 ;
        RECT -17.870 573.090 -16.690 574.270 ;
        RECT -19.470 394.690 -18.290 395.870 ;
        RECT -17.870 394.690 -16.690 395.870 ;
        RECT -19.470 393.090 -18.290 394.270 ;
        RECT -17.870 393.090 -16.690 394.270 ;
        RECT -19.470 214.690 -18.290 215.870 ;
        RECT -17.870 214.690 -16.690 215.870 ;
        RECT -19.470 213.090 -18.290 214.270 ;
        RECT -17.870 213.090 -16.690 214.270 ;
        RECT -19.470 34.690 -18.290 35.870 ;
        RECT -17.870 34.690 -16.690 35.870 ;
        RECT -19.470 33.090 -18.290 34.270 ;
        RECT -17.870 33.090 -16.690 34.270 ;
        RECT -19.470 -12.510 -18.290 -11.330 ;
        RECT -17.870 -12.510 -16.690 -11.330 ;
        RECT -19.470 -14.110 -18.290 -12.930 ;
        RECT -17.870 -14.110 -16.690 -12.930 ;
        RECT 27.730 3532.610 28.910 3533.790 ;
        RECT 29.330 3532.610 30.510 3533.790 ;
        RECT 27.730 3531.010 28.910 3532.190 ;
        RECT 29.330 3531.010 30.510 3532.190 ;
        RECT 27.730 3454.690 28.910 3455.870 ;
        RECT 29.330 3454.690 30.510 3455.870 ;
        RECT 27.730 3453.090 28.910 3454.270 ;
        RECT 29.330 3453.090 30.510 3454.270 ;
        RECT 27.730 3274.690 28.910 3275.870 ;
        RECT 29.330 3274.690 30.510 3275.870 ;
        RECT 27.730 3273.090 28.910 3274.270 ;
        RECT 29.330 3273.090 30.510 3274.270 ;
        RECT 27.730 3094.690 28.910 3095.870 ;
        RECT 29.330 3094.690 30.510 3095.870 ;
        RECT 27.730 3093.090 28.910 3094.270 ;
        RECT 29.330 3093.090 30.510 3094.270 ;
        RECT 27.730 2914.690 28.910 2915.870 ;
        RECT 29.330 2914.690 30.510 2915.870 ;
        RECT 27.730 2913.090 28.910 2914.270 ;
        RECT 29.330 2913.090 30.510 2914.270 ;
        RECT 27.730 2734.690 28.910 2735.870 ;
        RECT 29.330 2734.690 30.510 2735.870 ;
        RECT 27.730 2733.090 28.910 2734.270 ;
        RECT 29.330 2733.090 30.510 2734.270 ;
        RECT 27.730 2554.690 28.910 2555.870 ;
        RECT 29.330 2554.690 30.510 2555.870 ;
        RECT 27.730 2553.090 28.910 2554.270 ;
        RECT 29.330 2553.090 30.510 2554.270 ;
        RECT 27.730 2374.690 28.910 2375.870 ;
        RECT 29.330 2374.690 30.510 2375.870 ;
        RECT 27.730 2373.090 28.910 2374.270 ;
        RECT 29.330 2373.090 30.510 2374.270 ;
        RECT 27.730 2194.690 28.910 2195.870 ;
        RECT 29.330 2194.690 30.510 2195.870 ;
        RECT 27.730 2193.090 28.910 2194.270 ;
        RECT 29.330 2193.090 30.510 2194.270 ;
        RECT 27.730 2014.690 28.910 2015.870 ;
        RECT 29.330 2014.690 30.510 2015.870 ;
        RECT 27.730 2013.090 28.910 2014.270 ;
        RECT 29.330 2013.090 30.510 2014.270 ;
        RECT 27.730 1834.690 28.910 1835.870 ;
        RECT 29.330 1834.690 30.510 1835.870 ;
        RECT 27.730 1833.090 28.910 1834.270 ;
        RECT 29.330 1833.090 30.510 1834.270 ;
        RECT 27.730 1654.690 28.910 1655.870 ;
        RECT 29.330 1654.690 30.510 1655.870 ;
        RECT 27.730 1653.090 28.910 1654.270 ;
        RECT 29.330 1653.090 30.510 1654.270 ;
        RECT 27.730 1474.690 28.910 1475.870 ;
        RECT 29.330 1474.690 30.510 1475.870 ;
        RECT 27.730 1473.090 28.910 1474.270 ;
        RECT 29.330 1473.090 30.510 1474.270 ;
        RECT 27.730 1294.690 28.910 1295.870 ;
        RECT 29.330 1294.690 30.510 1295.870 ;
        RECT 27.730 1293.090 28.910 1294.270 ;
        RECT 29.330 1293.090 30.510 1294.270 ;
        RECT 27.730 1114.690 28.910 1115.870 ;
        RECT 29.330 1114.690 30.510 1115.870 ;
        RECT 27.730 1113.090 28.910 1114.270 ;
        RECT 29.330 1113.090 30.510 1114.270 ;
        RECT 207.730 3532.610 208.910 3533.790 ;
        RECT 209.330 3532.610 210.510 3533.790 ;
        RECT 207.730 3531.010 208.910 3532.190 ;
        RECT 209.330 3531.010 210.510 3532.190 ;
        RECT 207.730 3454.690 208.910 3455.870 ;
        RECT 209.330 3454.690 210.510 3455.870 ;
        RECT 207.730 3453.090 208.910 3454.270 ;
        RECT 209.330 3453.090 210.510 3454.270 ;
        RECT 207.730 3274.690 208.910 3275.870 ;
        RECT 209.330 3274.690 210.510 3275.870 ;
        RECT 207.730 3273.090 208.910 3274.270 ;
        RECT 209.330 3273.090 210.510 3274.270 ;
        RECT 207.730 3094.690 208.910 3095.870 ;
        RECT 209.330 3094.690 210.510 3095.870 ;
        RECT 207.730 3093.090 208.910 3094.270 ;
        RECT 209.330 3093.090 210.510 3094.270 ;
        RECT 207.730 2914.690 208.910 2915.870 ;
        RECT 209.330 2914.690 210.510 2915.870 ;
        RECT 207.730 2913.090 208.910 2914.270 ;
        RECT 209.330 2913.090 210.510 2914.270 ;
        RECT 207.730 2734.690 208.910 2735.870 ;
        RECT 209.330 2734.690 210.510 2735.870 ;
        RECT 207.730 2733.090 208.910 2734.270 ;
        RECT 209.330 2733.090 210.510 2734.270 ;
        RECT 207.730 2554.690 208.910 2555.870 ;
        RECT 209.330 2554.690 210.510 2555.870 ;
        RECT 207.730 2553.090 208.910 2554.270 ;
        RECT 209.330 2553.090 210.510 2554.270 ;
        RECT 207.730 2374.690 208.910 2375.870 ;
        RECT 209.330 2374.690 210.510 2375.870 ;
        RECT 207.730 2373.090 208.910 2374.270 ;
        RECT 209.330 2373.090 210.510 2374.270 ;
        RECT 207.730 2194.690 208.910 2195.870 ;
        RECT 209.330 2194.690 210.510 2195.870 ;
        RECT 207.730 2193.090 208.910 2194.270 ;
        RECT 209.330 2193.090 210.510 2194.270 ;
        RECT 207.730 2014.690 208.910 2015.870 ;
        RECT 209.330 2014.690 210.510 2015.870 ;
        RECT 207.730 2013.090 208.910 2014.270 ;
        RECT 209.330 2013.090 210.510 2014.270 ;
        RECT 207.730 1834.690 208.910 1835.870 ;
        RECT 209.330 1834.690 210.510 1835.870 ;
        RECT 207.730 1833.090 208.910 1834.270 ;
        RECT 209.330 1833.090 210.510 1834.270 ;
        RECT 207.730 1654.690 208.910 1655.870 ;
        RECT 209.330 1654.690 210.510 1655.870 ;
        RECT 207.730 1653.090 208.910 1654.270 ;
        RECT 209.330 1653.090 210.510 1654.270 ;
        RECT 207.730 1474.690 208.910 1475.870 ;
        RECT 209.330 1474.690 210.510 1475.870 ;
        RECT 207.730 1473.090 208.910 1474.270 ;
        RECT 209.330 1473.090 210.510 1474.270 ;
        RECT 207.730 1294.690 208.910 1295.870 ;
        RECT 209.330 1294.690 210.510 1295.870 ;
        RECT 207.730 1293.090 208.910 1294.270 ;
        RECT 209.330 1293.090 210.510 1294.270 ;
        RECT 207.730 1114.690 208.910 1115.870 ;
        RECT 209.330 1114.690 210.510 1115.870 ;
        RECT 207.730 1113.090 208.910 1114.270 ;
        RECT 209.330 1113.090 210.510 1114.270 ;
        RECT 387.730 3532.610 388.910 3533.790 ;
        RECT 389.330 3532.610 390.510 3533.790 ;
        RECT 387.730 3531.010 388.910 3532.190 ;
        RECT 389.330 3531.010 390.510 3532.190 ;
        RECT 387.730 3454.690 388.910 3455.870 ;
        RECT 389.330 3454.690 390.510 3455.870 ;
        RECT 387.730 3453.090 388.910 3454.270 ;
        RECT 389.330 3453.090 390.510 3454.270 ;
        RECT 387.730 3274.690 388.910 3275.870 ;
        RECT 389.330 3274.690 390.510 3275.870 ;
        RECT 387.730 3273.090 388.910 3274.270 ;
        RECT 389.330 3273.090 390.510 3274.270 ;
        RECT 387.730 3094.690 388.910 3095.870 ;
        RECT 389.330 3094.690 390.510 3095.870 ;
        RECT 387.730 3093.090 388.910 3094.270 ;
        RECT 389.330 3093.090 390.510 3094.270 ;
        RECT 387.730 2914.690 388.910 2915.870 ;
        RECT 389.330 2914.690 390.510 2915.870 ;
        RECT 387.730 2913.090 388.910 2914.270 ;
        RECT 389.330 2913.090 390.510 2914.270 ;
        RECT 387.730 2734.690 388.910 2735.870 ;
        RECT 389.330 2734.690 390.510 2735.870 ;
        RECT 387.730 2733.090 388.910 2734.270 ;
        RECT 389.330 2733.090 390.510 2734.270 ;
        RECT 387.730 2554.690 388.910 2555.870 ;
        RECT 389.330 2554.690 390.510 2555.870 ;
        RECT 387.730 2553.090 388.910 2554.270 ;
        RECT 389.330 2553.090 390.510 2554.270 ;
        RECT 387.730 2374.690 388.910 2375.870 ;
        RECT 389.330 2374.690 390.510 2375.870 ;
        RECT 387.730 2373.090 388.910 2374.270 ;
        RECT 389.330 2373.090 390.510 2374.270 ;
        RECT 387.730 2194.690 388.910 2195.870 ;
        RECT 389.330 2194.690 390.510 2195.870 ;
        RECT 387.730 2193.090 388.910 2194.270 ;
        RECT 389.330 2193.090 390.510 2194.270 ;
        RECT 387.730 2014.690 388.910 2015.870 ;
        RECT 389.330 2014.690 390.510 2015.870 ;
        RECT 387.730 2013.090 388.910 2014.270 ;
        RECT 389.330 2013.090 390.510 2014.270 ;
        RECT 387.730 1834.690 388.910 1835.870 ;
        RECT 389.330 1834.690 390.510 1835.870 ;
        RECT 387.730 1833.090 388.910 1834.270 ;
        RECT 389.330 1833.090 390.510 1834.270 ;
        RECT 387.730 1654.690 388.910 1655.870 ;
        RECT 389.330 1654.690 390.510 1655.870 ;
        RECT 387.730 1653.090 388.910 1654.270 ;
        RECT 389.330 1653.090 390.510 1654.270 ;
        RECT 387.730 1474.690 388.910 1475.870 ;
        RECT 389.330 1474.690 390.510 1475.870 ;
        RECT 387.730 1473.090 388.910 1474.270 ;
        RECT 389.330 1473.090 390.510 1474.270 ;
        RECT 387.730 1294.690 388.910 1295.870 ;
        RECT 389.330 1294.690 390.510 1295.870 ;
        RECT 387.730 1293.090 388.910 1294.270 ;
        RECT 389.330 1293.090 390.510 1294.270 ;
        RECT 387.730 1114.690 388.910 1115.870 ;
        RECT 389.330 1114.690 390.510 1115.870 ;
        RECT 387.730 1113.090 388.910 1114.270 ;
        RECT 389.330 1113.090 390.510 1114.270 ;
        RECT 567.730 3532.610 568.910 3533.790 ;
        RECT 569.330 3532.610 570.510 3533.790 ;
        RECT 567.730 3531.010 568.910 3532.190 ;
        RECT 569.330 3531.010 570.510 3532.190 ;
        RECT 567.730 3454.690 568.910 3455.870 ;
        RECT 569.330 3454.690 570.510 3455.870 ;
        RECT 567.730 3453.090 568.910 3454.270 ;
        RECT 569.330 3453.090 570.510 3454.270 ;
        RECT 567.730 3274.690 568.910 3275.870 ;
        RECT 569.330 3274.690 570.510 3275.870 ;
        RECT 567.730 3273.090 568.910 3274.270 ;
        RECT 569.330 3273.090 570.510 3274.270 ;
        RECT 567.730 3094.690 568.910 3095.870 ;
        RECT 569.330 3094.690 570.510 3095.870 ;
        RECT 567.730 3093.090 568.910 3094.270 ;
        RECT 569.330 3093.090 570.510 3094.270 ;
        RECT 567.730 2914.690 568.910 2915.870 ;
        RECT 569.330 2914.690 570.510 2915.870 ;
        RECT 567.730 2913.090 568.910 2914.270 ;
        RECT 569.330 2913.090 570.510 2914.270 ;
        RECT 567.730 2734.690 568.910 2735.870 ;
        RECT 569.330 2734.690 570.510 2735.870 ;
        RECT 567.730 2733.090 568.910 2734.270 ;
        RECT 569.330 2733.090 570.510 2734.270 ;
        RECT 567.730 2554.690 568.910 2555.870 ;
        RECT 569.330 2554.690 570.510 2555.870 ;
        RECT 567.730 2553.090 568.910 2554.270 ;
        RECT 569.330 2553.090 570.510 2554.270 ;
        RECT 567.730 2374.690 568.910 2375.870 ;
        RECT 569.330 2374.690 570.510 2375.870 ;
        RECT 567.730 2373.090 568.910 2374.270 ;
        RECT 569.330 2373.090 570.510 2374.270 ;
        RECT 567.730 2194.690 568.910 2195.870 ;
        RECT 569.330 2194.690 570.510 2195.870 ;
        RECT 567.730 2193.090 568.910 2194.270 ;
        RECT 569.330 2193.090 570.510 2194.270 ;
        RECT 567.730 2014.690 568.910 2015.870 ;
        RECT 569.330 2014.690 570.510 2015.870 ;
        RECT 567.730 2013.090 568.910 2014.270 ;
        RECT 569.330 2013.090 570.510 2014.270 ;
        RECT 567.730 1834.690 568.910 1835.870 ;
        RECT 569.330 1834.690 570.510 1835.870 ;
        RECT 567.730 1833.090 568.910 1834.270 ;
        RECT 569.330 1833.090 570.510 1834.270 ;
        RECT 567.730 1654.690 568.910 1655.870 ;
        RECT 569.330 1654.690 570.510 1655.870 ;
        RECT 567.730 1653.090 568.910 1654.270 ;
        RECT 569.330 1653.090 570.510 1654.270 ;
        RECT 567.730 1474.690 568.910 1475.870 ;
        RECT 569.330 1474.690 570.510 1475.870 ;
        RECT 567.730 1473.090 568.910 1474.270 ;
        RECT 569.330 1473.090 570.510 1474.270 ;
        RECT 567.730 1294.690 568.910 1295.870 ;
        RECT 569.330 1294.690 570.510 1295.870 ;
        RECT 567.730 1293.090 568.910 1294.270 ;
        RECT 569.330 1293.090 570.510 1294.270 ;
        RECT 567.730 1114.690 568.910 1115.870 ;
        RECT 569.330 1114.690 570.510 1115.870 ;
        RECT 567.730 1113.090 568.910 1114.270 ;
        RECT 569.330 1113.090 570.510 1114.270 ;
        RECT 747.730 3532.610 748.910 3533.790 ;
        RECT 749.330 3532.610 750.510 3533.790 ;
        RECT 747.730 3531.010 748.910 3532.190 ;
        RECT 749.330 3531.010 750.510 3532.190 ;
        RECT 747.730 3454.690 748.910 3455.870 ;
        RECT 749.330 3454.690 750.510 3455.870 ;
        RECT 747.730 3453.090 748.910 3454.270 ;
        RECT 749.330 3453.090 750.510 3454.270 ;
        RECT 747.730 3274.690 748.910 3275.870 ;
        RECT 749.330 3274.690 750.510 3275.870 ;
        RECT 747.730 3273.090 748.910 3274.270 ;
        RECT 749.330 3273.090 750.510 3274.270 ;
        RECT 747.730 3094.690 748.910 3095.870 ;
        RECT 749.330 3094.690 750.510 3095.870 ;
        RECT 747.730 3093.090 748.910 3094.270 ;
        RECT 749.330 3093.090 750.510 3094.270 ;
        RECT 747.730 2914.690 748.910 2915.870 ;
        RECT 749.330 2914.690 750.510 2915.870 ;
        RECT 747.730 2913.090 748.910 2914.270 ;
        RECT 749.330 2913.090 750.510 2914.270 ;
        RECT 747.730 2734.690 748.910 2735.870 ;
        RECT 749.330 2734.690 750.510 2735.870 ;
        RECT 747.730 2733.090 748.910 2734.270 ;
        RECT 749.330 2733.090 750.510 2734.270 ;
        RECT 747.730 2554.690 748.910 2555.870 ;
        RECT 749.330 2554.690 750.510 2555.870 ;
        RECT 747.730 2553.090 748.910 2554.270 ;
        RECT 749.330 2553.090 750.510 2554.270 ;
        RECT 747.730 2374.690 748.910 2375.870 ;
        RECT 749.330 2374.690 750.510 2375.870 ;
        RECT 747.730 2373.090 748.910 2374.270 ;
        RECT 749.330 2373.090 750.510 2374.270 ;
        RECT 747.730 2194.690 748.910 2195.870 ;
        RECT 749.330 2194.690 750.510 2195.870 ;
        RECT 747.730 2193.090 748.910 2194.270 ;
        RECT 749.330 2193.090 750.510 2194.270 ;
        RECT 747.730 2014.690 748.910 2015.870 ;
        RECT 749.330 2014.690 750.510 2015.870 ;
        RECT 747.730 2013.090 748.910 2014.270 ;
        RECT 749.330 2013.090 750.510 2014.270 ;
        RECT 747.730 1834.690 748.910 1835.870 ;
        RECT 749.330 1834.690 750.510 1835.870 ;
        RECT 747.730 1833.090 748.910 1834.270 ;
        RECT 749.330 1833.090 750.510 1834.270 ;
        RECT 747.730 1654.690 748.910 1655.870 ;
        RECT 749.330 1654.690 750.510 1655.870 ;
        RECT 747.730 1653.090 748.910 1654.270 ;
        RECT 749.330 1653.090 750.510 1654.270 ;
        RECT 747.730 1474.690 748.910 1475.870 ;
        RECT 749.330 1474.690 750.510 1475.870 ;
        RECT 747.730 1473.090 748.910 1474.270 ;
        RECT 749.330 1473.090 750.510 1474.270 ;
        RECT 747.730 1294.690 748.910 1295.870 ;
        RECT 749.330 1294.690 750.510 1295.870 ;
        RECT 747.730 1293.090 748.910 1294.270 ;
        RECT 749.330 1293.090 750.510 1294.270 ;
        RECT 747.730 1114.690 748.910 1115.870 ;
        RECT 749.330 1114.690 750.510 1115.870 ;
        RECT 747.730 1113.090 748.910 1114.270 ;
        RECT 749.330 1113.090 750.510 1114.270 ;
        RECT 927.730 3532.610 928.910 3533.790 ;
        RECT 929.330 3532.610 930.510 3533.790 ;
        RECT 927.730 3531.010 928.910 3532.190 ;
        RECT 929.330 3531.010 930.510 3532.190 ;
        RECT 927.730 3454.690 928.910 3455.870 ;
        RECT 929.330 3454.690 930.510 3455.870 ;
        RECT 927.730 3453.090 928.910 3454.270 ;
        RECT 929.330 3453.090 930.510 3454.270 ;
        RECT 927.730 3274.690 928.910 3275.870 ;
        RECT 929.330 3274.690 930.510 3275.870 ;
        RECT 927.730 3273.090 928.910 3274.270 ;
        RECT 929.330 3273.090 930.510 3274.270 ;
        RECT 927.730 3094.690 928.910 3095.870 ;
        RECT 929.330 3094.690 930.510 3095.870 ;
        RECT 927.730 3093.090 928.910 3094.270 ;
        RECT 929.330 3093.090 930.510 3094.270 ;
        RECT 927.730 2914.690 928.910 2915.870 ;
        RECT 929.330 2914.690 930.510 2915.870 ;
        RECT 927.730 2913.090 928.910 2914.270 ;
        RECT 929.330 2913.090 930.510 2914.270 ;
        RECT 927.730 2734.690 928.910 2735.870 ;
        RECT 929.330 2734.690 930.510 2735.870 ;
        RECT 927.730 2733.090 928.910 2734.270 ;
        RECT 929.330 2733.090 930.510 2734.270 ;
        RECT 927.730 2554.690 928.910 2555.870 ;
        RECT 929.330 2554.690 930.510 2555.870 ;
        RECT 927.730 2553.090 928.910 2554.270 ;
        RECT 929.330 2553.090 930.510 2554.270 ;
        RECT 927.730 2374.690 928.910 2375.870 ;
        RECT 929.330 2374.690 930.510 2375.870 ;
        RECT 927.730 2373.090 928.910 2374.270 ;
        RECT 929.330 2373.090 930.510 2374.270 ;
        RECT 927.730 2194.690 928.910 2195.870 ;
        RECT 929.330 2194.690 930.510 2195.870 ;
        RECT 927.730 2193.090 928.910 2194.270 ;
        RECT 929.330 2193.090 930.510 2194.270 ;
        RECT 927.730 2014.690 928.910 2015.870 ;
        RECT 929.330 2014.690 930.510 2015.870 ;
        RECT 927.730 2013.090 928.910 2014.270 ;
        RECT 929.330 2013.090 930.510 2014.270 ;
        RECT 927.730 1834.690 928.910 1835.870 ;
        RECT 929.330 1834.690 930.510 1835.870 ;
        RECT 927.730 1833.090 928.910 1834.270 ;
        RECT 929.330 1833.090 930.510 1834.270 ;
        RECT 927.730 1654.690 928.910 1655.870 ;
        RECT 929.330 1654.690 930.510 1655.870 ;
        RECT 927.730 1653.090 928.910 1654.270 ;
        RECT 929.330 1653.090 930.510 1654.270 ;
        RECT 927.730 1474.690 928.910 1475.870 ;
        RECT 929.330 1474.690 930.510 1475.870 ;
        RECT 927.730 1473.090 928.910 1474.270 ;
        RECT 929.330 1473.090 930.510 1474.270 ;
        RECT 927.730 1294.690 928.910 1295.870 ;
        RECT 929.330 1294.690 930.510 1295.870 ;
        RECT 927.730 1293.090 928.910 1294.270 ;
        RECT 929.330 1293.090 930.510 1294.270 ;
        RECT 927.730 1114.690 928.910 1115.870 ;
        RECT 929.330 1114.690 930.510 1115.870 ;
        RECT 927.730 1113.090 928.910 1114.270 ;
        RECT 929.330 1113.090 930.510 1114.270 ;
        RECT 1107.730 3532.610 1108.910 3533.790 ;
        RECT 1109.330 3532.610 1110.510 3533.790 ;
        RECT 1107.730 3531.010 1108.910 3532.190 ;
        RECT 1109.330 3531.010 1110.510 3532.190 ;
        RECT 1107.730 3454.690 1108.910 3455.870 ;
        RECT 1109.330 3454.690 1110.510 3455.870 ;
        RECT 1107.730 3453.090 1108.910 3454.270 ;
        RECT 1109.330 3453.090 1110.510 3454.270 ;
        RECT 1107.730 3274.690 1108.910 3275.870 ;
        RECT 1109.330 3274.690 1110.510 3275.870 ;
        RECT 1107.730 3273.090 1108.910 3274.270 ;
        RECT 1109.330 3273.090 1110.510 3274.270 ;
        RECT 1107.730 3094.690 1108.910 3095.870 ;
        RECT 1109.330 3094.690 1110.510 3095.870 ;
        RECT 1107.730 3093.090 1108.910 3094.270 ;
        RECT 1109.330 3093.090 1110.510 3094.270 ;
        RECT 1107.730 2914.690 1108.910 2915.870 ;
        RECT 1109.330 2914.690 1110.510 2915.870 ;
        RECT 1107.730 2913.090 1108.910 2914.270 ;
        RECT 1109.330 2913.090 1110.510 2914.270 ;
        RECT 1107.730 2734.690 1108.910 2735.870 ;
        RECT 1109.330 2734.690 1110.510 2735.870 ;
        RECT 1107.730 2733.090 1108.910 2734.270 ;
        RECT 1109.330 2733.090 1110.510 2734.270 ;
        RECT 1107.730 2554.690 1108.910 2555.870 ;
        RECT 1109.330 2554.690 1110.510 2555.870 ;
        RECT 1107.730 2553.090 1108.910 2554.270 ;
        RECT 1109.330 2553.090 1110.510 2554.270 ;
        RECT 1107.730 2374.690 1108.910 2375.870 ;
        RECT 1109.330 2374.690 1110.510 2375.870 ;
        RECT 1107.730 2373.090 1108.910 2374.270 ;
        RECT 1109.330 2373.090 1110.510 2374.270 ;
        RECT 1107.730 2194.690 1108.910 2195.870 ;
        RECT 1109.330 2194.690 1110.510 2195.870 ;
        RECT 1107.730 2193.090 1108.910 2194.270 ;
        RECT 1109.330 2193.090 1110.510 2194.270 ;
        RECT 1107.730 2014.690 1108.910 2015.870 ;
        RECT 1109.330 2014.690 1110.510 2015.870 ;
        RECT 1107.730 2013.090 1108.910 2014.270 ;
        RECT 1109.330 2013.090 1110.510 2014.270 ;
        RECT 1107.730 1834.690 1108.910 1835.870 ;
        RECT 1109.330 1834.690 1110.510 1835.870 ;
        RECT 1107.730 1833.090 1108.910 1834.270 ;
        RECT 1109.330 1833.090 1110.510 1834.270 ;
        RECT 1107.730 1654.690 1108.910 1655.870 ;
        RECT 1109.330 1654.690 1110.510 1655.870 ;
        RECT 1107.730 1653.090 1108.910 1654.270 ;
        RECT 1109.330 1653.090 1110.510 1654.270 ;
        RECT 1107.730 1474.690 1108.910 1475.870 ;
        RECT 1109.330 1474.690 1110.510 1475.870 ;
        RECT 1107.730 1473.090 1108.910 1474.270 ;
        RECT 1109.330 1473.090 1110.510 1474.270 ;
        RECT 1107.730 1294.690 1108.910 1295.870 ;
        RECT 1109.330 1294.690 1110.510 1295.870 ;
        RECT 1107.730 1293.090 1108.910 1294.270 ;
        RECT 1109.330 1293.090 1110.510 1294.270 ;
        RECT 1107.730 1114.690 1108.910 1115.870 ;
        RECT 1109.330 1114.690 1110.510 1115.870 ;
        RECT 1107.730 1113.090 1108.910 1114.270 ;
        RECT 1109.330 1113.090 1110.510 1114.270 ;
        RECT 1287.730 3532.610 1288.910 3533.790 ;
        RECT 1289.330 3532.610 1290.510 3533.790 ;
        RECT 1287.730 3531.010 1288.910 3532.190 ;
        RECT 1289.330 3531.010 1290.510 3532.190 ;
        RECT 1287.730 3454.690 1288.910 3455.870 ;
        RECT 1289.330 3454.690 1290.510 3455.870 ;
        RECT 1287.730 3453.090 1288.910 3454.270 ;
        RECT 1289.330 3453.090 1290.510 3454.270 ;
        RECT 1287.730 3274.690 1288.910 3275.870 ;
        RECT 1289.330 3274.690 1290.510 3275.870 ;
        RECT 1287.730 3273.090 1288.910 3274.270 ;
        RECT 1289.330 3273.090 1290.510 3274.270 ;
        RECT 1287.730 3094.690 1288.910 3095.870 ;
        RECT 1289.330 3094.690 1290.510 3095.870 ;
        RECT 1287.730 3093.090 1288.910 3094.270 ;
        RECT 1289.330 3093.090 1290.510 3094.270 ;
        RECT 1287.730 2914.690 1288.910 2915.870 ;
        RECT 1289.330 2914.690 1290.510 2915.870 ;
        RECT 1287.730 2913.090 1288.910 2914.270 ;
        RECT 1289.330 2913.090 1290.510 2914.270 ;
        RECT 1287.730 2734.690 1288.910 2735.870 ;
        RECT 1289.330 2734.690 1290.510 2735.870 ;
        RECT 1287.730 2733.090 1288.910 2734.270 ;
        RECT 1289.330 2733.090 1290.510 2734.270 ;
        RECT 1287.730 2554.690 1288.910 2555.870 ;
        RECT 1289.330 2554.690 1290.510 2555.870 ;
        RECT 1287.730 2553.090 1288.910 2554.270 ;
        RECT 1289.330 2553.090 1290.510 2554.270 ;
        RECT 1287.730 2374.690 1288.910 2375.870 ;
        RECT 1289.330 2374.690 1290.510 2375.870 ;
        RECT 1287.730 2373.090 1288.910 2374.270 ;
        RECT 1289.330 2373.090 1290.510 2374.270 ;
        RECT 1287.730 2194.690 1288.910 2195.870 ;
        RECT 1289.330 2194.690 1290.510 2195.870 ;
        RECT 1287.730 2193.090 1288.910 2194.270 ;
        RECT 1289.330 2193.090 1290.510 2194.270 ;
        RECT 1287.730 2014.690 1288.910 2015.870 ;
        RECT 1289.330 2014.690 1290.510 2015.870 ;
        RECT 1287.730 2013.090 1288.910 2014.270 ;
        RECT 1289.330 2013.090 1290.510 2014.270 ;
        RECT 1287.730 1834.690 1288.910 1835.870 ;
        RECT 1289.330 1834.690 1290.510 1835.870 ;
        RECT 1287.730 1833.090 1288.910 1834.270 ;
        RECT 1289.330 1833.090 1290.510 1834.270 ;
        RECT 1287.730 1654.690 1288.910 1655.870 ;
        RECT 1289.330 1654.690 1290.510 1655.870 ;
        RECT 1287.730 1653.090 1288.910 1654.270 ;
        RECT 1289.330 1653.090 1290.510 1654.270 ;
        RECT 1287.730 1474.690 1288.910 1475.870 ;
        RECT 1289.330 1474.690 1290.510 1475.870 ;
        RECT 1287.730 1473.090 1288.910 1474.270 ;
        RECT 1289.330 1473.090 1290.510 1474.270 ;
        RECT 1287.730 1294.690 1288.910 1295.870 ;
        RECT 1289.330 1294.690 1290.510 1295.870 ;
        RECT 1287.730 1293.090 1288.910 1294.270 ;
        RECT 1289.330 1293.090 1290.510 1294.270 ;
        RECT 1287.730 1114.690 1288.910 1115.870 ;
        RECT 1289.330 1114.690 1290.510 1115.870 ;
        RECT 1287.730 1113.090 1288.910 1114.270 ;
        RECT 1289.330 1113.090 1290.510 1114.270 ;
        RECT 27.730 934.690 28.910 935.870 ;
        RECT 29.330 934.690 30.510 935.870 ;
        RECT 27.730 933.090 28.910 934.270 ;
        RECT 29.330 933.090 30.510 934.270 ;
        RECT 27.730 754.690 28.910 755.870 ;
        RECT 29.330 754.690 30.510 755.870 ;
        RECT 27.730 753.090 28.910 754.270 ;
        RECT 29.330 753.090 30.510 754.270 ;
        RECT 27.730 574.690 28.910 575.870 ;
        RECT 29.330 574.690 30.510 575.870 ;
        RECT 27.730 573.090 28.910 574.270 ;
        RECT 29.330 573.090 30.510 574.270 ;
        RECT 27.730 394.690 28.910 395.870 ;
        RECT 29.330 394.690 30.510 395.870 ;
        RECT 27.730 393.090 28.910 394.270 ;
        RECT 29.330 393.090 30.510 394.270 ;
        RECT 1287.730 934.690 1288.910 935.870 ;
        RECT 1289.330 934.690 1290.510 935.870 ;
        RECT 1287.730 933.090 1288.910 934.270 ;
        RECT 1289.330 933.090 1290.510 934.270 ;
        RECT 1287.730 754.690 1288.910 755.870 ;
        RECT 1289.330 754.690 1290.510 755.870 ;
        RECT 1287.730 753.090 1288.910 754.270 ;
        RECT 1289.330 753.090 1290.510 754.270 ;
        RECT 1287.730 574.690 1288.910 575.870 ;
        RECT 1289.330 574.690 1290.510 575.870 ;
        RECT 1287.730 573.090 1288.910 574.270 ;
        RECT 1289.330 573.090 1290.510 574.270 ;
        RECT 1287.730 394.690 1288.910 395.870 ;
        RECT 1289.330 394.690 1290.510 395.870 ;
        RECT 1287.730 393.090 1288.910 394.270 ;
        RECT 1289.330 393.090 1290.510 394.270 ;
        RECT 27.730 214.690 28.910 215.870 ;
        RECT 29.330 214.690 30.510 215.870 ;
        RECT 27.730 213.090 28.910 214.270 ;
        RECT 29.330 213.090 30.510 214.270 ;
        RECT 27.730 34.690 28.910 35.870 ;
        RECT 29.330 34.690 30.510 35.870 ;
        RECT 27.730 33.090 28.910 34.270 ;
        RECT 29.330 33.090 30.510 34.270 ;
        RECT 27.730 -12.510 28.910 -11.330 ;
        RECT 29.330 -12.510 30.510 -11.330 ;
        RECT 27.730 -14.110 28.910 -12.930 ;
        RECT 29.330 -14.110 30.510 -12.930 ;
        RECT 207.730 214.690 208.910 215.870 ;
        RECT 209.330 214.690 210.510 215.870 ;
        RECT 207.730 213.090 208.910 214.270 ;
        RECT 209.330 213.090 210.510 214.270 ;
        RECT 207.730 34.690 208.910 35.870 ;
        RECT 209.330 34.690 210.510 35.870 ;
        RECT 207.730 33.090 208.910 34.270 ;
        RECT 209.330 33.090 210.510 34.270 ;
        RECT 207.730 -12.510 208.910 -11.330 ;
        RECT 209.330 -12.510 210.510 -11.330 ;
        RECT 207.730 -14.110 208.910 -12.930 ;
        RECT 209.330 -14.110 210.510 -12.930 ;
        RECT 387.730 214.690 388.910 215.870 ;
        RECT 389.330 214.690 390.510 215.870 ;
        RECT 387.730 213.090 388.910 214.270 ;
        RECT 389.330 213.090 390.510 214.270 ;
        RECT 387.730 34.690 388.910 35.870 ;
        RECT 389.330 34.690 390.510 35.870 ;
        RECT 387.730 33.090 388.910 34.270 ;
        RECT 389.330 33.090 390.510 34.270 ;
        RECT 387.730 -12.510 388.910 -11.330 ;
        RECT 389.330 -12.510 390.510 -11.330 ;
        RECT 387.730 -14.110 388.910 -12.930 ;
        RECT 389.330 -14.110 390.510 -12.930 ;
        RECT 567.730 214.690 568.910 215.870 ;
        RECT 569.330 214.690 570.510 215.870 ;
        RECT 567.730 213.090 568.910 214.270 ;
        RECT 569.330 213.090 570.510 214.270 ;
        RECT 567.730 34.690 568.910 35.870 ;
        RECT 569.330 34.690 570.510 35.870 ;
        RECT 567.730 33.090 568.910 34.270 ;
        RECT 569.330 33.090 570.510 34.270 ;
        RECT 567.730 -12.510 568.910 -11.330 ;
        RECT 569.330 -12.510 570.510 -11.330 ;
        RECT 567.730 -14.110 568.910 -12.930 ;
        RECT 569.330 -14.110 570.510 -12.930 ;
        RECT 747.730 214.690 748.910 215.870 ;
        RECT 749.330 214.690 750.510 215.870 ;
        RECT 747.730 213.090 748.910 214.270 ;
        RECT 749.330 213.090 750.510 214.270 ;
        RECT 747.730 34.690 748.910 35.870 ;
        RECT 749.330 34.690 750.510 35.870 ;
        RECT 747.730 33.090 748.910 34.270 ;
        RECT 749.330 33.090 750.510 34.270 ;
        RECT 747.730 -12.510 748.910 -11.330 ;
        RECT 749.330 -12.510 750.510 -11.330 ;
        RECT 747.730 -14.110 748.910 -12.930 ;
        RECT 749.330 -14.110 750.510 -12.930 ;
        RECT 927.730 214.690 928.910 215.870 ;
        RECT 929.330 214.690 930.510 215.870 ;
        RECT 927.730 213.090 928.910 214.270 ;
        RECT 929.330 213.090 930.510 214.270 ;
        RECT 927.730 34.690 928.910 35.870 ;
        RECT 929.330 34.690 930.510 35.870 ;
        RECT 927.730 33.090 928.910 34.270 ;
        RECT 929.330 33.090 930.510 34.270 ;
        RECT 927.730 -12.510 928.910 -11.330 ;
        RECT 929.330 -12.510 930.510 -11.330 ;
        RECT 927.730 -14.110 928.910 -12.930 ;
        RECT 929.330 -14.110 930.510 -12.930 ;
        RECT 1107.730 214.690 1108.910 215.870 ;
        RECT 1109.330 214.690 1110.510 215.870 ;
        RECT 1107.730 213.090 1108.910 214.270 ;
        RECT 1109.330 213.090 1110.510 214.270 ;
        RECT 1107.730 34.690 1108.910 35.870 ;
        RECT 1109.330 34.690 1110.510 35.870 ;
        RECT 1107.730 33.090 1108.910 34.270 ;
        RECT 1109.330 33.090 1110.510 34.270 ;
        RECT 1107.730 -12.510 1108.910 -11.330 ;
        RECT 1109.330 -12.510 1110.510 -11.330 ;
        RECT 1107.730 -14.110 1108.910 -12.930 ;
        RECT 1109.330 -14.110 1110.510 -12.930 ;
        RECT 1287.730 214.690 1288.910 215.870 ;
        RECT 1289.330 214.690 1290.510 215.870 ;
        RECT 1287.730 213.090 1288.910 214.270 ;
        RECT 1289.330 213.090 1290.510 214.270 ;
        RECT 1287.730 34.690 1288.910 35.870 ;
        RECT 1289.330 34.690 1290.510 35.870 ;
        RECT 1287.730 33.090 1288.910 34.270 ;
        RECT 1289.330 33.090 1290.510 34.270 ;
        RECT 1287.730 -12.510 1288.910 -11.330 ;
        RECT 1289.330 -12.510 1290.510 -11.330 ;
        RECT 1287.730 -14.110 1288.910 -12.930 ;
        RECT 1289.330 -14.110 1290.510 -12.930 ;
        RECT 1467.730 3532.610 1468.910 3533.790 ;
        RECT 1469.330 3532.610 1470.510 3533.790 ;
        RECT 1467.730 3531.010 1468.910 3532.190 ;
        RECT 1469.330 3531.010 1470.510 3532.190 ;
        RECT 1467.730 3454.690 1468.910 3455.870 ;
        RECT 1469.330 3454.690 1470.510 3455.870 ;
        RECT 1467.730 3453.090 1468.910 3454.270 ;
        RECT 1469.330 3453.090 1470.510 3454.270 ;
        RECT 1467.730 3274.690 1468.910 3275.870 ;
        RECT 1469.330 3274.690 1470.510 3275.870 ;
        RECT 1467.730 3273.090 1468.910 3274.270 ;
        RECT 1469.330 3273.090 1470.510 3274.270 ;
        RECT 1467.730 3094.690 1468.910 3095.870 ;
        RECT 1469.330 3094.690 1470.510 3095.870 ;
        RECT 1467.730 3093.090 1468.910 3094.270 ;
        RECT 1469.330 3093.090 1470.510 3094.270 ;
        RECT 1467.730 2914.690 1468.910 2915.870 ;
        RECT 1469.330 2914.690 1470.510 2915.870 ;
        RECT 1467.730 2913.090 1468.910 2914.270 ;
        RECT 1469.330 2913.090 1470.510 2914.270 ;
        RECT 1467.730 2734.690 1468.910 2735.870 ;
        RECT 1469.330 2734.690 1470.510 2735.870 ;
        RECT 1467.730 2733.090 1468.910 2734.270 ;
        RECT 1469.330 2733.090 1470.510 2734.270 ;
        RECT 1467.730 2554.690 1468.910 2555.870 ;
        RECT 1469.330 2554.690 1470.510 2555.870 ;
        RECT 1467.730 2553.090 1468.910 2554.270 ;
        RECT 1469.330 2553.090 1470.510 2554.270 ;
        RECT 1467.730 2374.690 1468.910 2375.870 ;
        RECT 1469.330 2374.690 1470.510 2375.870 ;
        RECT 1467.730 2373.090 1468.910 2374.270 ;
        RECT 1469.330 2373.090 1470.510 2374.270 ;
        RECT 1467.730 2194.690 1468.910 2195.870 ;
        RECT 1469.330 2194.690 1470.510 2195.870 ;
        RECT 1467.730 2193.090 1468.910 2194.270 ;
        RECT 1469.330 2193.090 1470.510 2194.270 ;
        RECT 1467.730 2014.690 1468.910 2015.870 ;
        RECT 1469.330 2014.690 1470.510 2015.870 ;
        RECT 1467.730 2013.090 1468.910 2014.270 ;
        RECT 1469.330 2013.090 1470.510 2014.270 ;
        RECT 1467.730 1834.690 1468.910 1835.870 ;
        RECT 1469.330 1834.690 1470.510 1835.870 ;
        RECT 1467.730 1833.090 1468.910 1834.270 ;
        RECT 1469.330 1833.090 1470.510 1834.270 ;
        RECT 1467.730 1654.690 1468.910 1655.870 ;
        RECT 1469.330 1654.690 1470.510 1655.870 ;
        RECT 1467.730 1653.090 1468.910 1654.270 ;
        RECT 1469.330 1653.090 1470.510 1654.270 ;
        RECT 1467.730 1474.690 1468.910 1475.870 ;
        RECT 1469.330 1474.690 1470.510 1475.870 ;
        RECT 1467.730 1473.090 1468.910 1474.270 ;
        RECT 1469.330 1473.090 1470.510 1474.270 ;
        RECT 1467.730 1294.690 1468.910 1295.870 ;
        RECT 1469.330 1294.690 1470.510 1295.870 ;
        RECT 1467.730 1293.090 1468.910 1294.270 ;
        RECT 1469.330 1293.090 1470.510 1294.270 ;
        RECT 1467.730 1114.690 1468.910 1115.870 ;
        RECT 1469.330 1114.690 1470.510 1115.870 ;
        RECT 1467.730 1113.090 1468.910 1114.270 ;
        RECT 1469.330 1113.090 1470.510 1114.270 ;
        RECT 1467.730 934.690 1468.910 935.870 ;
        RECT 1469.330 934.690 1470.510 935.870 ;
        RECT 1467.730 933.090 1468.910 934.270 ;
        RECT 1469.330 933.090 1470.510 934.270 ;
        RECT 1467.730 754.690 1468.910 755.870 ;
        RECT 1469.330 754.690 1470.510 755.870 ;
        RECT 1467.730 753.090 1468.910 754.270 ;
        RECT 1469.330 753.090 1470.510 754.270 ;
        RECT 1467.730 574.690 1468.910 575.870 ;
        RECT 1469.330 574.690 1470.510 575.870 ;
        RECT 1467.730 573.090 1468.910 574.270 ;
        RECT 1469.330 573.090 1470.510 574.270 ;
        RECT 1467.730 394.690 1468.910 395.870 ;
        RECT 1469.330 394.690 1470.510 395.870 ;
        RECT 1467.730 393.090 1468.910 394.270 ;
        RECT 1469.330 393.090 1470.510 394.270 ;
        RECT 1467.730 214.690 1468.910 215.870 ;
        RECT 1469.330 214.690 1470.510 215.870 ;
        RECT 1467.730 213.090 1468.910 214.270 ;
        RECT 1469.330 213.090 1470.510 214.270 ;
        RECT 1467.730 34.690 1468.910 35.870 ;
        RECT 1469.330 34.690 1470.510 35.870 ;
        RECT 1467.730 33.090 1468.910 34.270 ;
        RECT 1469.330 33.090 1470.510 34.270 ;
        RECT 1467.730 -12.510 1468.910 -11.330 ;
        RECT 1469.330 -12.510 1470.510 -11.330 ;
        RECT 1467.730 -14.110 1468.910 -12.930 ;
        RECT 1469.330 -14.110 1470.510 -12.930 ;
        RECT 1647.730 3532.610 1648.910 3533.790 ;
        RECT 1649.330 3532.610 1650.510 3533.790 ;
        RECT 1647.730 3531.010 1648.910 3532.190 ;
        RECT 1649.330 3531.010 1650.510 3532.190 ;
        RECT 1647.730 3454.690 1648.910 3455.870 ;
        RECT 1649.330 3454.690 1650.510 3455.870 ;
        RECT 1647.730 3453.090 1648.910 3454.270 ;
        RECT 1649.330 3453.090 1650.510 3454.270 ;
        RECT 1647.730 3274.690 1648.910 3275.870 ;
        RECT 1649.330 3274.690 1650.510 3275.870 ;
        RECT 1647.730 3273.090 1648.910 3274.270 ;
        RECT 1649.330 3273.090 1650.510 3274.270 ;
        RECT 1647.730 3094.690 1648.910 3095.870 ;
        RECT 1649.330 3094.690 1650.510 3095.870 ;
        RECT 1647.730 3093.090 1648.910 3094.270 ;
        RECT 1649.330 3093.090 1650.510 3094.270 ;
        RECT 1647.730 2914.690 1648.910 2915.870 ;
        RECT 1649.330 2914.690 1650.510 2915.870 ;
        RECT 1647.730 2913.090 1648.910 2914.270 ;
        RECT 1649.330 2913.090 1650.510 2914.270 ;
        RECT 1647.730 2734.690 1648.910 2735.870 ;
        RECT 1649.330 2734.690 1650.510 2735.870 ;
        RECT 1647.730 2733.090 1648.910 2734.270 ;
        RECT 1649.330 2733.090 1650.510 2734.270 ;
        RECT 1647.730 2554.690 1648.910 2555.870 ;
        RECT 1649.330 2554.690 1650.510 2555.870 ;
        RECT 1647.730 2553.090 1648.910 2554.270 ;
        RECT 1649.330 2553.090 1650.510 2554.270 ;
        RECT 1647.730 2374.690 1648.910 2375.870 ;
        RECT 1649.330 2374.690 1650.510 2375.870 ;
        RECT 1647.730 2373.090 1648.910 2374.270 ;
        RECT 1649.330 2373.090 1650.510 2374.270 ;
        RECT 1647.730 2194.690 1648.910 2195.870 ;
        RECT 1649.330 2194.690 1650.510 2195.870 ;
        RECT 1647.730 2193.090 1648.910 2194.270 ;
        RECT 1649.330 2193.090 1650.510 2194.270 ;
        RECT 1647.730 2014.690 1648.910 2015.870 ;
        RECT 1649.330 2014.690 1650.510 2015.870 ;
        RECT 1647.730 2013.090 1648.910 2014.270 ;
        RECT 1649.330 2013.090 1650.510 2014.270 ;
        RECT 1647.730 1834.690 1648.910 1835.870 ;
        RECT 1649.330 1834.690 1650.510 1835.870 ;
        RECT 1647.730 1833.090 1648.910 1834.270 ;
        RECT 1649.330 1833.090 1650.510 1834.270 ;
        RECT 1647.730 1654.690 1648.910 1655.870 ;
        RECT 1649.330 1654.690 1650.510 1655.870 ;
        RECT 1647.730 1653.090 1648.910 1654.270 ;
        RECT 1649.330 1653.090 1650.510 1654.270 ;
        RECT 1647.730 1474.690 1648.910 1475.870 ;
        RECT 1649.330 1474.690 1650.510 1475.870 ;
        RECT 1647.730 1473.090 1648.910 1474.270 ;
        RECT 1649.330 1473.090 1650.510 1474.270 ;
        RECT 1647.730 1294.690 1648.910 1295.870 ;
        RECT 1649.330 1294.690 1650.510 1295.870 ;
        RECT 1647.730 1293.090 1648.910 1294.270 ;
        RECT 1649.330 1293.090 1650.510 1294.270 ;
        RECT 1647.730 1114.690 1648.910 1115.870 ;
        RECT 1649.330 1114.690 1650.510 1115.870 ;
        RECT 1647.730 1113.090 1648.910 1114.270 ;
        RECT 1649.330 1113.090 1650.510 1114.270 ;
        RECT 1647.730 934.690 1648.910 935.870 ;
        RECT 1649.330 934.690 1650.510 935.870 ;
        RECT 1647.730 933.090 1648.910 934.270 ;
        RECT 1649.330 933.090 1650.510 934.270 ;
        RECT 1647.730 754.690 1648.910 755.870 ;
        RECT 1649.330 754.690 1650.510 755.870 ;
        RECT 1647.730 753.090 1648.910 754.270 ;
        RECT 1649.330 753.090 1650.510 754.270 ;
        RECT 1647.730 574.690 1648.910 575.870 ;
        RECT 1649.330 574.690 1650.510 575.870 ;
        RECT 1647.730 573.090 1648.910 574.270 ;
        RECT 1649.330 573.090 1650.510 574.270 ;
        RECT 1647.730 394.690 1648.910 395.870 ;
        RECT 1649.330 394.690 1650.510 395.870 ;
        RECT 1647.730 393.090 1648.910 394.270 ;
        RECT 1649.330 393.090 1650.510 394.270 ;
        RECT 1647.730 214.690 1648.910 215.870 ;
        RECT 1649.330 214.690 1650.510 215.870 ;
        RECT 1647.730 213.090 1648.910 214.270 ;
        RECT 1649.330 213.090 1650.510 214.270 ;
        RECT 1647.730 34.690 1648.910 35.870 ;
        RECT 1649.330 34.690 1650.510 35.870 ;
        RECT 1647.730 33.090 1648.910 34.270 ;
        RECT 1649.330 33.090 1650.510 34.270 ;
        RECT 1647.730 -12.510 1648.910 -11.330 ;
        RECT 1649.330 -12.510 1650.510 -11.330 ;
        RECT 1647.730 -14.110 1648.910 -12.930 ;
        RECT 1649.330 -14.110 1650.510 -12.930 ;
        RECT 1827.730 3532.610 1828.910 3533.790 ;
        RECT 1829.330 3532.610 1830.510 3533.790 ;
        RECT 1827.730 3531.010 1828.910 3532.190 ;
        RECT 1829.330 3531.010 1830.510 3532.190 ;
        RECT 1827.730 3454.690 1828.910 3455.870 ;
        RECT 1829.330 3454.690 1830.510 3455.870 ;
        RECT 1827.730 3453.090 1828.910 3454.270 ;
        RECT 1829.330 3453.090 1830.510 3454.270 ;
        RECT 1827.730 3274.690 1828.910 3275.870 ;
        RECT 1829.330 3274.690 1830.510 3275.870 ;
        RECT 1827.730 3273.090 1828.910 3274.270 ;
        RECT 1829.330 3273.090 1830.510 3274.270 ;
        RECT 1827.730 3094.690 1828.910 3095.870 ;
        RECT 1829.330 3094.690 1830.510 3095.870 ;
        RECT 1827.730 3093.090 1828.910 3094.270 ;
        RECT 1829.330 3093.090 1830.510 3094.270 ;
        RECT 1827.730 2914.690 1828.910 2915.870 ;
        RECT 1829.330 2914.690 1830.510 2915.870 ;
        RECT 1827.730 2913.090 1828.910 2914.270 ;
        RECT 1829.330 2913.090 1830.510 2914.270 ;
        RECT 1827.730 2734.690 1828.910 2735.870 ;
        RECT 1829.330 2734.690 1830.510 2735.870 ;
        RECT 1827.730 2733.090 1828.910 2734.270 ;
        RECT 1829.330 2733.090 1830.510 2734.270 ;
        RECT 1827.730 2554.690 1828.910 2555.870 ;
        RECT 1829.330 2554.690 1830.510 2555.870 ;
        RECT 1827.730 2553.090 1828.910 2554.270 ;
        RECT 1829.330 2553.090 1830.510 2554.270 ;
        RECT 1827.730 2374.690 1828.910 2375.870 ;
        RECT 1829.330 2374.690 1830.510 2375.870 ;
        RECT 1827.730 2373.090 1828.910 2374.270 ;
        RECT 1829.330 2373.090 1830.510 2374.270 ;
        RECT 1827.730 2194.690 1828.910 2195.870 ;
        RECT 1829.330 2194.690 1830.510 2195.870 ;
        RECT 1827.730 2193.090 1828.910 2194.270 ;
        RECT 1829.330 2193.090 1830.510 2194.270 ;
        RECT 1827.730 2014.690 1828.910 2015.870 ;
        RECT 1829.330 2014.690 1830.510 2015.870 ;
        RECT 1827.730 2013.090 1828.910 2014.270 ;
        RECT 1829.330 2013.090 1830.510 2014.270 ;
        RECT 1827.730 1834.690 1828.910 1835.870 ;
        RECT 1829.330 1834.690 1830.510 1835.870 ;
        RECT 1827.730 1833.090 1828.910 1834.270 ;
        RECT 1829.330 1833.090 1830.510 1834.270 ;
        RECT 1827.730 1654.690 1828.910 1655.870 ;
        RECT 1829.330 1654.690 1830.510 1655.870 ;
        RECT 1827.730 1653.090 1828.910 1654.270 ;
        RECT 1829.330 1653.090 1830.510 1654.270 ;
        RECT 1827.730 1474.690 1828.910 1475.870 ;
        RECT 1829.330 1474.690 1830.510 1475.870 ;
        RECT 1827.730 1473.090 1828.910 1474.270 ;
        RECT 1829.330 1473.090 1830.510 1474.270 ;
        RECT 1827.730 1294.690 1828.910 1295.870 ;
        RECT 1829.330 1294.690 1830.510 1295.870 ;
        RECT 1827.730 1293.090 1828.910 1294.270 ;
        RECT 1829.330 1293.090 1830.510 1294.270 ;
        RECT 1827.730 1114.690 1828.910 1115.870 ;
        RECT 1829.330 1114.690 1830.510 1115.870 ;
        RECT 1827.730 1113.090 1828.910 1114.270 ;
        RECT 1829.330 1113.090 1830.510 1114.270 ;
        RECT 1827.730 934.690 1828.910 935.870 ;
        RECT 1829.330 934.690 1830.510 935.870 ;
        RECT 1827.730 933.090 1828.910 934.270 ;
        RECT 1829.330 933.090 1830.510 934.270 ;
        RECT 1827.730 754.690 1828.910 755.870 ;
        RECT 1829.330 754.690 1830.510 755.870 ;
        RECT 1827.730 753.090 1828.910 754.270 ;
        RECT 1829.330 753.090 1830.510 754.270 ;
        RECT 1827.730 574.690 1828.910 575.870 ;
        RECT 1829.330 574.690 1830.510 575.870 ;
        RECT 1827.730 573.090 1828.910 574.270 ;
        RECT 1829.330 573.090 1830.510 574.270 ;
        RECT 1827.730 394.690 1828.910 395.870 ;
        RECT 1829.330 394.690 1830.510 395.870 ;
        RECT 1827.730 393.090 1828.910 394.270 ;
        RECT 1829.330 393.090 1830.510 394.270 ;
        RECT 1827.730 214.690 1828.910 215.870 ;
        RECT 1829.330 214.690 1830.510 215.870 ;
        RECT 1827.730 213.090 1828.910 214.270 ;
        RECT 1829.330 213.090 1830.510 214.270 ;
        RECT 1827.730 34.690 1828.910 35.870 ;
        RECT 1829.330 34.690 1830.510 35.870 ;
        RECT 1827.730 33.090 1828.910 34.270 ;
        RECT 1829.330 33.090 1830.510 34.270 ;
        RECT 1827.730 -12.510 1828.910 -11.330 ;
        RECT 1829.330 -12.510 1830.510 -11.330 ;
        RECT 1827.730 -14.110 1828.910 -12.930 ;
        RECT 1829.330 -14.110 1830.510 -12.930 ;
        RECT 2007.730 3532.610 2008.910 3533.790 ;
        RECT 2009.330 3532.610 2010.510 3533.790 ;
        RECT 2007.730 3531.010 2008.910 3532.190 ;
        RECT 2009.330 3531.010 2010.510 3532.190 ;
        RECT 2007.730 3454.690 2008.910 3455.870 ;
        RECT 2009.330 3454.690 2010.510 3455.870 ;
        RECT 2007.730 3453.090 2008.910 3454.270 ;
        RECT 2009.330 3453.090 2010.510 3454.270 ;
        RECT 2007.730 3274.690 2008.910 3275.870 ;
        RECT 2009.330 3274.690 2010.510 3275.870 ;
        RECT 2007.730 3273.090 2008.910 3274.270 ;
        RECT 2009.330 3273.090 2010.510 3274.270 ;
        RECT 2007.730 3094.690 2008.910 3095.870 ;
        RECT 2009.330 3094.690 2010.510 3095.870 ;
        RECT 2007.730 3093.090 2008.910 3094.270 ;
        RECT 2009.330 3093.090 2010.510 3094.270 ;
        RECT 2007.730 2914.690 2008.910 2915.870 ;
        RECT 2009.330 2914.690 2010.510 2915.870 ;
        RECT 2007.730 2913.090 2008.910 2914.270 ;
        RECT 2009.330 2913.090 2010.510 2914.270 ;
        RECT 2007.730 2734.690 2008.910 2735.870 ;
        RECT 2009.330 2734.690 2010.510 2735.870 ;
        RECT 2007.730 2733.090 2008.910 2734.270 ;
        RECT 2009.330 2733.090 2010.510 2734.270 ;
        RECT 2007.730 2554.690 2008.910 2555.870 ;
        RECT 2009.330 2554.690 2010.510 2555.870 ;
        RECT 2007.730 2553.090 2008.910 2554.270 ;
        RECT 2009.330 2553.090 2010.510 2554.270 ;
        RECT 2007.730 2374.690 2008.910 2375.870 ;
        RECT 2009.330 2374.690 2010.510 2375.870 ;
        RECT 2007.730 2373.090 2008.910 2374.270 ;
        RECT 2009.330 2373.090 2010.510 2374.270 ;
        RECT 2007.730 2194.690 2008.910 2195.870 ;
        RECT 2009.330 2194.690 2010.510 2195.870 ;
        RECT 2007.730 2193.090 2008.910 2194.270 ;
        RECT 2009.330 2193.090 2010.510 2194.270 ;
        RECT 2007.730 2014.690 2008.910 2015.870 ;
        RECT 2009.330 2014.690 2010.510 2015.870 ;
        RECT 2007.730 2013.090 2008.910 2014.270 ;
        RECT 2009.330 2013.090 2010.510 2014.270 ;
        RECT 2007.730 1834.690 2008.910 1835.870 ;
        RECT 2009.330 1834.690 2010.510 1835.870 ;
        RECT 2007.730 1833.090 2008.910 1834.270 ;
        RECT 2009.330 1833.090 2010.510 1834.270 ;
        RECT 2007.730 1654.690 2008.910 1655.870 ;
        RECT 2009.330 1654.690 2010.510 1655.870 ;
        RECT 2007.730 1653.090 2008.910 1654.270 ;
        RECT 2009.330 1653.090 2010.510 1654.270 ;
        RECT 2007.730 1474.690 2008.910 1475.870 ;
        RECT 2009.330 1474.690 2010.510 1475.870 ;
        RECT 2007.730 1473.090 2008.910 1474.270 ;
        RECT 2009.330 1473.090 2010.510 1474.270 ;
        RECT 2007.730 1294.690 2008.910 1295.870 ;
        RECT 2009.330 1294.690 2010.510 1295.870 ;
        RECT 2007.730 1293.090 2008.910 1294.270 ;
        RECT 2009.330 1293.090 2010.510 1294.270 ;
        RECT 2007.730 1114.690 2008.910 1115.870 ;
        RECT 2009.330 1114.690 2010.510 1115.870 ;
        RECT 2007.730 1113.090 2008.910 1114.270 ;
        RECT 2009.330 1113.090 2010.510 1114.270 ;
        RECT 2007.730 934.690 2008.910 935.870 ;
        RECT 2009.330 934.690 2010.510 935.870 ;
        RECT 2007.730 933.090 2008.910 934.270 ;
        RECT 2009.330 933.090 2010.510 934.270 ;
        RECT 2007.730 754.690 2008.910 755.870 ;
        RECT 2009.330 754.690 2010.510 755.870 ;
        RECT 2007.730 753.090 2008.910 754.270 ;
        RECT 2009.330 753.090 2010.510 754.270 ;
        RECT 2007.730 574.690 2008.910 575.870 ;
        RECT 2009.330 574.690 2010.510 575.870 ;
        RECT 2007.730 573.090 2008.910 574.270 ;
        RECT 2009.330 573.090 2010.510 574.270 ;
        RECT 2007.730 394.690 2008.910 395.870 ;
        RECT 2009.330 394.690 2010.510 395.870 ;
        RECT 2007.730 393.090 2008.910 394.270 ;
        RECT 2009.330 393.090 2010.510 394.270 ;
        RECT 2007.730 214.690 2008.910 215.870 ;
        RECT 2009.330 214.690 2010.510 215.870 ;
        RECT 2007.730 213.090 2008.910 214.270 ;
        RECT 2009.330 213.090 2010.510 214.270 ;
        RECT 2007.730 34.690 2008.910 35.870 ;
        RECT 2009.330 34.690 2010.510 35.870 ;
        RECT 2007.730 33.090 2008.910 34.270 ;
        RECT 2009.330 33.090 2010.510 34.270 ;
        RECT 2007.730 -12.510 2008.910 -11.330 ;
        RECT 2009.330 -12.510 2010.510 -11.330 ;
        RECT 2007.730 -14.110 2008.910 -12.930 ;
        RECT 2009.330 -14.110 2010.510 -12.930 ;
        RECT 2187.730 3532.610 2188.910 3533.790 ;
        RECT 2189.330 3532.610 2190.510 3533.790 ;
        RECT 2187.730 3531.010 2188.910 3532.190 ;
        RECT 2189.330 3531.010 2190.510 3532.190 ;
        RECT 2187.730 3454.690 2188.910 3455.870 ;
        RECT 2189.330 3454.690 2190.510 3455.870 ;
        RECT 2187.730 3453.090 2188.910 3454.270 ;
        RECT 2189.330 3453.090 2190.510 3454.270 ;
        RECT 2187.730 3274.690 2188.910 3275.870 ;
        RECT 2189.330 3274.690 2190.510 3275.870 ;
        RECT 2187.730 3273.090 2188.910 3274.270 ;
        RECT 2189.330 3273.090 2190.510 3274.270 ;
        RECT 2187.730 3094.690 2188.910 3095.870 ;
        RECT 2189.330 3094.690 2190.510 3095.870 ;
        RECT 2187.730 3093.090 2188.910 3094.270 ;
        RECT 2189.330 3093.090 2190.510 3094.270 ;
        RECT 2187.730 2914.690 2188.910 2915.870 ;
        RECT 2189.330 2914.690 2190.510 2915.870 ;
        RECT 2187.730 2913.090 2188.910 2914.270 ;
        RECT 2189.330 2913.090 2190.510 2914.270 ;
        RECT 2187.730 2734.690 2188.910 2735.870 ;
        RECT 2189.330 2734.690 2190.510 2735.870 ;
        RECT 2187.730 2733.090 2188.910 2734.270 ;
        RECT 2189.330 2733.090 2190.510 2734.270 ;
        RECT 2187.730 2554.690 2188.910 2555.870 ;
        RECT 2189.330 2554.690 2190.510 2555.870 ;
        RECT 2187.730 2553.090 2188.910 2554.270 ;
        RECT 2189.330 2553.090 2190.510 2554.270 ;
        RECT 2187.730 2374.690 2188.910 2375.870 ;
        RECT 2189.330 2374.690 2190.510 2375.870 ;
        RECT 2187.730 2373.090 2188.910 2374.270 ;
        RECT 2189.330 2373.090 2190.510 2374.270 ;
        RECT 2187.730 2194.690 2188.910 2195.870 ;
        RECT 2189.330 2194.690 2190.510 2195.870 ;
        RECT 2187.730 2193.090 2188.910 2194.270 ;
        RECT 2189.330 2193.090 2190.510 2194.270 ;
        RECT 2187.730 2014.690 2188.910 2015.870 ;
        RECT 2189.330 2014.690 2190.510 2015.870 ;
        RECT 2187.730 2013.090 2188.910 2014.270 ;
        RECT 2189.330 2013.090 2190.510 2014.270 ;
        RECT 2187.730 1834.690 2188.910 1835.870 ;
        RECT 2189.330 1834.690 2190.510 1835.870 ;
        RECT 2187.730 1833.090 2188.910 1834.270 ;
        RECT 2189.330 1833.090 2190.510 1834.270 ;
        RECT 2187.730 1654.690 2188.910 1655.870 ;
        RECT 2189.330 1654.690 2190.510 1655.870 ;
        RECT 2187.730 1653.090 2188.910 1654.270 ;
        RECT 2189.330 1653.090 2190.510 1654.270 ;
        RECT 2187.730 1474.690 2188.910 1475.870 ;
        RECT 2189.330 1474.690 2190.510 1475.870 ;
        RECT 2187.730 1473.090 2188.910 1474.270 ;
        RECT 2189.330 1473.090 2190.510 1474.270 ;
        RECT 2187.730 1294.690 2188.910 1295.870 ;
        RECT 2189.330 1294.690 2190.510 1295.870 ;
        RECT 2187.730 1293.090 2188.910 1294.270 ;
        RECT 2189.330 1293.090 2190.510 1294.270 ;
        RECT 2187.730 1114.690 2188.910 1115.870 ;
        RECT 2189.330 1114.690 2190.510 1115.870 ;
        RECT 2187.730 1113.090 2188.910 1114.270 ;
        RECT 2189.330 1113.090 2190.510 1114.270 ;
        RECT 2187.730 934.690 2188.910 935.870 ;
        RECT 2189.330 934.690 2190.510 935.870 ;
        RECT 2187.730 933.090 2188.910 934.270 ;
        RECT 2189.330 933.090 2190.510 934.270 ;
        RECT 2187.730 754.690 2188.910 755.870 ;
        RECT 2189.330 754.690 2190.510 755.870 ;
        RECT 2187.730 753.090 2188.910 754.270 ;
        RECT 2189.330 753.090 2190.510 754.270 ;
        RECT 2187.730 574.690 2188.910 575.870 ;
        RECT 2189.330 574.690 2190.510 575.870 ;
        RECT 2187.730 573.090 2188.910 574.270 ;
        RECT 2189.330 573.090 2190.510 574.270 ;
        RECT 2187.730 394.690 2188.910 395.870 ;
        RECT 2189.330 394.690 2190.510 395.870 ;
        RECT 2187.730 393.090 2188.910 394.270 ;
        RECT 2189.330 393.090 2190.510 394.270 ;
        RECT 2187.730 214.690 2188.910 215.870 ;
        RECT 2189.330 214.690 2190.510 215.870 ;
        RECT 2187.730 213.090 2188.910 214.270 ;
        RECT 2189.330 213.090 2190.510 214.270 ;
        RECT 2187.730 34.690 2188.910 35.870 ;
        RECT 2189.330 34.690 2190.510 35.870 ;
        RECT 2187.730 33.090 2188.910 34.270 ;
        RECT 2189.330 33.090 2190.510 34.270 ;
        RECT 2187.730 -12.510 2188.910 -11.330 ;
        RECT 2189.330 -12.510 2190.510 -11.330 ;
        RECT 2187.730 -14.110 2188.910 -12.930 ;
        RECT 2189.330 -14.110 2190.510 -12.930 ;
        RECT 2367.730 3532.610 2368.910 3533.790 ;
        RECT 2369.330 3532.610 2370.510 3533.790 ;
        RECT 2367.730 3531.010 2368.910 3532.190 ;
        RECT 2369.330 3531.010 2370.510 3532.190 ;
        RECT 2367.730 3454.690 2368.910 3455.870 ;
        RECT 2369.330 3454.690 2370.510 3455.870 ;
        RECT 2367.730 3453.090 2368.910 3454.270 ;
        RECT 2369.330 3453.090 2370.510 3454.270 ;
        RECT 2367.730 3274.690 2368.910 3275.870 ;
        RECT 2369.330 3274.690 2370.510 3275.870 ;
        RECT 2367.730 3273.090 2368.910 3274.270 ;
        RECT 2369.330 3273.090 2370.510 3274.270 ;
        RECT 2367.730 3094.690 2368.910 3095.870 ;
        RECT 2369.330 3094.690 2370.510 3095.870 ;
        RECT 2367.730 3093.090 2368.910 3094.270 ;
        RECT 2369.330 3093.090 2370.510 3094.270 ;
        RECT 2367.730 2914.690 2368.910 2915.870 ;
        RECT 2369.330 2914.690 2370.510 2915.870 ;
        RECT 2367.730 2913.090 2368.910 2914.270 ;
        RECT 2369.330 2913.090 2370.510 2914.270 ;
        RECT 2367.730 2734.690 2368.910 2735.870 ;
        RECT 2369.330 2734.690 2370.510 2735.870 ;
        RECT 2367.730 2733.090 2368.910 2734.270 ;
        RECT 2369.330 2733.090 2370.510 2734.270 ;
        RECT 2367.730 2554.690 2368.910 2555.870 ;
        RECT 2369.330 2554.690 2370.510 2555.870 ;
        RECT 2367.730 2553.090 2368.910 2554.270 ;
        RECT 2369.330 2553.090 2370.510 2554.270 ;
        RECT 2367.730 2374.690 2368.910 2375.870 ;
        RECT 2369.330 2374.690 2370.510 2375.870 ;
        RECT 2367.730 2373.090 2368.910 2374.270 ;
        RECT 2369.330 2373.090 2370.510 2374.270 ;
        RECT 2367.730 2194.690 2368.910 2195.870 ;
        RECT 2369.330 2194.690 2370.510 2195.870 ;
        RECT 2367.730 2193.090 2368.910 2194.270 ;
        RECT 2369.330 2193.090 2370.510 2194.270 ;
        RECT 2367.730 2014.690 2368.910 2015.870 ;
        RECT 2369.330 2014.690 2370.510 2015.870 ;
        RECT 2367.730 2013.090 2368.910 2014.270 ;
        RECT 2369.330 2013.090 2370.510 2014.270 ;
        RECT 2367.730 1834.690 2368.910 1835.870 ;
        RECT 2369.330 1834.690 2370.510 1835.870 ;
        RECT 2367.730 1833.090 2368.910 1834.270 ;
        RECT 2369.330 1833.090 2370.510 1834.270 ;
        RECT 2367.730 1654.690 2368.910 1655.870 ;
        RECT 2369.330 1654.690 2370.510 1655.870 ;
        RECT 2367.730 1653.090 2368.910 1654.270 ;
        RECT 2369.330 1653.090 2370.510 1654.270 ;
        RECT 2367.730 1474.690 2368.910 1475.870 ;
        RECT 2369.330 1474.690 2370.510 1475.870 ;
        RECT 2367.730 1473.090 2368.910 1474.270 ;
        RECT 2369.330 1473.090 2370.510 1474.270 ;
        RECT 2367.730 1294.690 2368.910 1295.870 ;
        RECT 2369.330 1294.690 2370.510 1295.870 ;
        RECT 2367.730 1293.090 2368.910 1294.270 ;
        RECT 2369.330 1293.090 2370.510 1294.270 ;
        RECT 2367.730 1114.690 2368.910 1115.870 ;
        RECT 2369.330 1114.690 2370.510 1115.870 ;
        RECT 2367.730 1113.090 2368.910 1114.270 ;
        RECT 2369.330 1113.090 2370.510 1114.270 ;
        RECT 2367.730 934.690 2368.910 935.870 ;
        RECT 2369.330 934.690 2370.510 935.870 ;
        RECT 2367.730 933.090 2368.910 934.270 ;
        RECT 2369.330 933.090 2370.510 934.270 ;
        RECT 2367.730 754.690 2368.910 755.870 ;
        RECT 2369.330 754.690 2370.510 755.870 ;
        RECT 2367.730 753.090 2368.910 754.270 ;
        RECT 2369.330 753.090 2370.510 754.270 ;
        RECT 2367.730 574.690 2368.910 575.870 ;
        RECT 2369.330 574.690 2370.510 575.870 ;
        RECT 2367.730 573.090 2368.910 574.270 ;
        RECT 2369.330 573.090 2370.510 574.270 ;
        RECT 2367.730 394.690 2368.910 395.870 ;
        RECT 2369.330 394.690 2370.510 395.870 ;
        RECT 2367.730 393.090 2368.910 394.270 ;
        RECT 2369.330 393.090 2370.510 394.270 ;
        RECT 2367.730 214.690 2368.910 215.870 ;
        RECT 2369.330 214.690 2370.510 215.870 ;
        RECT 2367.730 213.090 2368.910 214.270 ;
        RECT 2369.330 213.090 2370.510 214.270 ;
        RECT 2367.730 34.690 2368.910 35.870 ;
        RECT 2369.330 34.690 2370.510 35.870 ;
        RECT 2367.730 33.090 2368.910 34.270 ;
        RECT 2369.330 33.090 2370.510 34.270 ;
        RECT 2367.730 -12.510 2368.910 -11.330 ;
        RECT 2369.330 -12.510 2370.510 -11.330 ;
        RECT 2367.730 -14.110 2368.910 -12.930 ;
        RECT 2369.330 -14.110 2370.510 -12.930 ;
        RECT 2547.730 3532.610 2548.910 3533.790 ;
        RECT 2549.330 3532.610 2550.510 3533.790 ;
        RECT 2547.730 3531.010 2548.910 3532.190 ;
        RECT 2549.330 3531.010 2550.510 3532.190 ;
        RECT 2547.730 3454.690 2548.910 3455.870 ;
        RECT 2549.330 3454.690 2550.510 3455.870 ;
        RECT 2547.730 3453.090 2548.910 3454.270 ;
        RECT 2549.330 3453.090 2550.510 3454.270 ;
        RECT 2547.730 3274.690 2548.910 3275.870 ;
        RECT 2549.330 3274.690 2550.510 3275.870 ;
        RECT 2547.730 3273.090 2548.910 3274.270 ;
        RECT 2549.330 3273.090 2550.510 3274.270 ;
        RECT 2547.730 3094.690 2548.910 3095.870 ;
        RECT 2549.330 3094.690 2550.510 3095.870 ;
        RECT 2547.730 3093.090 2548.910 3094.270 ;
        RECT 2549.330 3093.090 2550.510 3094.270 ;
        RECT 2547.730 2914.690 2548.910 2915.870 ;
        RECT 2549.330 2914.690 2550.510 2915.870 ;
        RECT 2547.730 2913.090 2548.910 2914.270 ;
        RECT 2549.330 2913.090 2550.510 2914.270 ;
        RECT 2547.730 2734.690 2548.910 2735.870 ;
        RECT 2549.330 2734.690 2550.510 2735.870 ;
        RECT 2547.730 2733.090 2548.910 2734.270 ;
        RECT 2549.330 2733.090 2550.510 2734.270 ;
        RECT 2547.730 2554.690 2548.910 2555.870 ;
        RECT 2549.330 2554.690 2550.510 2555.870 ;
        RECT 2547.730 2553.090 2548.910 2554.270 ;
        RECT 2549.330 2553.090 2550.510 2554.270 ;
        RECT 2547.730 2374.690 2548.910 2375.870 ;
        RECT 2549.330 2374.690 2550.510 2375.870 ;
        RECT 2547.730 2373.090 2548.910 2374.270 ;
        RECT 2549.330 2373.090 2550.510 2374.270 ;
        RECT 2547.730 2194.690 2548.910 2195.870 ;
        RECT 2549.330 2194.690 2550.510 2195.870 ;
        RECT 2547.730 2193.090 2548.910 2194.270 ;
        RECT 2549.330 2193.090 2550.510 2194.270 ;
        RECT 2547.730 2014.690 2548.910 2015.870 ;
        RECT 2549.330 2014.690 2550.510 2015.870 ;
        RECT 2547.730 2013.090 2548.910 2014.270 ;
        RECT 2549.330 2013.090 2550.510 2014.270 ;
        RECT 2547.730 1834.690 2548.910 1835.870 ;
        RECT 2549.330 1834.690 2550.510 1835.870 ;
        RECT 2547.730 1833.090 2548.910 1834.270 ;
        RECT 2549.330 1833.090 2550.510 1834.270 ;
        RECT 2547.730 1654.690 2548.910 1655.870 ;
        RECT 2549.330 1654.690 2550.510 1655.870 ;
        RECT 2547.730 1653.090 2548.910 1654.270 ;
        RECT 2549.330 1653.090 2550.510 1654.270 ;
        RECT 2547.730 1474.690 2548.910 1475.870 ;
        RECT 2549.330 1474.690 2550.510 1475.870 ;
        RECT 2547.730 1473.090 2548.910 1474.270 ;
        RECT 2549.330 1473.090 2550.510 1474.270 ;
        RECT 2547.730 1294.690 2548.910 1295.870 ;
        RECT 2549.330 1294.690 2550.510 1295.870 ;
        RECT 2547.730 1293.090 2548.910 1294.270 ;
        RECT 2549.330 1293.090 2550.510 1294.270 ;
        RECT 2547.730 1114.690 2548.910 1115.870 ;
        RECT 2549.330 1114.690 2550.510 1115.870 ;
        RECT 2547.730 1113.090 2548.910 1114.270 ;
        RECT 2549.330 1113.090 2550.510 1114.270 ;
        RECT 2547.730 934.690 2548.910 935.870 ;
        RECT 2549.330 934.690 2550.510 935.870 ;
        RECT 2547.730 933.090 2548.910 934.270 ;
        RECT 2549.330 933.090 2550.510 934.270 ;
        RECT 2547.730 754.690 2548.910 755.870 ;
        RECT 2549.330 754.690 2550.510 755.870 ;
        RECT 2547.730 753.090 2548.910 754.270 ;
        RECT 2549.330 753.090 2550.510 754.270 ;
        RECT 2547.730 574.690 2548.910 575.870 ;
        RECT 2549.330 574.690 2550.510 575.870 ;
        RECT 2547.730 573.090 2548.910 574.270 ;
        RECT 2549.330 573.090 2550.510 574.270 ;
        RECT 2547.730 394.690 2548.910 395.870 ;
        RECT 2549.330 394.690 2550.510 395.870 ;
        RECT 2547.730 393.090 2548.910 394.270 ;
        RECT 2549.330 393.090 2550.510 394.270 ;
        RECT 2547.730 214.690 2548.910 215.870 ;
        RECT 2549.330 214.690 2550.510 215.870 ;
        RECT 2547.730 213.090 2548.910 214.270 ;
        RECT 2549.330 213.090 2550.510 214.270 ;
        RECT 2547.730 34.690 2548.910 35.870 ;
        RECT 2549.330 34.690 2550.510 35.870 ;
        RECT 2547.730 33.090 2548.910 34.270 ;
        RECT 2549.330 33.090 2550.510 34.270 ;
        RECT 2547.730 -12.510 2548.910 -11.330 ;
        RECT 2549.330 -12.510 2550.510 -11.330 ;
        RECT 2547.730 -14.110 2548.910 -12.930 ;
        RECT 2549.330 -14.110 2550.510 -12.930 ;
        RECT 2727.730 3532.610 2728.910 3533.790 ;
        RECT 2729.330 3532.610 2730.510 3533.790 ;
        RECT 2727.730 3531.010 2728.910 3532.190 ;
        RECT 2729.330 3531.010 2730.510 3532.190 ;
        RECT 2727.730 3454.690 2728.910 3455.870 ;
        RECT 2729.330 3454.690 2730.510 3455.870 ;
        RECT 2727.730 3453.090 2728.910 3454.270 ;
        RECT 2729.330 3453.090 2730.510 3454.270 ;
        RECT 2727.730 3274.690 2728.910 3275.870 ;
        RECT 2729.330 3274.690 2730.510 3275.870 ;
        RECT 2727.730 3273.090 2728.910 3274.270 ;
        RECT 2729.330 3273.090 2730.510 3274.270 ;
        RECT 2727.730 3094.690 2728.910 3095.870 ;
        RECT 2729.330 3094.690 2730.510 3095.870 ;
        RECT 2727.730 3093.090 2728.910 3094.270 ;
        RECT 2729.330 3093.090 2730.510 3094.270 ;
        RECT 2727.730 2914.690 2728.910 2915.870 ;
        RECT 2729.330 2914.690 2730.510 2915.870 ;
        RECT 2727.730 2913.090 2728.910 2914.270 ;
        RECT 2729.330 2913.090 2730.510 2914.270 ;
        RECT 2727.730 2734.690 2728.910 2735.870 ;
        RECT 2729.330 2734.690 2730.510 2735.870 ;
        RECT 2727.730 2733.090 2728.910 2734.270 ;
        RECT 2729.330 2733.090 2730.510 2734.270 ;
        RECT 2727.730 2554.690 2728.910 2555.870 ;
        RECT 2729.330 2554.690 2730.510 2555.870 ;
        RECT 2727.730 2553.090 2728.910 2554.270 ;
        RECT 2729.330 2553.090 2730.510 2554.270 ;
        RECT 2727.730 2374.690 2728.910 2375.870 ;
        RECT 2729.330 2374.690 2730.510 2375.870 ;
        RECT 2727.730 2373.090 2728.910 2374.270 ;
        RECT 2729.330 2373.090 2730.510 2374.270 ;
        RECT 2727.730 2194.690 2728.910 2195.870 ;
        RECT 2729.330 2194.690 2730.510 2195.870 ;
        RECT 2727.730 2193.090 2728.910 2194.270 ;
        RECT 2729.330 2193.090 2730.510 2194.270 ;
        RECT 2727.730 2014.690 2728.910 2015.870 ;
        RECT 2729.330 2014.690 2730.510 2015.870 ;
        RECT 2727.730 2013.090 2728.910 2014.270 ;
        RECT 2729.330 2013.090 2730.510 2014.270 ;
        RECT 2727.730 1834.690 2728.910 1835.870 ;
        RECT 2729.330 1834.690 2730.510 1835.870 ;
        RECT 2727.730 1833.090 2728.910 1834.270 ;
        RECT 2729.330 1833.090 2730.510 1834.270 ;
        RECT 2727.730 1654.690 2728.910 1655.870 ;
        RECT 2729.330 1654.690 2730.510 1655.870 ;
        RECT 2727.730 1653.090 2728.910 1654.270 ;
        RECT 2729.330 1653.090 2730.510 1654.270 ;
        RECT 2727.730 1474.690 2728.910 1475.870 ;
        RECT 2729.330 1474.690 2730.510 1475.870 ;
        RECT 2727.730 1473.090 2728.910 1474.270 ;
        RECT 2729.330 1473.090 2730.510 1474.270 ;
        RECT 2727.730 1294.690 2728.910 1295.870 ;
        RECT 2729.330 1294.690 2730.510 1295.870 ;
        RECT 2727.730 1293.090 2728.910 1294.270 ;
        RECT 2729.330 1293.090 2730.510 1294.270 ;
        RECT 2727.730 1114.690 2728.910 1115.870 ;
        RECT 2729.330 1114.690 2730.510 1115.870 ;
        RECT 2727.730 1113.090 2728.910 1114.270 ;
        RECT 2729.330 1113.090 2730.510 1114.270 ;
        RECT 2727.730 934.690 2728.910 935.870 ;
        RECT 2729.330 934.690 2730.510 935.870 ;
        RECT 2727.730 933.090 2728.910 934.270 ;
        RECT 2729.330 933.090 2730.510 934.270 ;
        RECT 2727.730 754.690 2728.910 755.870 ;
        RECT 2729.330 754.690 2730.510 755.870 ;
        RECT 2727.730 753.090 2728.910 754.270 ;
        RECT 2729.330 753.090 2730.510 754.270 ;
        RECT 2727.730 574.690 2728.910 575.870 ;
        RECT 2729.330 574.690 2730.510 575.870 ;
        RECT 2727.730 573.090 2728.910 574.270 ;
        RECT 2729.330 573.090 2730.510 574.270 ;
        RECT 2727.730 394.690 2728.910 395.870 ;
        RECT 2729.330 394.690 2730.510 395.870 ;
        RECT 2727.730 393.090 2728.910 394.270 ;
        RECT 2729.330 393.090 2730.510 394.270 ;
        RECT 2727.730 214.690 2728.910 215.870 ;
        RECT 2729.330 214.690 2730.510 215.870 ;
        RECT 2727.730 213.090 2728.910 214.270 ;
        RECT 2729.330 213.090 2730.510 214.270 ;
        RECT 2727.730 34.690 2728.910 35.870 ;
        RECT 2729.330 34.690 2730.510 35.870 ;
        RECT 2727.730 33.090 2728.910 34.270 ;
        RECT 2729.330 33.090 2730.510 34.270 ;
        RECT 2727.730 -12.510 2728.910 -11.330 ;
        RECT 2729.330 -12.510 2730.510 -11.330 ;
        RECT 2727.730 -14.110 2728.910 -12.930 ;
        RECT 2729.330 -14.110 2730.510 -12.930 ;
        RECT 2907.730 3532.610 2908.910 3533.790 ;
        RECT 2909.330 3532.610 2910.510 3533.790 ;
        RECT 2907.730 3531.010 2908.910 3532.190 ;
        RECT 2909.330 3531.010 2910.510 3532.190 ;
        RECT 2907.730 3454.690 2908.910 3455.870 ;
        RECT 2909.330 3454.690 2910.510 3455.870 ;
        RECT 2907.730 3453.090 2908.910 3454.270 ;
        RECT 2909.330 3453.090 2910.510 3454.270 ;
        RECT 2907.730 3274.690 2908.910 3275.870 ;
        RECT 2909.330 3274.690 2910.510 3275.870 ;
        RECT 2907.730 3273.090 2908.910 3274.270 ;
        RECT 2909.330 3273.090 2910.510 3274.270 ;
        RECT 2907.730 3094.690 2908.910 3095.870 ;
        RECT 2909.330 3094.690 2910.510 3095.870 ;
        RECT 2907.730 3093.090 2908.910 3094.270 ;
        RECT 2909.330 3093.090 2910.510 3094.270 ;
        RECT 2907.730 2914.690 2908.910 2915.870 ;
        RECT 2909.330 2914.690 2910.510 2915.870 ;
        RECT 2907.730 2913.090 2908.910 2914.270 ;
        RECT 2909.330 2913.090 2910.510 2914.270 ;
        RECT 2907.730 2734.690 2908.910 2735.870 ;
        RECT 2909.330 2734.690 2910.510 2735.870 ;
        RECT 2907.730 2733.090 2908.910 2734.270 ;
        RECT 2909.330 2733.090 2910.510 2734.270 ;
        RECT 2907.730 2554.690 2908.910 2555.870 ;
        RECT 2909.330 2554.690 2910.510 2555.870 ;
        RECT 2907.730 2553.090 2908.910 2554.270 ;
        RECT 2909.330 2553.090 2910.510 2554.270 ;
        RECT 2907.730 2374.690 2908.910 2375.870 ;
        RECT 2909.330 2374.690 2910.510 2375.870 ;
        RECT 2907.730 2373.090 2908.910 2374.270 ;
        RECT 2909.330 2373.090 2910.510 2374.270 ;
        RECT 2907.730 2194.690 2908.910 2195.870 ;
        RECT 2909.330 2194.690 2910.510 2195.870 ;
        RECT 2907.730 2193.090 2908.910 2194.270 ;
        RECT 2909.330 2193.090 2910.510 2194.270 ;
        RECT 2907.730 2014.690 2908.910 2015.870 ;
        RECT 2909.330 2014.690 2910.510 2015.870 ;
        RECT 2907.730 2013.090 2908.910 2014.270 ;
        RECT 2909.330 2013.090 2910.510 2014.270 ;
        RECT 2907.730 1834.690 2908.910 1835.870 ;
        RECT 2909.330 1834.690 2910.510 1835.870 ;
        RECT 2907.730 1833.090 2908.910 1834.270 ;
        RECT 2909.330 1833.090 2910.510 1834.270 ;
        RECT 2907.730 1654.690 2908.910 1655.870 ;
        RECT 2909.330 1654.690 2910.510 1655.870 ;
        RECT 2907.730 1653.090 2908.910 1654.270 ;
        RECT 2909.330 1653.090 2910.510 1654.270 ;
        RECT 2907.730 1474.690 2908.910 1475.870 ;
        RECT 2909.330 1474.690 2910.510 1475.870 ;
        RECT 2907.730 1473.090 2908.910 1474.270 ;
        RECT 2909.330 1473.090 2910.510 1474.270 ;
        RECT 2907.730 1294.690 2908.910 1295.870 ;
        RECT 2909.330 1294.690 2910.510 1295.870 ;
        RECT 2907.730 1293.090 2908.910 1294.270 ;
        RECT 2909.330 1293.090 2910.510 1294.270 ;
        RECT 2907.730 1114.690 2908.910 1115.870 ;
        RECT 2909.330 1114.690 2910.510 1115.870 ;
        RECT 2907.730 1113.090 2908.910 1114.270 ;
        RECT 2909.330 1113.090 2910.510 1114.270 ;
        RECT 2907.730 934.690 2908.910 935.870 ;
        RECT 2909.330 934.690 2910.510 935.870 ;
        RECT 2907.730 933.090 2908.910 934.270 ;
        RECT 2909.330 933.090 2910.510 934.270 ;
        RECT 2907.730 754.690 2908.910 755.870 ;
        RECT 2909.330 754.690 2910.510 755.870 ;
        RECT 2907.730 753.090 2908.910 754.270 ;
        RECT 2909.330 753.090 2910.510 754.270 ;
        RECT 2907.730 574.690 2908.910 575.870 ;
        RECT 2909.330 574.690 2910.510 575.870 ;
        RECT 2907.730 573.090 2908.910 574.270 ;
        RECT 2909.330 573.090 2910.510 574.270 ;
        RECT 2907.730 394.690 2908.910 395.870 ;
        RECT 2909.330 394.690 2910.510 395.870 ;
        RECT 2907.730 393.090 2908.910 394.270 ;
        RECT 2909.330 393.090 2910.510 394.270 ;
        RECT 2907.730 214.690 2908.910 215.870 ;
        RECT 2909.330 214.690 2910.510 215.870 ;
        RECT 2907.730 213.090 2908.910 214.270 ;
        RECT 2909.330 213.090 2910.510 214.270 ;
        RECT 2907.730 34.690 2908.910 35.870 ;
        RECT 2909.330 34.690 2910.510 35.870 ;
        RECT 2907.730 33.090 2908.910 34.270 ;
        RECT 2909.330 33.090 2910.510 34.270 ;
        RECT 2907.730 -12.510 2908.910 -11.330 ;
        RECT 2909.330 -12.510 2910.510 -11.330 ;
        RECT 2907.730 -14.110 2908.910 -12.930 ;
        RECT 2909.330 -14.110 2910.510 -12.930 ;
        RECT 2936.310 3532.610 2937.490 3533.790 ;
        RECT 2937.910 3532.610 2939.090 3533.790 ;
        RECT 2936.310 3531.010 2937.490 3532.190 ;
        RECT 2937.910 3531.010 2939.090 3532.190 ;
        RECT 2936.310 3454.690 2937.490 3455.870 ;
        RECT 2937.910 3454.690 2939.090 3455.870 ;
        RECT 2936.310 3453.090 2937.490 3454.270 ;
        RECT 2937.910 3453.090 2939.090 3454.270 ;
        RECT 2936.310 3274.690 2937.490 3275.870 ;
        RECT 2937.910 3274.690 2939.090 3275.870 ;
        RECT 2936.310 3273.090 2937.490 3274.270 ;
        RECT 2937.910 3273.090 2939.090 3274.270 ;
        RECT 2936.310 3094.690 2937.490 3095.870 ;
        RECT 2937.910 3094.690 2939.090 3095.870 ;
        RECT 2936.310 3093.090 2937.490 3094.270 ;
        RECT 2937.910 3093.090 2939.090 3094.270 ;
        RECT 2936.310 2914.690 2937.490 2915.870 ;
        RECT 2937.910 2914.690 2939.090 2915.870 ;
        RECT 2936.310 2913.090 2937.490 2914.270 ;
        RECT 2937.910 2913.090 2939.090 2914.270 ;
        RECT 2936.310 2734.690 2937.490 2735.870 ;
        RECT 2937.910 2734.690 2939.090 2735.870 ;
        RECT 2936.310 2733.090 2937.490 2734.270 ;
        RECT 2937.910 2733.090 2939.090 2734.270 ;
        RECT 2936.310 2554.690 2937.490 2555.870 ;
        RECT 2937.910 2554.690 2939.090 2555.870 ;
        RECT 2936.310 2553.090 2937.490 2554.270 ;
        RECT 2937.910 2553.090 2939.090 2554.270 ;
        RECT 2936.310 2374.690 2937.490 2375.870 ;
        RECT 2937.910 2374.690 2939.090 2375.870 ;
        RECT 2936.310 2373.090 2937.490 2374.270 ;
        RECT 2937.910 2373.090 2939.090 2374.270 ;
        RECT 2936.310 2194.690 2937.490 2195.870 ;
        RECT 2937.910 2194.690 2939.090 2195.870 ;
        RECT 2936.310 2193.090 2937.490 2194.270 ;
        RECT 2937.910 2193.090 2939.090 2194.270 ;
        RECT 2936.310 2014.690 2937.490 2015.870 ;
        RECT 2937.910 2014.690 2939.090 2015.870 ;
        RECT 2936.310 2013.090 2937.490 2014.270 ;
        RECT 2937.910 2013.090 2939.090 2014.270 ;
        RECT 2936.310 1834.690 2937.490 1835.870 ;
        RECT 2937.910 1834.690 2939.090 1835.870 ;
        RECT 2936.310 1833.090 2937.490 1834.270 ;
        RECT 2937.910 1833.090 2939.090 1834.270 ;
        RECT 2936.310 1654.690 2937.490 1655.870 ;
        RECT 2937.910 1654.690 2939.090 1655.870 ;
        RECT 2936.310 1653.090 2937.490 1654.270 ;
        RECT 2937.910 1653.090 2939.090 1654.270 ;
        RECT 2936.310 1474.690 2937.490 1475.870 ;
        RECT 2937.910 1474.690 2939.090 1475.870 ;
        RECT 2936.310 1473.090 2937.490 1474.270 ;
        RECT 2937.910 1473.090 2939.090 1474.270 ;
        RECT 2936.310 1294.690 2937.490 1295.870 ;
        RECT 2937.910 1294.690 2939.090 1295.870 ;
        RECT 2936.310 1293.090 2937.490 1294.270 ;
        RECT 2937.910 1293.090 2939.090 1294.270 ;
        RECT 2936.310 1114.690 2937.490 1115.870 ;
        RECT 2937.910 1114.690 2939.090 1115.870 ;
        RECT 2936.310 1113.090 2937.490 1114.270 ;
        RECT 2937.910 1113.090 2939.090 1114.270 ;
        RECT 2936.310 934.690 2937.490 935.870 ;
        RECT 2937.910 934.690 2939.090 935.870 ;
        RECT 2936.310 933.090 2937.490 934.270 ;
        RECT 2937.910 933.090 2939.090 934.270 ;
        RECT 2936.310 754.690 2937.490 755.870 ;
        RECT 2937.910 754.690 2939.090 755.870 ;
        RECT 2936.310 753.090 2937.490 754.270 ;
        RECT 2937.910 753.090 2939.090 754.270 ;
        RECT 2936.310 574.690 2937.490 575.870 ;
        RECT 2937.910 574.690 2939.090 575.870 ;
        RECT 2936.310 573.090 2937.490 574.270 ;
        RECT 2937.910 573.090 2939.090 574.270 ;
        RECT 2936.310 394.690 2937.490 395.870 ;
        RECT 2937.910 394.690 2939.090 395.870 ;
        RECT 2936.310 393.090 2937.490 394.270 ;
        RECT 2937.910 393.090 2939.090 394.270 ;
        RECT 2936.310 214.690 2937.490 215.870 ;
        RECT 2937.910 214.690 2939.090 215.870 ;
        RECT 2936.310 213.090 2937.490 214.270 ;
        RECT 2937.910 213.090 2939.090 214.270 ;
        RECT 2936.310 34.690 2937.490 35.870 ;
        RECT 2937.910 34.690 2939.090 35.870 ;
        RECT 2936.310 33.090 2937.490 34.270 ;
        RECT 2937.910 33.090 2939.090 34.270 ;
        RECT 2936.310 -12.510 2937.490 -11.330 ;
        RECT 2937.910 -12.510 2939.090 -11.330 ;
        RECT 2936.310 -14.110 2937.490 -12.930 ;
        RECT 2937.910 -14.110 2939.090 -12.930 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
        RECT -24.430 932.930 2944.050 936.030 ;
        RECT -24.430 752.930 2944.050 756.030 ;
        RECT -24.430 572.930 2944.050 576.030 ;
        RECT -24.430 392.930 2944.050 396.030 ;
        RECT -24.430 212.930 2944.050 216.030 ;
        RECT -24.430 32.930 2944.050 36.030 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
        RECT 226.170 1010.000 229.270 3548.350 ;
        RECT 406.170 1010.000 409.270 3548.350 ;
        RECT 586.170 1010.000 589.270 3548.350 ;
        RECT 766.170 1010.000 769.270 3548.350 ;
        RECT 946.170 1010.000 949.270 3548.350 ;
        RECT 226.170 -28.670 229.270 390.000 ;
        RECT 406.170 -28.670 409.270 390.000 ;
        RECT 586.170 -28.670 589.270 390.000 ;
        RECT 766.170 -28.670 769.270 390.000 ;
        RECT 946.170 -28.670 949.270 390.000 ;
        RECT 1126.170 -28.670 1129.270 3548.350 ;
        RECT 1306.170 -28.670 1309.270 3548.350 ;
        RECT 1486.170 -28.670 1489.270 3548.350 ;
        RECT 1666.170 -28.670 1669.270 3548.350 ;
        RECT 1846.170 -28.670 1849.270 3548.350 ;
        RECT 2026.170 -28.670 2029.270 3548.350 ;
        RECT 2206.170 -28.670 2209.270 3548.350 ;
        RECT 2386.170 -28.670 2389.270 3548.350 ;
        RECT 2566.170 -28.670 2569.270 3548.350 ;
        RECT 2746.170 -28.670 2749.270 3548.350 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER via4 ;
        RECT -29.070 3542.210 -27.890 3543.390 ;
        RECT -27.470 3542.210 -26.290 3543.390 ;
        RECT -29.070 3540.610 -27.890 3541.790 ;
        RECT -27.470 3540.610 -26.290 3541.790 ;
        RECT -29.070 3473.290 -27.890 3474.470 ;
        RECT -27.470 3473.290 -26.290 3474.470 ;
        RECT -29.070 3471.690 -27.890 3472.870 ;
        RECT -27.470 3471.690 -26.290 3472.870 ;
        RECT -29.070 3293.290 -27.890 3294.470 ;
        RECT -27.470 3293.290 -26.290 3294.470 ;
        RECT -29.070 3291.690 -27.890 3292.870 ;
        RECT -27.470 3291.690 -26.290 3292.870 ;
        RECT -29.070 3113.290 -27.890 3114.470 ;
        RECT -27.470 3113.290 -26.290 3114.470 ;
        RECT -29.070 3111.690 -27.890 3112.870 ;
        RECT -27.470 3111.690 -26.290 3112.870 ;
        RECT -29.070 2933.290 -27.890 2934.470 ;
        RECT -27.470 2933.290 -26.290 2934.470 ;
        RECT -29.070 2931.690 -27.890 2932.870 ;
        RECT -27.470 2931.690 -26.290 2932.870 ;
        RECT -29.070 2753.290 -27.890 2754.470 ;
        RECT -27.470 2753.290 -26.290 2754.470 ;
        RECT -29.070 2751.690 -27.890 2752.870 ;
        RECT -27.470 2751.690 -26.290 2752.870 ;
        RECT -29.070 2573.290 -27.890 2574.470 ;
        RECT -27.470 2573.290 -26.290 2574.470 ;
        RECT -29.070 2571.690 -27.890 2572.870 ;
        RECT -27.470 2571.690 -26.290 2572.870 ;
        RECT -29.070 2393.290 -27.890 2394.470 ;
        RECT -27.470 2393.290 -26.290 2394.470 ;
        RECT -29.070 2391.690 -27.890 2392.870 ;
        RECT -27.470 2391.690 -26.290 2392.870 ;
        RECT -29.070 2213.290 -27.890 2214.470 ;
        RECT -27.470 2213.290 -26.290 2214.470 ;
        RECT -29.070 2211.690 -27.890 2212.870 ;
        RECT -27.470 2211.690 -26.290 2212.870 ;
        RECT -29.070 2033.290 -27.890 2034.470 ;
        RECT -27.470 2033.290 -26.290 2034.470 ;
        RECT -29.070 2031.690 -27.890 2032.870 ;
        RECT -27.470 2031.690 -26.290 2032.870 ;
        RECT -29.070 1853.290 -27.890 1854.470 ;
        RECT -27.470 1853.290 -26.290 1854.470 ;
        RECT -29.070 1851.690 -27.890 1852.870 ;
        RECT -27.470 1851.690 -26.290 1852.870 ;
        RECT -29.070 1673.290 -27.890 1674.470 ;
        RECT -27.470 1673.290 -26.290 1674.470 ;
        RECT -29.070 1671.690 -27.890 1672.870 ;
        RECT -27.470 1671.690 -26.290 1672.870 ;
        RECT -29.070 1493.290 -27.890 1494.470 ;
        RECT -27.470 1493.290 -26.290 1494.470 ;
        RECT -29.070 1491.690 -27.890 1492.870 ;
        RECT -27.470 1491.690 -26.290 1492.870 ;
        RECT -29.070 1313.290 -27.890 1314.470 ;
        RECT -27.470 1313.290 -26.290 1314.470 ;
        RECT -29.070 1311.690 -27.890 1312.870 ;
        RECT -27.470 1311.690 -26.290 1312.870 ;
        RECT -29.070 1133.290 -27.890 1134.470 ;
        RECT -27.470 1133.290 -26.290 1134.470 ;
        RECT -29.070 1131.690 -27.890 1132.870 ;
        RECT -27.470 1131.690 -26.290 1132.870 ;
        RECT -29.070 953.290 -27.890 954.470 ;
        RECT -27.470 953.290 -26.290 954.470 ;
        RECT -29.070 951.690 -27.890 952.870 ;
        RECT -27.470 951.690 -26.290 952.870 ;
        RECT -29.070 773.290 -27.890 774.470 ;
        RECT -27.470 773.290 -26.290 774.470 ;
        RECT -29.070 771.690 -27.890 772.870 ;
        RECT -27.470 771.690 -26.290 772.870 ;
        RECT -29.070 593.290 -27.890 594.470 ;
        RECT -27.470 593.290 -26.290 594.470 ;
        RECT -29.070 591.690 -27.890 592.870 ;
        RECT -27.470 591.690 -26.290 592.870 ;
        RECT -29.070 413.290 -27.890 414.470 ;
        RECT -27.470 413.290 -26.290 414.470 ;
        RECT -29.070 411.690 -27.890 412.870 ;
        RECT -27.470 411.690 -26.290 412.870 ;
        RECT -29.070 233.290 -27.890 234.470 ;
        RECT -27.470 233.290 -26.290 234.470 ;
        RECT -29.070 231.690 -27.890 232.870 ;
        RECT -27.470 231.690 -26.290 232.870 ;
        RECT -29.070 53.290 -27.890 54.470 ;
        RECT -27.470 53.290 -26.290 54.470 ;
        RECT -29.070 51.690 -27.890 52.870 ;
        RECT -27.470 51.690 -26.290 52.870 ;
        RECT -29.070 -22.110 -27.890 -20.930 ;
        RECT -27.470 -22.110 -26.290 -20.930 ;
        RECT -29.070 -23.710 -27.890 -22.530 ;
        RECT -27.470 -23.710 -26.290 -22.530 ;
        RECT 46.330 3542.210 47.510 3543.390 ;
        RECT 47.930 3542.210 49.110 3543.390 ;
        RECT 46.330 3540.610 47.510 3541.790 ;
        RECT 47.930 3540.610 49.110 3541.790 ;
        RECT 46.330 3473.290 47.510 3474.470 ;
        RECT 47.930 3473.290 49.110 3474.470 ;
        RECT 46.330 3471.690 47.510 3472.870 ;
        RECT 47.930 3471.690 49.110 3472.870 ;
        RECT 46.330 3293.290 47.510 3294.470 ;
        RECT 47.930 3293.290 49.110 3294.470 ;
        RECT 46.330 3291.690 47.510 3292.870 ;
        RECT 47.930 3291.690 49.110 3292.870 ;
        RECT 46.330 3113.290 47.510 3114.470 ;
        RECT 47.930 3113.290 49.110 3114.470 ;
        RECT 46.330 3111.690 47.510 3112.870 ;
        RECT 47.930 3111.690 49.110 3112.870 ;
        RECT 46.330 2933.290 47.510 2934.470 ;
        RECT 47.930 2933.290 49.110 2934.470 ;
        RECT 46.330 2931.690 47.510 2932.870 ;
        RECT 47.930 2931.690 49.110 2932.870 ;
        RECT 46.330 2753.290 47.510 2754.470 ;
        RECT 47.930 2753.290 49.110 2754.470 ;
        RECT 46.330 2751.690 47.510 2752.870 ;
        RECT 47.930 2751.690 49.110 2752.870 ;
        RECT 46.330 2573.290 47.510 2574.470 ;
        RECT 47.930 2573.290 49.110 2574.470 ;
        RECT 46.330 2571.690 47.510 2572.870 ;
        RECT 47.930 2571.690 49.110 2572.870 ;
        RECT 46.330 2393.290 47.510 2394.470 ;
        RECT 47.930 2393.290 49.110 2394.470 ;
        RECT 46.330 2391.690 47.510 2392.870 ;
        RECT 47.930 2391.690 49.110 2392.870 ;
        RECT 46.330 2213.290 47.510 2214.470 ;
        RECT 47.930 2213.290 49.110 2214.470 ;
        RECT 46.330 2211.690 47.510 2212.870 ;
        RECT 47.930 2211.690 49.110 2212.870 ;
        RECT 46.330 2033.290 47.510 2034.470 ;
        RECT 47.930 2033.290 49.110 2034.470 ;
        RECT 46.330 2031.690 47.510 2032.870 ;
        RECT 47.930 2031.690 49.110 2032.870 ;
        RECT 46.330 1853.290 47.510 1854.470 ;
        RECT 47.930 1853.290 49.110 1854.470 ;
        RECT 46.330 1851.690 47.510 1852.870 ;
        RECT 47.930 1851.690 49.110 1852.870 ;
        RECT 46.330 1673.290 47.510 1674.470 ;
        RECT 47.930 1673.290 49.110 1674.470 ;
        RECT 46.330 1671.690 47.510 1672.870 ;
        RECT 47.930 1671.690 49.110 1672.870 ;
        RECT 46.330 1493.290 47.510 1494.470 ;
        RECT 47.930 1493.290 49.110 1494.470 ;
        RECT 46.330 1491.690 47.510 1492.870 ;
        RECT 47.930 1491.690 49.110 1492.870 ;
        RECT 46.330 1313.290 47.510 1314.470 ;
        RECT 47.930 1313.290 49.110 1314.470 ;
        RECT 46.330 1311.690 47.510 1312.870 ;
        RECT 47.930 1311.690 49.110 1312.870 ;
        RECT 46.330 1133.290 47.510 1134.470 ;
        RECT 47.930 1133.290 49.110 1134.470 ;
        RECT 46.330 1131.690 47.510 1132.870 ;
        RECT 47.930 1131.690 49.110 1132.870 ;
        RECT 226.330 3542.210 227.510 3543.390 ;
        RECT 227.930 3542.210 229.110 3543.390 ;
        RECT 226.330 3540.610 227.510 3541.790 ;
        RECT 227.930 3540.610 229.110 3541.790 ;
        RECT 226.330 3473.290 227.510 3474.470 ;
        RECT 227.930 3473.290 229.110 3474.470 ;
        RECT 226.330 3471.690 227.510 3472.870 ;
        RECT 227.930 3471.690 229.110 3472.870 ;
        RECT 226.330 3293.290 227.510 3294.470 ;
        RECT 227.930 3293.290 229.110 3294.470 ;
        RECT 226.330 3291.690 227.510 3292.870 ;
        RECT 227.930 3291.690 229.110 3292.870 ;
        RECT 226.330 3113.290 227.510 3114.470 ;
        RECT 227.930 3113.290 229.110 3114.470 ;
        RECT 226.330 3111.690 227.510 3112.870 ;
        RECT 227.930 3111.690 229.110 3112.870 ;
        RECT 226.330 2933.290 227.510 2934.470 ;
        RECT 227.930 2933.290 229.110 2934.470 ;
        RECT 226.330 2931.690 227.510 2932.870 ;
        RECT 227.930 2931.690 229.110 2932.870 ;
        RECT 226.330 2753.290 227.510 2754.470 ;
        RECT 227.930 2753.290 229.110 2754.470 ;
        RECT 226.330 2751.690 227.510 2752.870 ;
        RECT 227.930 2751.690 229.110 2752.870 ;
        RECT 226.330 2573.290 227.510 2574.470 ;
        RECT 227.930 2573.290 229.110 2574.470 ;
        RECT 226.330 2571.690 227.510 2572.870 ;
        RECT 227.930 2571.690 229.110 2572.870 ;
        RECT 226.330 2393.290 227.510 2394.470 ;
        RECT 227.930 2393.290 229.110 2394.470 ;
        RECT 226.330 2391.690 227.510 2392.870 ;
        RECT 227.930 2391.690 229.110 2392.870 ;
        RECT 226.330 2213.290 227.510 2214.470 ;
        RECT 227.930 2213.290 229.110 2214.470 ;
        RECT 226.330 2211.690 227.510 2212.870 ;
        RECT 227.930 2211.690 229.110 2212.870 ;
        RECT 226.330 2033.290 227.510 2034.470 ;
        RECT 227.930 2033.290 229.110 2034.470 ;
        RECT 226.330 2031.690 227.510 2032.870 ;
        RECT 227.930 2031.690 229.110 2032.870 ;
        RECT 226.330 1853.290 227.510 1854.470 ;
        RECT 227.930 1853.290 229.110 1854.470 ;
        RECT 226.330 1851.690 227.510 1852.870 ;
        RECT 227.930 1851.690 229.110 1852.870 ;
        RECT 226.330 1673.290 227.510 1674.470 ;
        RECT 227.930 1673.290 229.110 1674.470 ;
        RECT 226.330 1671.690 227.510 1672.870 ;
        RECT 227.930 1671.690 229.110 1672.870 ;
        RECT 226.330 1493.290 227.510 1494.470 ;
        RECT 227.930 1493.290 229.110 1494.470 ;
        RECT 226.330 1491.690 227.510 1492.870 ;
        RECT 227.930 1491.690 229.110 1492.870 ;
        RECT 226.330 1313.290 227.510 1314.470 ;
        RECT 227.930 1313.290 229.110 1314.470 ;
        RECT 226.330 1311.690 227.510 1312.870 ;
        RECT 227.930 1311.690 229.110 1312.870 ;
        RECT 226.330 1133.290 227.510 1134.470 ;
        RECT 227.930 1133.290 229.110 1134.470 ;
        RECT 226.330 1131.690 227.510 1132.870 ;
        RECT 227.930 1131.690 229.110 1132.870 ;
        RECT 406.330 3542.210 407.510 3543.390 ;
        RECT 407.930 3542.210 409.110 3543.390 ;
        RECT 406.330 3540.610 407.510 3541.790 ;
        RECT 407.930 3540.610 409.110 3541.790 ;
        RECT 406.330 3473.290 407.510 3474.470 ;
        RECT 407.930 3473.290 409.110 3474.470 ;
        RECT 406.330 3471.690 407.510 3472.870 ;
        RECT 407.930 3471.690 409.110 3472.870 ;
        RECT 406.330 3293.290 407.510 3294.470 ;
        RECT 407.930 3293.290 409.110 3294.470 ;
        RECT 406.330 3291.690 407.510 3292.870 ;
        RECT 407.930 3291.690 409.110 3292.870 ;
        RECT 406.330 3113.290 407.510 3114.470 ;
        RECT 407.930 3113.290 409.110 3114.470 ;
        RECT 406.330 3111.690 407.510 3112.870 ;
        RECT 407.930 3111.690 409.110 3112.870 ;
        RECT 406.330 2933.290 407.510 2934.470 ;
        RECT 407.930 2933.290 409.110 2934.470 ;
        RECT 406.330 2931.690 407.510 2932.870 ;
        RECT 407.930 2931.690 409.110 2932.870 ;
        RECT 406.330 2753.290 407.510 2754.470 ;
        RECT 407.930 2753.290 409.110 2754.470 ;
        RECT 406.330 2751.690 407.510 2752.870 ;
        RECT 407.930 2751.690 409.110 2752.870 ;
        RECT 406.330 2573.290 407.510 2574.470 ;
        RECT 407.930 2573.290 409.110 2574.470 ;
        RECT 406.330 2571.690 407.510 2572.870 ;
        RECT 407.930 2571.690 409.110 2572.870 ;
        RECT 406.330 2393.290 407.510 2394.470 ;
        RECT 407.930 2393.290 409.110 2394.470 ;
        RECT 406.330 2391.690 407.510 2392.870 ;
        RECT 407.930 2391.690 409.110 2392.870 ;
        RECT 406.330 2213.290 407.510 2214.470 ;
        RECT 407.930 2213.290 409.110 2214.470 ;
        RECT 406.330 2211.690 407.510 2212.870 ;
        RECT 407.930 2211.690 409.110 2212.870 ;
        RECT 406.330 2033.290 407.510 2034.470 ;
        RECT 407.930 2033.290 409.110 2034.470 ;
        RECT 406.330 2031.690 407.510 2032.870 ;
        RECT 407.930 2031.690 409.110 2032.870 ;
        RECT 406.330 1853.290 407.510 1854.470 ;
        RECT 407.930 1853.290 409.110 1854.470 ;
        RECT 406.330 1851.690 407.510 1852.870 ;
        RECT 407.930 1851.690 409.110 1852.870 ;
        RECT 406.330 1673.290 407.510 1674.470 ;
        RECT 407.930 1673.290 409.110 1674.470 ;
        RECT 406.330 1671.690 407.510 1672.870 ;
        RECT 407.930 1671.690 409.110 1672.870 ;
        RECT 406.330 1493.290 407.510 1494.470 ;
        RECT 407.930 1493.290 409.110 1494.470 ;
        RECT 406.330 1491.690 407.510 1492.870 ;
        RECT 407.930 1491.690 409.110 1492.870 ;
        RECT 406.330 1313.290 407.510 1314.470 ;
        RECT 407.930 1313.290 409.110 1314.470 ;
        RECT 406.330 1311.690 407.510 1312.870 ;
        RECT 407.930 1311.690 409.110 1312.870 ;
        RECT 406.330 1133.290 407.510 1134.470 ;
        RECT 407.930 1133.290 409.110 1134.470 ;
        RECT 406.330 1131.690 407.510 1132.870 ;
        RECT 407.930 1131.690 409.110 1132.870 ;
        RECT 586.330 3542.210 587.510 3543.390 ;
        RECT 587.930 3542.210 589.110 3543.390 ;
        RECT 586.330 3540.610 587.510 3541.790 ;
        RECT 587.930 3540.610 589.110 3541.790 ;
        RECT 586.330 3473.290 587.510 3474.470 ;
        RECT 587.930 3473.290 589.110 3474.470 ;
        RECT 586.330 3471.690 587.510 3472.870 ;
        RECT 587.930 3471.690 589.110 3472.870 ;
        RECT 586.330 3293.290 587.510 3294.470 ;
        RECT 587.930 3293.290 589.110 3294.470 ;
        RECT 586.330 3291.690 587.510 3292.870 ;
        RECT 587.930 3291.690 589.110 3292.870 ;
        RECT 586.330 3113.290 587.510 3114.470 ;
        RECT 587.930 3113.290 589.110 3114.470 ;
        RECT 586.330 3111.690 587.510 3112.870 ;
        RECT 587.930 3111.690 589.110 3112.870 ;
        RECT 586.330 2933.290 587.510 2934.470 ;
        RECT 587.930 2933.290 589.110 2934.470 ;
        RECT 586.330 2931.690 587.510 2932.870 ;
        RECT 587.930 2931.690 589.110 2932.870 ;
        RECT 586.330 2753.290 587.510 2754.470 ;
        RECT 587.930 2753.290 589.110 2754.470 ;
        RECT 586.330 2751.690 587.510 2752.870 ;
        RECT 587.930 2751.690 589.110 2752.870 ;
        RECT 586.330 2573.290 587.510 2574.470 ;
        RECT 587.930 2573.290 589.110 2574.470 ;
        RECT 586.330 2571.690 587.510 2572.870 ;
        RECT 587.930 2571.690 589.110 2572.870 ;
        RECT 586.330 2393.290 587.510 2394.470 ;
        RECT 587.930 2393.290 589.110 2394.470 ;
        RECT 586.330 2391.690 587.510 2392.870 ;
        RECT 587.930 2391.690 589.110 2392.870 ;
        RECT 586.330 2213.290 587.510 2214.470 ;
        RECT 587.930 2213.290 589.110 2214.470 ;
        RECT 586.330 2211.690 587.510 2212.870 ;
        RECT 587.930 2211.690 589.110 2212.870 ;
        RECT 586.330 2033.290 587.510 2034.470 ;
        RECT 587.930 2033.290 589.110 2034.470 ;
        RECT 586.330 2031.690 587.510 2032.870 ;
        RECT 587.930 2031.690 589.110 2032.870 ;
        RECT 586.330 1853.290 587.510 1854.470 ;
        RECT 587.930 1853.290 589.110 1854.470 ;
        RECT 586.330 1851.690 587.510 1852.870 ;
        RECT 587.930 1851.690 589.110 1852.870 ;
        RECT 586.330 1673.290 587.510 1674.470 ;
        RECT 587.930 1673.290 589.110 1674.470 ;
        RECT 586.330 1671.690 587.510 1672.870 ;
        RECT 587.930 1671.690 589.110 1672.870 ;
        RECT 586.330 1493.290 587.510 1494.470 ;
        RECT 587.930 1493.290 589.110 1494.470 ;
        RECT 586.330 1491.690 587.510 1492.870 ;
        RECT 587.930 1491.690 589.110 1492.870 ;
        RECT 586.330 1313.290 587.510 1314.470 ;
        RECT 587.930 1313.290 589.110 1314.470 ;
        RECT 586.330 1311.690 587.510 1312.870 ;
        RECT 587.930 1311.690 589.110 1312.870 ;
        RECT 586.330 1133.290 587.510 1134.470 ;
        RECT 587.930 1133.290 589.110 1134.470 ;
        RECT 586.330 1131.690 587.510 1132.870 ;
        RECT 587.930 1131.690 589.110 1132.870 ;
        RECT 766.330 3542.210 767.510 3543.390 ;
        RECT 767.930 3542.210 769.110 3543.390 ;
        RECT 766.330 3540.610 767.510 3541.790 ;
        RECT 767.930 3540.610 769.110 3541.790 ;
        RECT 766.330 3473.290 767.510 3474.470 ;
        RECT 767.930 3473.290 769.110 3474.470 ;
        RECT 766.330 3471.690 767.510 3472.870 ;
        RECT 767.930 3471.690 769.110 3472.870 ;
        RECT 766.330 3293.290 767.510 3294.470 ;
        RECT 767.930 3293.290 769.110 3294.470 ;
        RECT 766.330 3291.690 767.510 3292.870 ;
        RECT 767.930 3291.690 769.110 3292.870 ;
        RECT 766.330 3113.290 767.510 3114.470 ;
        RECT 767.930 3113.290 769.110 3114.470 ;
        RECT 766.330 3111.690 767.510 3112.870 ;
        RECT 767.930 3111.690 769.110 3112.870 ;
        RECT 766.330 2933.290 767.510 2934.470 ;
        RECT 767.930 2933.290 769.110 2934.470 ;
        RECT 766.330 2931.690 767.510 2932.870 ;
        RECT 767.930 2931.690 769.110 2932.870 ;
        RECT 766.330 2753.290 767.510 2754.470 ;
        RECT 767.930 2753.290 769.110 2754.470 ;
        RECT 766.330 2751.690 767.510 2752.870 ;
        RECT 767.930 2751.690 769.110 2752.870 ;
        RECT 766.330 2573.290 767.510 2574.470 ;
        RECT 767.930 2573.290 769.110 2574.470 ;
        RECT 766.330 2571.690 767.510 2572.870 ;
        RECT 767.930 2571.690 769.110 2572.870 ;
        RECT 766.330 2393.290 767.510 2394.470 ;
        RECT 767.930 2393.290 769.110 2394.470 ;
        RECT 766.330 2391.690 767.510 2392.870 ;
        RECT 767.930 2391.690 769.110 2392.870 ;
        RECT 766.330 2213.290 767.510 2214.470 ;
        RECT 767.930 2213.290 769.110 2214.470 ;
        RECT 766.330 2211.690 767.510 2212.870 ;
        RECT 767.930 2211.690 769.110 2212.870 ;
        RECT 766.330 2033.290 767.510 2034.470 ;
        RECT 767.930 2033.290 769.110 2034.470 ;
        RECT 766.330 2031.690 767.510 2032.870 ;
        RECT 767.930 2031.690 769.110 2032.870 ;
        RECT 766.330 1853.290 767.510 1854.470 ;
        RECT 767.930 1853.290 769.110 1854.470 ;
        RECT 766.330 1851.690 767.510 1852.870 ;
        RECT 767.930 1851.690 769.110 1852.870 ;
        RECT 766.330 1673.290 767.510 1674.470 ;
        RECT 767.930 1673.290 769.110 1674.470 ;
        RECT 766.330 1671.690 767.510 1672.870 ;
        RECT 767.930 1671.690 769.110 1672.870 ;
        RECT 766.330 1493.290 767.510 1494.470 ;
        RECT 767.930 1493.290 769.110 1494.470 ;
        RECT 766.330 1491.690 767.510 1492.870 ;
        RECT 767.930 1491.690 769.110 1492.870 ;
        RECT 766.330 1313.290 767.510 1314.470 ;
        RECT 767.930 1313.290 769.110 1314.470 ;
        RECT 766.330 1311.690 767.510 1312.870 ;
        RECT 767.930 1311.690 769.110 1312.870 ;
        RECT 766.330 1133.290 767.510 1134.470 ;
        RECT 767.930 1133.290 769.110 1134.470 ;
        RECT 766.330 1131.690 767.510 1132.870 ;
        RECT 767.930 1131.690 769.110 1132.870 ;
        RECT 946.330 3542.210 947.510 3543.390 ;
        RECT 947.930 3542.210 949.110 3543.390 ;
        RECT 946.330 3540.610 947.510 3541.790 ;
        RECT 947.930 3540.610 949.110 3541.790 ;
        RECT 946.330 3473.290 947.510 3474.470 ;
        RECT 947.930 3473.290 949.110 3474.470 ;
        RECT 946.330 3471.690 947.510 3472.870 ;
        RECT 947.930 3471.690 949.110 3472.870 ;
        RECT 946.330 3293.290 947.510 3294.470 ;
        RECT 947.930 3293.290 949.110 3294.470 ;
        RECT 946.330 3291.690 947.510 3292.870 ;
        RECT 947.930 3291.690 949.110 3292.870 ;
        RECT 946.330 3113.290 947.510 3114.470 ;
        RECT 947.930 3113.290 949.110 3114.470 ;
        RECT 946.330 3111.690 947.510 3112.870 ;
        RECT 947.930 3111.690 949.110 3112.870 ;
        RECT 946.330 2933.290 947.510 2934.470 ;
        RECT 947.930 2933.290 949.110 2934.470 ;
        RECT 946.330 2931.690 947.510 2932.870 ;
        RECT 947.930 2931.690 949.110 2932.870 ;
        RECT 946.330 2753.290 947.510 2754.470 ;
        RECT 947.930 2753.290 949.110 2754.470 ;
        RECT 946.330 2751.690 947.510 2752.870 ;
        RECT 947.930 2751.690 949.110 2752.870 ;
        RECT 946.330 2573.290 947.510 2574.470 ;
        RECT 947.930 2573.290 949.110 2574.470 ;
        RECT 946.330 2571.690 947.510 2572.870 ;
        RECT 947.930 2571.690 949.110 2572.870 ;
        RECT 946.330 2393.290 947.510 2394.470 ;
        RECT 947.930 2393.290 949.110 2394.470 ;
        RECT 946.330 2391.690 947.510 2392.870 ;
        RECT 947.930 2391.690 949.110 2392.870 ;
        RECT 946.330 2213.290 947.510 2214.470 ;
        RECT 947.930 2213.290 949.110 2214.470 ;
        RECT 946.330 2211.690 947.510 2212.870 ;
        RECT 947.930 2211.690 949.110 2212.870 ;
        RECT 946.330 2033.290 947.510 2034.470 ;
        RECT 947.930 2033.290 949.110 2034.470 ;
        RECT 946.330 2031.690 947.510 2032.870 ;
        RECT 947.930 2031.690 949.110 2032.870 ;
        RECT 946.330 1853.290 947.510 1854.470 ;
        RECT 947.930 1853.290 949.110 1854.470 ;
        RECT 946.330 1851.690 947.510 1852.870 ;
        RECT 947.930 1851.690 949.110 1852.870 ;
        RECT 946.330 1673.290 947.510 1674.470 ;
        RECT 947.930 1673.290 949.110 1674.470 ;
        RECT 946.330 1671.690 947.510 1672.870 ;
        RECT 947.930 1671.690 949.110 1672.870 ;
        RECT 946.330 1493.290 947.510 1494.470 ;
        RECT 947.930 1493.290 949.110 1494.470 ;
        RECT 946.330 1491.690 947.510 1492.870 ;
        RECT 947.930 1491.690 949.110 1492.870 ;
        RECT 946.330 1313.290 947.510 1314.470 ;
        RECT 947.930 1313.290 949.110 1314.470 ;
        RECT 946.330 1311.690 947.510 1312.870 ;
        RECT 947.930 1311.690 949.110 1312.870 ;
        RECT 946.330 1133.290 947.510 1134.470 ;
        RECT 947.930 1133.290 949.110 1134.470 ;
        RECT 946.330 1131.690 947.510 1132.870 ;
        RECT 947.930 1131.690 949.110 1132.870 ;
        RECT 1126.330 3542.210 1127.510 3543.390 ;
        RECT 1127.930 3542.210 1129.110 3543.390 ;
        RECT 1126.330 3540.610 1127.510 3541.790 ;
        RECT 1127.930 3540.610 1129.110 3541.790 ;
        RECT 1126.330 3473.290 1127.510 3474.470 ;
        RECT 1127.930 3473.290 1129.110 3474.470 ;
        RECT 1126.330 3471.690 1127.510 3472.870 ;
        RECT 1127.930 3471.690 1129.110 3472.870 ;
        RECT 1126.330 3293.290 1127.510 3294.470 ;
        RECT 1127.930 3293.290 1129.110 3294.470 ;
        RECT 1126.330 3291.690 1127.510 3292.870 ;
        RECT 1127.930 3291.690 1129.110 3292.870 ;
        RECT 1126.330 3113.290 1127.510 3114.470 ;
        RECT 1127.930 3113.290 1129.110 3114.470 ;
        RECT 1126.330 3111.690 1127.510 3112.870 ;
        RECT 1127.930 3111.690 1129.110 3112.870 ;
        RECT 1126.330 2933.290 1127.510 2934.470 ;
        RECT 1127.930 2933.290 1129.110 2934.470 ;
        RECT 1126.330 2931.690 1127.510 2932.870 ;
        RECT 1127.930 2931.690 1129.110 2932.870 ;
        RECT 1126.330 2753.290 1127.510 2754.470 ;
        RECT 1127.930 2753.290 1129.110 2754.470 ;
        RECT 1126.330 2751.690 1127.510 2752.870 ;
        RECT 1127.930 2751.690 1129.110 2752.870 ;
        RECT 1126.330 2573.290 1127.510 2574.470 ;
        RECT 1127.930 2573.290 1129.110 2574.470 ;
        RECT 1126.330 2571.690 1127.510 2572.870 ;
        RECT 1127.930 2571.690 1129.110 2572.870 ;
        RECT 1126.330 2393.290 1127.510 2394.470 ;
        RECT 1127.930 2393.290 1129.110 2394.470 ;
        RECT 1126.330 2391.690 1127.510 2392.870 ;
        RECT 1127.930 2391.690 1129.110 2392.870 ;
        RECT 1126.330 2213.290 1127.510 2214.470 ;
        RECT 1127.930 2213.290 1129.110 2214.470 ;
        RECT 1126.330 2211.690 1127.510 2212.870 ;
        RECT 1127.930 2211.690 1129.110 2212.870 ;
        RECT 1126.330 2033.290 1127.510 2034.470 ;
        RECT 1127.930 2033.290 1129.110 2034.470 ;
        RECT 1126.330 2031.690 1127.510 2032.870 ;
        RECT 1127.930 2031.690 1129.110 2032.870 ;
        RECT 1126.330 1853.290 1127.510 1854.470 ;
        RECT 1127.930 1853.290 1129.110 1854.470 ;
        RECT 1126.330 1851.690 1127.510 1852.870 ;
        RECT 1127.930 1851.690 1129.110 1852.870 ;
        RECT 1126.330 1673.290 1127.510 1674.470 ;
        RECT 1127.930 1673.290 1129.110 1674.470 ;
        RECT 1126.330 1671.690 1127.510 1672.870 ;
        RECT 1127.930 1671.690 1129.110 1672.870 ;
        RECT 1126.330 1493.290 1127.510 1494.470 ;
        RECT 1127.930 1493.290 1129.110 1494.470 ;
        RECT 1126.330 1491.690 1127.510 1492.870 ;
        RECT 1127.930 1491.690 1129.110 1492.870 ;
        RECT 1126.330 1313.290 1127.510 1314.470 ;
        RECT 1127.930 1313.290 1129.110 1314.470 ;
        RECT 1126.330 1311.690 1127.510 1312.870 ;
        RECT 1127.930 1311.690 1129.110 1312.870 ;
        RECT 1126.330 1133.290 1127.510 1134.470 ;
        RECT 1127.930 1133.290 1129.110 1134.470 ;
        RECT 1126.330 1131.690 1127.510 1132.870 ;
        RECT 1127.930 1131.690 1129.110 1132.870 ;
        RECT 46.330 953.290 47.510 954.470 ;
        RECT 47.930 953.290 49.110 954.470 ;
        RECT 46.330 951.690 47.510 952.870 ;
        RECT 47.930 951.690 49.110 952.870 ;
        RECT 46.330 773.290 47.510 774.470 ;
        RECT 47.930 773.290 49.110 774.470 ;
        RECT 46.330 771.690 47.510 772.870 ;
        RECT 47.930 771.690 49.110 772.870 ;
        RECT 46.330 593.290 47.510 594.470 ;
        RECT 47.930 593.290 49.110 594.470 ;
        RECT 46.330 591.690 47.510 592.870 ;
        RECT 47.930 591.690 49.110 592.870 ;
        RECT 46.330 413.290 47.510 414.470 ;
        RECT 47.930 413.290 49.110 414.470 ;
        RECT 46.330 411.690 47.510 412.870 ;
        RECT 47.930 411.690 49.110 412.870 ;
        RECT 1126.330 953.290 1127.510 954.470 ;
        RECT 1127.930 953.290 1129.110 954.470 ;
        RECT 1126.330 951.690 1127.510 952.870 ;
        RECT 1127.930 951.690 1129.110 952.870 ;
        RECT 1126.330 773.290 1127.510 774.470 ;
        RECT 1127.930 773.290 1129.110 774.470 ;
        RECT 1126.330 771.690 1127.510 772.870 ;
        RECT 1127.930 771.690 1129.110 772.870 ;
        RECT 1126.330 593.290 1127.510 594.470 ;
        RECT 1127.930 593.290 1129.110 594.470 ;
        RECT 1126.330 591.690 1127.510 592.870 ;
        RECT 1127.930 591.690 1129.110 592.870 ;
        RECT 1126.330 413.290 1127.510 414.470 ;
        RECT 1127.930 413.290 1129.110 414.470 ;
        RECT 1126.330 411.690 1127.510 412.870 ;
        RECT 1127.930 411.690 1129.110 412.870 ;
        RECT 46.330 233.290 47.510 234.470 ;
        RECT 47.930 233.290 49.110 234.470 ;
        RECT 46.330 231.690 47.510 232.870 ;
        RECT 47.930 231.690 49.110 232.870 ;
        RECT 46.330 53.290 47.510 54.470 ;
        RECT 47.930 53.290 49.110 54.470 ;
        RECT 46.330 51.690 47.510 52.870 ;
        RECT 47.930 51.690 49.110 52.870 ;
        RECT 46.330 -22.110 47.510 -20.930 ;
        RECT 47.930 -22.110 49.110 -20.930 ;
        RECT 46.330 -23.710 47.510 -22.530 ;
        RECT 47.930 -23.710 49.110 -22.530 ;
        RECT 226.330 233.290 227.510 234.470 ;
        RECT 227.930 233.290 229.110 234.470 ;
        RECT 226.330 231.690 227.510 232.870 ;
        RECT 227.930 231.690 229.110 232.870 ;
        RECT 226.330 53.290 227.510 54.470 ;
        RECT 227.930 53.290 229.110 54.470 ;
        RECT 226.330 51.690 227.510 52.870 ;
        RECT 227.930 51.690 229.110 52.870 ;
        RECT 226.330 -22.110 227.510 -20.930 ;
        RECT 227.930 -22.110 229.110 -20.930 ;
        RECT 226.330 -23.710 227.510 -22.530 ;
        RECT 227.930 -23.710 229.110 -22.530 ;
        RECT 406.330 233.290 407.510 234.470 ;
        RECT 407.930 233.290 409.110 234.470 ;
        RECT 406.330 231.690 407.510 232.870 ;
        RECT 407.930 231.690 409.110 232.870 ;
        RECT 406.330 53.290 407.510 54.470 ;
        RECT 407.930 53.290 409.110 54.470 ;
        RECT 406.330 51.690 407.510 52.870 ;
        RECT 407.930 51.690 409.110 52.870 ;
        RECT 406.330 -22.110 407.510 -20.930 ;
        RECT 407.930 -22.110 409.110 -20.930 ;
        RECT 406.330 -23.710 407.510 -22.530 ;
        RECT 407.930 -23.710 409.110 -22.530 ;
        RECT 586.330 233.290 587.510 234.470 ;
        RECT 587.930 233.290 589.110 234.470 ;
        RECT 586.330 231.690 587.510 232.870 ;
        RECT 587.930 231.690 589.110 232.870 ;
        RECT 586.330 53.290 587.510 54.470 ;
        RECT 587.930 53.290 589.110 54.470 ;
        RECT 586.330 51.690 587.510 52.870 ;
        RECT 587.930 51.690 589.110 52.870 ;
        RECT 586.330 -22.110 587.510 -20.930 ;
        RECT 587.930 -22.110 589.110 -20.930 ;
        RECT 586.330 -23.710 587.510 -22.530 ;
        RECT 587.930 -23.710 589.110 -22.530 ;
        RECT 766.330 233.290 767.510 234.470 ;
        RECT 767.930 233.290 769.110 234.470 ;
        RECT 766.330 231.690 767.510 232.870 ;
        RECT 767.930 231.690 769.110 232.870 ;
        RECT 766.330 53.290 767.510 54.470 ;
        RECT 767.930 53.290 769.110 54.470 ;
        RECT 766.330 51.690 767.510 52.870 ;
        RECT 767.930 51.690 769.110 52.870 ;
        RECT 766.330 -22.110 767.510 -20.930 ;
        RECT 767.930 -22.110 769.110 -20.930 ;
        RECT 766.330 -23.710 767.510 -22.530 ;
        RECT 767.930 -23.710 769.110 -22.530 ;
        RECT 946.330 233.290 947.510 234.470 ;
        RECT 947.930 233.290 949.110 234.470 ;
        RECT 946.330 231.690 947.510 232.870 ;
        RECT 947.930 231.690 949.110 232.870 ;
        RECT 946.330 53.290 947.510 54.470 ;
        RECT 947.930 53.290 949.110 54.470 ;
        RECT 946.330 51.690 947.510 52.870 ;
        RECT 947.930 51.690 949.110 52.870 ;
        RECT 946.330 -22.110 947.510 -20.930 ;
        RECT 947.930 -22.110 949.110 -20.930 ;
        RECT 946.330 -23.710 947.510 -22.530 ;
        RECT 947.930 -23.710 949.110 -22.530 ;
        RECT 1126.330 233.290 1127.510 234.470 ;
        RECT 1127.930 233.290 1129.110 234.470 ;
        RECT 1126.330 231.690 1127.510 232.870 ;
        RECT 1127.930 231.690 1129.110 232.870 ;
        RECT 1126.330 53.290 1127.510 54.470 ;
        RECT 1127.930 53.290 1129.110 54.470 ;
        RECT 1126.330 51.690 1127.510 52.870 ;
        RECT 1127.930 51.690 1129.110 52.870 ;
        RECT 1126.330 -22.110 1127.510 -20.930 ;
        RECT 1127.930 -22.110 1129.110 -20.930 ;
        RECT 1126.330 -23.710 1127.510 -22.530 ;
        RECT 1127.930 -23.710 1129.110 -22.530 ;
        RECT 1306.330 3542.210 1307.510 3543.390 ;
        RECT 1307.930 3542.210 1309.110 3543.390 ;
        RECT 1306.330 3540.610 1307.510 3541.790 ;
        RECT 1307.930 3540.610 1309.110 3541.790 ;
        RECT 1306.330 3473.290 1307.510 3474.470 ;
        RECT 1307.930 3473.290 1309.110 3474.470 ;
        RECT 1306.330 3471.690 1307.510 3472.870 ;
        RECT 1307.930 3471.690 1309.110 3472.870 ;
        RECT 1306.330 3293.290 1307.510 3294.470 ;
        RECT 1307.930 3293.290 1309.110 3294.470 ;
        RECT 1306.330 3291.690 1307.510 3292.870 ;
        RECT 1307.930 3291.690 1309.110 3292.870 ;
        RECT 1306.330 3113.290 1307.510 3114.470 ;
        RECT 1307.930 3113.290 1309.110 3114.470 ;
        RECT 1306.330 3111.690 1307.510 3112.870 ;
        RECT 1307.930 3111.690 1309.110 3112.870 ;
        RECT 1306.330 2933.290 1307.510 2934.470 ;
        RECT 1307.930 2933.290 1309.110 2934.470 ;
        RECT 1306.330 2931.690 1307.510 2932.870 ;
        RECT 1307.930 2931.690 1309.110 2932.870 ;
        RECT 1306.330 2753.290 1307.510 2754.470 ;
        RECT 1307.930 2753.290 1309.110 2754.470 ;
        RECT 1306.330 2751.690 1307.510 2752.870 ;
        RECT 1307.930 2751.690 1309.110 2752.870 ;
        RECT 1306.330 2573.290 1307.510 2574.470 ;
        RECT 1307.930 2573.290 1309.110 2574.470 ;
        RECT 1306.330 2571.690 1307.510 2572.870 ;
        RECT 1307.930 2571.690 1309.110 2572.870 ;
        RECT 1306.330 2393.290 1307.510 2394.470 ;
        RECT 1307.930 2393.290 1309.110 2394.470 ;
        RECT 1306.330 2391.690 1307.510 2392.870 ;
        RECT 1307.930 2391.690 1309.110 2392.870 ;
        RECT 1306.330 2213.290 1307.510 2214.470 ;
        RECT 1307.930 2213.290 1309.110 2214.470 ;
        RECT 1306.330 2211.690 1307.510 2212.870 ;
        RECT 1307.930 2211.690 1309.110 2212.870 ;
        RECT 1306.330 2033.290 1307.510 2034.470 ;
        RECT 1307.930 2033.290 1309.110 2034.470 ;
        RECT 1306.330 2031.690 1307.510 2032.870 ;
        RECT 1307.930 2031.690 1309.110 2032.870 ;
        RECT 1306.330 1853.290 1307.510 1854.470 ;
        RECT 1307.930 1853.290 1309.110 1854.470 ;
        RECT 1306.330 1851.690 1307.510 1852.870 ;
        RECT 1307.930 1851.690 1309.110 1852.870 ;
        RECT 1306.330 1673.290 1307.510 1674.470 ;
        RECT 1307.930 1673.290 1309.110 1674.470 ;
        RECT 1306.330 1671.690 1307.510 1672.870 ;
        RECT 1307.930 1671.690 1309.110 1672.870 ;
        RECT 1306.330 1493.290 1307.510 1494.470 ;
        RECT 1307.930 1493.290 1309.110 1494.470 ;
        RECT 1306.330 1491.690 1307.510 1492.870 ;
        RECT 1307.930 1491.690 1309.110 1492.870 ;
        RECT 1306.330 1313.290 1307.510 1314.470 ;
        RECT 1307.930 1313.290 1309.110 1314.470 ;
        RECT 1306.330 1311.690 1307.510 1312.870 ;
        RECT 1307.930 1311.690 1309.110 1312.870 ;
        RECT 1306.330 1133.290 1307.510 1134.470 ;
        RECT 1307.930 1133.290 1309.110 1134.470 ;
        RECT 1306.330 1131.690 1307.510 1132.870 ;
        RECT 1307.930 1131.690 1309.110 1132.870 ;
        RECT 1306.330 953.290 1307.510 954.470 ;
        RECT 1307.930 953.290 1309.110 954.470 ;
        RECT 1306.330 951.690 1307.510 952.870 ;
        RECT 1307.930 951.690 1309.110 952.870 ;
        RECT 1306.330 773.290 1307.510 774.470 ;
        RECT 1307.930 773.290 1309.110 774.470 ;
        RECT 1306.330 771.690 1307.510 772.870 ;
        RECT 1307.930 771.690 1309.110 772.870 ;
        RECT 1306.330 593.290 1307.510 594.470 ;
        RECT 1307.930 593.290 1309.110 594.470 ;
        RECT 1306.330 591.690 1307.510 592.870 ;
        RECT 1307.930 591.690 1309.110 592.870 ;
        RECT 1306.330 413.290 1307.510 414.470 ;
        RECT 1307.930 413.290 1309.110 414.470 ;
        RECT 1306.330 411.690 1307.510 412.870 ;
        RECT 1307.930 411.690 1309.110 412.870 ;
        RECT 1306.330 233.290 1307.510 234.470 ;
        RECT 1307.930 233.290 1309.110 234.470 ;
        RECT 1306.330 231.690 1307.510 232.870 ;
        RECT 1307.930 231.690 1309.110 232.870 ;
        RECT 1306.330 53.290 1307.510 54.470 ;
        RECT 1307.930 53.290 1309.110 54.470 ;
        RECT 1306.330 51.690 1307.510 52.870 ;
        RECT 1307.930 51.690 1309.110 52.870 ;
        RECT 1306.330 -22.110 1307.510 -20.930 ;
        RECT 1307.930 -22.110 1309.110 -20.930 ;
        RECT 1306.330 -23.710 1307.510 -22.530 ;
        RECT 1307.930 -23.710 1309.110 -22.530 ;
        RECT 1486.330 3542.210 1487.510 3543.390 ;
        RECT 1487.930 3542.210 1489.110 3543.390 ;
        RECT 1486.330 3540.610 1487.510 3541.790 ;
        RECT 1487.930 3540.610 1489.110 3541.790 ;
        RECT 1486.330 3473.290 1487.510 3474.470 ;
        RECT 1487.930 3473.290 1489.110 3474.470 ;
        RECT 1486.330 3471.690 1487.510 3472.870 ;
        RECT 1487.930 3471.690 1489.110 3472.870 ;
        RECT 1486.330 3293.290 1487.510 3294.470 ;
        RECT 1487.930 3293.290 1489.110 3294.470 ;
        RECT 1486.330 3291.690 1487.510 3292.870 ;
        RECT 1487.930 3291.690 1489.110 3292.870 ;
        RECT 1486.330 3113.290 1487.510 3114.470 ;
        RECT 1487.930 3113.290 1489.110 3114.470 ;
        RECT 1486.330 3111.690 1487.510 3112.870 ;
        RECT 1487.930 3111.690 1489.110 3112.870 ;
        RECT 1486.330 2933.290 1487.510 2934.470 ;
        RECT 1487.930 2933.290 1489.110 2934.470 ;
        RECT 1486.330 2931.690 1487.510 2932.870 ;
        RECT 1487.930 2931.690 1489.110 2932.870 ;
        RECT 1486.330 2753.290 1487.510 2754.470 ;
        RECT 1487.930 2753.290 1489.110 2754.470 ;
        RECT 1486.330 2751.690 1487.510 2752.870 ;
        RECT 1487.930 2751.690 1489.110 2752.870 ;
        RECT 1486.330 2573.290 1487.510 2574.470 ;
        RECT 1487.930 2573.290 1489.110 2574.470 ;
        RECT 1486.330 2571.690 1487.510 2572.870 ;
        RECT 1487.930 2571.690 1489.110 2572.870 ;
        RECT 1486.330 2393.290 1487.510 2394.470 ;
        RECT 1487.930 2393.290 1489.110 2394.470 ;
        RECT 1486.330 2391.690 1487.510 2392.870 ;
        RECT 1487.930 2391.690 1489.110 2392.870 ;
        RECT 1486.330 2213.290 1487.510 2214.470 ;
        RECT 1487.930 2213.290 1489.110 2214.470 ;
        RECT 1486.330 2211.690 1487.510 2212.870 ;
        RECT 1487.930 2211.690 1489.110 2212.870 ;
        RECT 1486.330 2033.290 1487.510 2034.470 ;
        RECT 1487.930 2033.290 1489.110 2034.470 ;
        RECT 1486.330 2031.690 1487.510 2032.870 ;
        RECT 1487.930 2031.690 1489.110 2032.870 ;
        RECT 1486.330 1853.290 1487.510 1854.470 ;
        RECT 1487.930 1853.290 1489.110 1854.470 ;
        RECT 1486.330 1851.690 1487.510 1852.870 ;
        RECT 1487.930 1851.690 1489.110 1852.870 ;
        RECT 1486.330 1673.290 1487.510 1674.470 ;
        RECT 1487.930 1673.290 1489.110 1674.470 ;
        RECT 1486.330 1671.690 1487.510 1672.870 ;
        RECT 1487.930 1671.690 1489.110 1672.870 ;
        RECT 1486.330 1493.290 1487.510 1494.470 ;
        RECT 1487.930 1493.290 1489.110 1494.470 ;
        RECT 1486.330 1491.690 1487.510 1492.870 ;
        RECT 1487.930 1491.690 1489.110 1492.870 ;
        RECT 1486.330 1313.290 1487.510 1314.470 ;
        RECT 1487.930 1313.290 1489.110 1314.470 ;
        RECT 1486.330 1311.690 1487.510 1312.870 ;
        RECT 1487.930 1311.690 1489.110 1312.870 ;
        RECT 1486.330 1133.290 1487.510 1134.470 ;
        RECT 1487.930 1133.290 1489.110 1134.470 ;
        RECT 1486.330 1131.690 1487.510 1132.870 ;
        RECT 1487.930 1131.690 1489.110 1132.870 ;
        RECT 1486.330 953.290 1487.510 954.470 ;
        RECT 1487.930 953.290 1489.110 954.470 ;
        RECT 1486.330 951.690 1487.510 952.870 ;
        RECT 1487.930 951.690 1489.110 952.870 ;
        RECT 1486.330 773.290 1487.510 774.470 ;
        RECT 1487.930 773.290 1489.110 774.470 ;
        RECT 1486.330 771.690 1487.510 772.870 ;
        RECT 1487.930 771.690 1489.110 772.870 ;
        RECT 1486.330 593.290 1487.510 594.470 ;
        RECT 1487.930 593.290 1489.110 594.470 ;
        RECT 1486.330 591.690 1487.510 592.870 ;
        RECT 1487.930 591.690 1489.110 592.870 ;
        RECT 1486.330 413.290 1487.510 414.470 ;
        RECT 1487.930 413.290 1489.110 414.470 ;
        RECT 1486.330 411.690 1487.510 412.870 ;
        RECT 1487.930 411.690 1489.110 412.870 ;
        RECT 1486.330 233.290 1487.510 234.470 ;
        RECT 1487.930 233.290 1489.110 234.470 ;
        RECT 1486.330 231.690 1487.510 232.870 ;
        RECT 1487.930 231.690 1489.110 232.870 ;
        RECT 1486.330 53.290 1487.510 54.470 ;
        RECT 1487.930 53.290 1489.110 54.470 ;
        RECT 1486.330 51.690 1487.510 52.870 ;
        RECT 1487.930 51.690 1489.110 52.870 ;
        RECT 1486.330 -22.110 1487.510 -20.930 ;
        RECT 1487.930 -22.110 1489.110 -20.930 ;
        RECT 1486.330 -23.710 1487.510 -22.530 ;
        RECT 1487.930 -23.710 1489.110 -22.530 ;
        RECT 1666.330 3542.210 1667.510 3543.390 ;
        RECT 1667.930 3542.210 1669.110 3543.390 ;
        RECT 1666.330 3540.610 1667.510 3541.790 ;
        RECT 1667.930 3540.610 1669.110 3541.790 ;
        RECT 1666.330 3473.290 1667.510 3474.470 ;
        RECT 1667.930 3473.290 1669.110 3474.470 ;
        RECT 1666.330 3471.690 1667.510 3472.870 ;
        RECT 1667.930 3471.690 1669.110 3472.870 ;
        RECT 1666.330 3293.290 1667.510 3294.470 ;
        RECT 1667.930 3293.290 1669.110 3294.470 ;
        RECT 1666.330 3291.690 1667.510 3292.870 ;
        RECT 1667.930 3291.690 1669.110 3292.870 ;
        RECT 1666.330 3113.290 1667.510 3114.470 ;
        RECT 1667.930 3113.290 1669.110 3114.470 ;
        RECT 1666.330 3111.690 1667.510 3112.870 ;
        RECT 1667.930 3111.690 1669.110 3112.870 ;
        RECT 1666.330 2933.290 1667.510 2934.470 ;
        RECT 1667.930 2933.290 1669.110 2934.470 ;
        RECT 1666.330 2931.690 1667.510 2932.870 ;
        RECT 1667.930 2931.690 1669.110 2932.870 ;
        RECT 1666.330 2753.290 1667.510 2754.470 ;
        RECT 1667.930 2753.290 1669.110 2754.470 ;
        RECT 1666.330 2751.690 1667.510 2752.870 ;
        RECT 1667.930 2751.690 1669.110 2752.870 ;
        RECT 1666.330 2573.290 1667.510 2574.470 ;
        RECT 1667.930 2573.290 1669.110 2574.470 ;
        RECT 1666.330 2571.690 1667.510 2572.870 ;
        RECT 1667.930 2571.690 1669.110 2572.870 ;
        RECT 1666.330 2393.290 1667.510 2394.470 ;
        RECT 1667.930 2393.290 1669.110 2394.470 ;
        RECT 1666.330 2391.690 1667.510 2392.870 ;
        RECT 1667.930 2391.690 1669.110 2392.870 ;
        RECT 1666.330 2213.290 1667.510 2214.470 ;
        RECT 1667.930 2213.290 1669.110 2214.470 ;
        RECT 1666.330 2211.690 1667.510 2212.870 ;
        RECT 1667.930 2211.690 1669.110 2212.870 ;
        RECT 1666.330 2033.290 1667.510 2034.470 ;
        RECT 1667.930 2033.290 1669.110 2034.470 ;
        RECT 1666.330 2031.690 1667.510 2032.870 ;
        RECT 1667.930 2031.690 1669.110 2032.870 ;
        RECT 1666.330 1853.290 1667.510 1854.470 ;
        RECT 1667.930 1853.290 1669.110 1854.470 ;
        RECT 1666.330 1851.690 1667.510 1852.870 ;
        RECT 1667.930 1851.690 1669.110 1852.870 ;
        RECT 1666.330 1673.290 1667.510 1674.470 ;
        RECT 1667.930 1673.290 1669.110 1674.470 ;
        RECT 1666.330 1671.690 1667.510 1672.870 ;
        RECT 1667.930 1671.690 1669.110 1672.870 ;
        RECT 1666.330 1493.290 1667.510 1494.470 ;
        RECT 1667.930 1493.290 1669.110 1494.470 ;
        RECT 1666.330 1491.690 1667.510 1492.870 ;
        RECT 1667.930 1491.690 1669.110 1492.870 ;
        RECT 1666.330 1313.290 1667.510 1314.470 ;
        RECT 1667.930 1313.290 1669.110 1314.470 ;
        RECT 1666.330 1311.690 1667.510 1312.870 ;
        RECT 1667.930 1311.690 1669.110 1312.870 ;
        RECT 1666.330 1133.290 1667.510 1134.470 ;
        RECT 1667.930 1133.290 1669.110 1134.470 ;
        RECT 1666.330 1131.690 1667.510 1132.870 ;
        RECT 1667.930 1131.690 1669.110 1132.870 ;
        RECT 1666.330 953.290 1667.510 954.470 ;
        RECT 1667.930 953.290 1669.110 954.470 ;
        RECT 1666.330 951.690 1667.510 952.870 ;
        RECT 1667.930 951.690 1669.110 952.870 ;
        RECT 1666.330 773.290 1667.510 774.470 ;
        RECT 1667.930 773.290 1669.110 774.470 ;
        RECT 1666.330 771.690 1667.510 772.870 ;
        RECT 1667.930 771.690 1669.110 772.870 ;
        RECT 1666.330 593.290 1667.510 594.470 ;
        RECT 1667.930 593.290 1669.110 594.470 ;
        RECT 1666.330 591.690 1667.510 592.870 ;
        RECT 1667.930 591.690 1669.110 592.870 ;
        RECT 1666.330 413.290 1667.510 414.470 ;
        RECT 1667.930 413.290 1669.110 414.470 ;
        RECT 1666.330 411.690 1667.510 412.870 ;
        RECT 1667.930 411.690 1669.110 412.870 ;
        RECT 1666.330 233.290 1667.510 234.470 ;
        RECT 1667.930 233.290 1669.110 234.470 ;
        RECT 1666.330 231.690 1667.510 232.870 ;
        RECT 1667.930 231.690 1669.110 232.870 ;
        RECT 1666.330 53.290 1667.510 54.470 ;
        RECT 1667.930 53.290 1669.110 54.470 ;
        RECT 1666.330 51.690 1667.510 52.870 ;
        RECT 1667.930 51.690 1669.110 52.870 ;
        RECT 1666.330 -22.110 1667.510 -20.930 ;
        RECT 1667.930 -22.110 1669.110 -20.930 ;
        RECT 1666.330 -23.710 1667.510 -22.530 ;
        RECT 1667.930 -23.710 1669.110 -22.530 ;
        RECT 1846.330 3542.210 1847.510 3543.390 ;
        RECT 1847.930 3542.210 1849.110 3543.390 ;
        RECT 1846.330 3540.610 1847.510 3541.790 ;
        RECT 1847.930 3540.610 1849.110 3541.790 ;
        RECT 1846.330 3473.290 1847.510 3474.470 ;
        RECT 1847.930 3473.290 1849.110 3474.470 ;
        RECT 1846.330 3471.690 1847.510 3472.870 ;
        RECT 1847.930 3471.690 1849.110 3472.870 ;
        RECT 1846.330 3293.290 1847.510 3294.470 ;
        RECT 1847.930 3293.290 1849.110 3294.470 ;
        RECT 1846.330 3291.690 1847.510 3292.870 ;
        RECT 1847.930 3291.690 1849.110 3292.870 ;
        RECT 1846.330 3113.290 1847.510 3114.470 ;
        RECT 1847.930 3113.290 1849.110 3114.470 ;
        RECT 1846.330 3111.690 1847.510 3112.870 ;
        RECT 1847.930 3111.690 1849.110 3112.870 ;
        RECT 1846.330 2933.290 1847.510 2934.470 ;
        RECT 1847.930 2933.290 1849.110 2934.470 ;
        RECT 1846.330 2931.690 1847.510 2932.870 ;
        RECT 1847.930 2931.690 1849.110 2932.870 ;
        RECT 1846.330 2753.290 1847.510 2754.470 ;
        RECT 1847.930 2753.290 1849.110 2754.470 ;
        RECT 1846.330 2751.690 1847.510 2752.870 ;
        RECT 1847.930 2751.690 1849.110 2752.870 ;
        RECT 1846.330 2573.290 1847.510 2574.470 ;
        RECT 1847.930 2573.290 1849.110 2574.470 ;
        RECT 1846.330 2571.690 1847.510 2572.870 ;
        RECT 1847.930 2571.690 1849.110 2572.870 ;
        RECT 1846.330 2393.290 1847.510 2394.470 ;
        RECT 1847.930 2393.290 1849.110 2394.470 ;
        RECT 1846.330 2391.690 1847.510 2392.870 ;
        RECT 1847.930 2391.690 1849.110 2392.870 ;
        RECT 1846.330 2213.290 1847.510 2214.470 ;
        RECT 1847.930 2213.290 1849.110 2214.470 ;
        RECT 1846.330 2211.690 1847.510 2212.870 ;
        RECT 1847.930 2211.690 1849.110 2212.870 ;
        RECT 1846.330 2033.290 1847.510 2034.470 ;
        RECT 1847.930 2033.290 1849.110 2034.470 ;
        RECT 1846.330 2031.690 1847.510 2032.870 ;
        RECT 1847.930 2031.690 1849.110 2032.870 ;
        RECT 1846.330 1853.290 1847.510 1854.470 ;
        RECT 1847.930 1853.290 1849.110 1854.470 ;
        RECT 1846.330 1851.690 1847.510 1852.870 ;
        RECT 1847.930 1851.690 1849.110 1852.870 ;
        RECT 1846.330 1673.290 1847.510 1674.470 ;
        RECT 1847.930 1673.290 1849.110 1674.470 ;
        RECT 1846.330 1671.690 1847.510 1672.870 ;
        RECT 1847.930 1671.690 1849.110 1672.870 ;
        RECT 1846.330 1493.290 1847.510 1494.470 ;
        RECT 1847.930 1493.290 1849.110 1494.470 ;
        RECT 1846.330 1491.690 1847.510 1492.870 ;
        RECT 1847.930 1491.690 1849.110 1492.870 ;
        RECT 1846.330 1313.290 1847.510 1314.470 ;
        RECT 1847.930 1313.290 1849.110 1314.470 ;
        RECT 1846.330 1311.690 1847.510 1312.870 ;
        RECT 1847.930 1311.690 1849.110 1312.870 ;
        RECT 1846.330 1133.290 1847.510 1134.470 ;
        RECT 1847.930 1133.290 1849.110 1134.470 ;
        RECT 1846.330 1131.690 1847.510 1132.870 ;
        RECT 1847.930 1131.690 1849.110 1132.870 ;
        RECT 1846.330 953.290 1847.510 954.470 ;
        RECT 1847.930 953.290 1849.110 954.470 ;
        RECT 1846.330 951.690 1847.510 952.870 ;
        RECT 1847.930 951.690 1849.110 952.870 ;
        RECT 1846.330 773.290 1847.510 774.470 ;
        RECT 1847.930 773.290 1849.110 774.470 ;
        RECT 1846.330 771.690 1847.510 772.870 ;
        RECT 1847.930 771.690 1849.110 772.870 ;
        RECT 1846.330 593.290 1847.510 594.470 ;
        RECT 1847.930 593.290 1849.110 594.470 ;
        RECT 1846.330 591.690 1847.510 592.870 ;
        RECT 1847.930 591.690 1849.110 592.870 ;
        RECT 1846.330 413.290 1847.510 414.470 ;
        RECT 1847.930 413.290 1849.110 414.470 ;
        RECT 1846.330 411.690 1847.510 412.870 ;
        RECT 1847.930 411.690 1849.110 412.870 ;
        RECT 1846.330 233.290 1847.510 234.470 ;
        RECT 1847.930 233.290 1849.110 234.470 ;
        RECT 1846.330 231.690 1847.510 232.870 ;
        RECT 1847.930 231.690 1849.110 232.870 ;
        RECT 1846.330 53.290 1847.510 54.470 ;
        RECT 1847.930 53.290 1849.110 54.470 ;
        RECT 1846.330 51.690 1847.510 52.870 ;
        RECT 1847.930 51.690 1849.110 52.870 ;
        RECT 1846.330 -22.110 1847.510 -20.930 ;
        RECT 1847.930 -22.110 1849.110 -20.930 ;
        RECT 1846.330 -23.710 1847.510 -22.530 ;
        RECT 1847.930 -23.710 1849.110 -22.530 ;
        RECT 2026.330 3542.210 2027.510 3543.390 ;
        RECT 2027.930 3542.210 2029.110 3543.390 ;
        RECT 2026.330 3540.610 2027.510 3541.790 ;
        RECT 2027.930 3540.610 2029.110 3541.790 ;
        RECT 2026.330 3473.290 2027.510 3474.470 ;
        RECT 2027.930 3473.290 2029.110 3474.470 ;
        RECT 2026.330 3471.690 2027.510 3472.870 ;
        RECT 2027.930 3471.690 2029.110 3472.870 ;
        RECT 2026.330 3293.290 2027.510 3294.470 ;
        RECT 2027.930 3293.290 2029.110 3294.470 ;
        RECT 2026.330 3291.690 2027.510 3292.870 ;
        RECT 2027.930 3291.690 2029.110 3292.870 ;
        RECT 2026.330 3113.290 2027.510 3114.470 ;
        RECT 2027.930 3113.290 2029.110 3114.470 ;
        RECT 2026.330 3111.690 2027.510 3112.870 ;
        RECT 2027.930 3111.690 2029.110 3112.870 ;
        RECT 2026.330 2933.290 2027.510 2934.470 ;
        RECT 2027.930 2933.290 2029.110 2934.470 ;
        RECT 2026.330 2931.690 2027.510 2932.870 ;
        RECT 2027.930 2931.690 2029.110 2932.870 ;
        RECT 2026.330 2753.290 2027.510 2754.470 ;
        RECT 2027.930 2753.290 2029.110 2754.470 ;
        RECT 2026.330 2751.690 2027.510 2752.870 ;
        RECT 2027.930 2751.690 2029.110 2752.870 ;
        RECT 2026.330 2573.290 2027.510 2574.470 ;
        RECT 2027.930 2573.290 2029.110 2574.470 ;
        RECT 2026.330 2571.690 2027.510 2572.870 ;
        RECT 2027.930 2571.690 2029.110 2572.870 ;
        RECT 2026.330 2393.290 2027.510 2394.470 ;
        RECT 2027.930 2393.290 2029.110 2394.470 ;
        RECT 2026.330 2391.690 2027.510 2392.870 ;
        RECT 2027.930 2391.690 2029.110 2392.870 ;
        RECT 2026.330 2213.290 2027.510 2214.470 ;
        RECT 2027.930 2213.290 2029.110 2214.470 ;
        RECT 2026.330 2211.690 2027.510 2212.870 ;
        RECT 2027.930 2211.690 2029.110 2212.870 ;
        RECT 2026.330 2033.290 2027.510 2034.470 ;
        RECT 2027.930 2033.290 2029.110 2034.470 ;
        RECT 2026.330 2031.690 2027.510 2032.870 ;
        RECT 2027.930 2031.690 2029.110 2032.870 ;
        RECT 2026.330 1853.290 2027.510 1854.470 ;
        RECT 2027.930 1853.290 2029.110 1854.470 ;
        RECT 2026.330 1851.690 2027.510 1852.870 ;
        RECT 2027.930 1851.690 2029.110 1852.870 ;
        RECT 2026.330 1673.290 2027.510 1674.470 ;
        RECT 2027.930 1673.290 2029.110 1674.470 ;
        RECT 2026.330 1671.690 2027.510 1672.870 ;
        RECT 2027.930 1671.690 2029.110 1672.870 ;
        RECT 2026.330 1493.290 2027.510 1494.470 ;
        RECT 2027.930 1493.290 2029.110 1494.470 ;
        RECT 2026.330 1491.690 2027.510 1492.870 ;
        RECT 2027.930 1491.690 2029.110 1492.870 ;
        RECT 2026.330 1313.290 2027.510 1314.470 ;
        RECT 2027.930 1313.290 2029.110 1314.470 ;
        RECT 2026.330 1311.690 2027.510 1312.870 ;
        RECT 2027.930 1311.690 2029.110 1312.870 ;
        RECT 2026.330 1133.290 2027.510 1134.470 ;
        RECT 2027.930 1133.290 2029.110 1134.470 ;
        RECT 2026.330 1131.690 2027.510 1132.870 ;
        RECT 2027.930 1131.690 2029.110 1132.870 ;
        RECT 2026.330 953.290 2027.510 954.470 ;
        RECT 2027.930 953.290 2029.110 954.470 ;
        RECT 2026.330 951.690 2027.510 952.870 ;
        RECT 2027.930 951.690 2029.110 952.870 ;
        RECT 2026.330 773.290 2027.510 774.470 ;
        RECT 2027.930 773.290 2029.110 774.470 ;
        RECT 2026.330 771.690 2027.510 772.870 ;
        RECT 2027.930 771.690 2029.110 772.870 ;
        RECT 2026.330 593.290 2027.510 594.470 ;
        RECT 2027.930 593.290 2029.110 594.470 ;
        RECT 2026.330 591.690 2027.510 592.870 ;
        RECT 2027.930 591.690 2029.110 592.870 ;
        RECT 2026.330 413.290 2027.510 414.470 ;
        RECT 2027.930 413.290 2029.110 414.470 ;
        RECT 2026.330 411.690 2027.510 412.870 ;
        RECT 2027.930 411.690 2029.110 412.870 ;
        RECT 2026.330 233.290 2027.510 234.470 ;
        RECT 2027.930 233.290 2029.110 234.470 ;
        RECT 2026.330 231.690 2027.510 232.870 ;
        RECT 2027.930 231.690 2029.110 232.870 ;
        RECT 2026.330 53.290 2027.510 54.470 ;
        RECT 2027.930 53.290 2029.110 54.470 ;
        RECT 2026.330 51.690 2027.510 52.870 ;
        RECT 2027.930 51.690 2029.110 52.870 ;
        RECT 2026.330 -22.110 2027.510 -20.930 ;
        RECT 2027.930 -22.110 2029.110 -20.930 ;
        RECT 2026.330 -23.710 2027.510 -22.530 ;
        RECT 2027.930 -23.710 2029.110 -22.530 ;
        RECT 2206.330 3542.210 2207.510 3543.390 ;
        RECT 2207.930 3542.210 2209.110 3543.390 ;
        RECT 2206.330 3540.610 2207.510 3541.790 ;
        RECT 2207.930 3540.610 2209.110 3541.790 ;
        RECT 2206.330 3473.290 2207.510 3474.470 ;
        RECT 2207.930 3473.290 2209.110 3474.470 ;
        RECT 2206.330 3471.690 2207.510 3472.870 ;
        RECT 2207.930 3471.690 2209.110 3472.870 ;
        RECT 2206.330 3293.290 2207.510 3294.470 ;
        RECT 2207.930 3293.290 2209.110 3294.470 ;
        RECT 2206.330 3291.690 2207.510 3292.870 ;
        RECT 2207.930 3291.690 2209.110 3292.870 ;
        RECT 2206.330 3113.290 2207.510 3114.470 ;
        RECT 2207.930 3113.290 2209.110 3114.470 ;
        RECT 2206.330 3111.690 2207.510 3112.870 ;
        RECT 2207.930 3111.690 2209.110 3112.870 ;
        RECT 2206.330 2933.290 2207.510 2934.470 ;
        RECT 2207.930 2933.290 2209.110 2934.470 ;
        RECT 2206.330 2931.690 2207.510 2932.870 ;
        RECT 2207.930 2931.690 2209.110 2932.870 ;
        RECT 2206.330 2753.290 2207.510 2754.470 ;
        RECT 2207.930 2753.290 2209.110 2754.470 ;
        RECT 2206.330 2751.690 2207.510 2752.870 ;
        RECT 2207.930 2751.690 2209.110 2752.870 ;
        RECT 2206.330 2573.290 2207.510 2574.470 ;
        RECT 2207.930 2573.290 2209.110 2574.470 ;
        RECT 2206.330 2571.690 2207.510 2572.870 ;
        RECT 2207.930 2571.690 2209.110 2572.870 ;
        RECT 2206.330 2393.290 2207.510 2394.470 ;
        RECT 2207.930 2393.290 2209.110 2394.470 ;
        RECT 2206.330 2391.690 2207.510 2392.870 ;
        RECT 2207.930 2391.690 2209.110 2392.870 ;
        RECT 2206.330 2213.290 2207.510 2214.470 ;
        RECT 2207.930 2213.290 2209.110 2214.470 ;
        RECT 2206.330 2211.690 2207.510 2212.870 ;
        RECT 2207.930 2211.690 2209.110 2212.870 ;
        RECT 2206.330 2033.290 2207.510 2034.470 ;
        RECT 2207.930 2033.290 2209.110 2034.470 ;
        RECT 2206.330 2031.690 2207.510 2032.870 ;
        RECT 2207.930 2031.690 2209.110 2032.870 ;
        RECT 2206.330 1853.290 2207.510 1854.470 ;
        RECT 2207.930 1853.290 2209.110 1854.470 ;
        RECT 2206.330 1851.690 2207.510 1852.870 ;
        RECT 2207.930 1851.690 2209.110 1852.870 ;
        RECT 2206.330 1673.290 2207.510 1674.470 ;
        RECT 2207.930 1673.290 2209.110 1674.470 ;
        RECT 2206.330 1671.690 2207.510 1672.870 ;
        RECT 2207.930 1671.690 2209.110 1672.870 ;
        RECT 2206.330 1493.290 2207.510 1494.470 ;
        RECT 2207.930 1493.290 2209.110 1494.470 ;
        RECT 2206.330 1491.690 2207.510 1492.870 ;
        RECT 2207.930 1491.690 2209.110 1492.870 ;
        RECT 2206.330 1313.290 2207.510 1314.470 ;
        RECT 2207.930 1313.290 2209.110 1314.470 ;
        RECT 2206.330 1311.690 2207.510 1312.870 ;
        RECT 2207.930 1311.690 2209.110 1312.870 ;
        RECT 2206.330 1133.290 2207.510 1134.470 ;
        RECT 2207.930 1133.290 2209.110 1134.470 ;
        RECT 2206.330 1131.690 2207.510 1132.870 ;
        RECT 2207.930 1131.690 2209.110 1132.870 ;
        RECT 2206.330 953.290 2207.510 954.470 ;
        RECT 2207.930 953.290 2209.110 954.470 ;
        RECT 2206.330 951.690 2207.510 952.870 ;
        RECT 2207.930 951.690 2209.110 952.870 ;
        RECT 2206.330 773.290 2207.510 774.470 ;
        RECT 2207.930 773.290 2209.110 774.470 ;
        RECT 2206.330 771.690 2207.510 772.870 ;
        RECT 2207.930 771.690 2209.110 772.870 ;
        RECT 2206.330 593.290 2207.510 594.470 ;
        RECT 2207.930 593.290 2209.110 594.470 ;
        RECT 2206.330 591.690 2207.510 592.870 ;
        RECT 2207.930 591.690 2209.110 592.870 ;
        RECT 2206.330 413.290 2207.510 414.470 ;
        RECT 2207.930 413.290 2209.110 414.470 ;
        RECT 2206.330 411.690 2207.510 412.870 ;
        RECT 2207.930 411.690 2209.110 412.870 ;
        RECT 2206.330 233.290 2207.510 234.470 ;
        RECT 2207.930 233.290 2209.110 234.470 ;
        RECT 2206.330 231.690 2207.510 232.870 ;
        RECT 2207.930 231.690 2209.110 232.870 ;
        RECT 2206.330 53.290 2207.510 54.470 ;
        RECT 2207.930 53.290 2209.110 54.470 ;
        RECT 2206.330 51.690 2207.510 52.870 ;
        RECT 2207.930 51.690 2209.110 52.870 ;
        RECT 2206.330 -22.110 2207.510 -20.930 ;
        RECT 2207.930 -22.110 2209.110 -20.930 ;
        RECT 2206.330 -23.710 2207.510 -22.530 ;
        RECT 2207.930 -23.710 2209.110 -22.530 ;
        RECT 2386.330 3542.210 2387.510 3543.390 ;
        RECT 2387.930 3542.210 2389.110 3543.390 ;
        RECT 2386.330 3540.610 2387.510 3541.790 ;
        RECT 2387.930 3540.610 2389.110 3541.790 ;
        RECT 2386.330 3473.290 2387.510 3474.470 ;
        RECT 2387.930 3473.290 2389.110 3474.470 ;
        RECT 2386.330 3471.690 2387.510 3472.870 ;
        RECT 2387.930 3471.690 2389.110 3472.870 ;
        RECT 2386.330 3293.290 2387.510 3294.470 ;
        RECT 2387.930 3293.290 2389.110 3294.470 ;
        RECT 2386.330 3291.690 2387.510 3292.870 ;
        RECT 2387.930 3291.690 2389.110 3292.870 ;
        RECT 2386.330 3113.290 2387.510 3114.470 ;
        RECT 2387.930 3113.290 2389.110 3114.470 ;
        RECT 2386.330 3111.690 2387.510 3112.870 ;
        RECT 2387.930 3111.690 2389.110 3112.870 ;
        RECT 2386.330 2933.290 2387.510 2934.470 ;
        RECT 2387.930 2933.290 2389.110 2934.470 ;
        RECT 2386.330 2931.690 2387.510 2932.870 ;
        RECT 2387.930 2931.690 2389.110 2932.870 ;
        RECT 2386.330 2753.290 2387.510 2754.470 ;
        RECT 2387.930 2753.290 2389.110 2754.470 ;
        RECT 2386.330 2751.690 2387.510 2752.870 ;
        RECT 2387.930 2751.690 2389.110 2752.870 ;
        RECT 2386.330 2573.290 2387.510 2574.470 ;
        RECT 2387.930 2573.290 2389.110 2574.470 ;
        RECT 2386.330 2571.690 2387.510 2572.870 ;
        RECT 2387.930 2571.690 2389.110 2572.870 ;
        RECT 2386.330 2393.290 2387.510 2394.470 ;
        RECT 2387.930 2393.290 2389.110 2394.470 ;
        RECT 2386.330 2391.690 2387.510 2392.870 ;
        RECT 2387.930 2391.690 2389.110 2392.870 ;
        RECT 2386.330 2213.290 2387.510 2214.470 ;
        RECT 2387.930 2213.290 2389.110 2214.470 ;
        RECT 2386.330 2211.690 2387.510 2212.870 ;
        RECT 2387.930 2211.690 2389.110 2212.870 ;
        RECT 2386.330 2033.290 2387.510 2034.470 ;
        RECT 2387.930 2033.290 2389.110 2034.470 ;
        RECT 2386.330 2031.690 2387.510 2032.870 ;
        RECT 2387.930 2031.690 2389.110 2032.870 ;
        RECT 2386.330 1853.290 2387.510 1854.470 ;
        RECT 2387.930 1853.290 2389.110 1854.470 ;
        RECT 2386.330 1851.690 2387.510 1852.870 ;
        RECT 2387.930 1851.690 2389.110 1852.870 ;
        RECT 2386.330 1673.290 2387.510 1674.470 ;
        RECT 2387.930 1673.290 2389.110 1674.470 ;
        RECT 2386.330 1671.690 2387.510 1672.870 ;
        RECT 2387.930 1671.690 2389.110 1672.870 ;
        RECT 2386.330 1493.290 2387.510 1494.470 ;
        RECT 2387.930 1493.290 2389.110 1494.470 ;
        RECT 2386.330 1491.690 2387.510 1492.870 ;
        RECT 2387.930 1491.690 2389.110 1492.870 ;
        RECT 2386.330 1313.290 2387.510 1314.470 ;
        RECT 2387.930 1313.290 2389.110 1314.470 ;
        RECT 2386.330 1311.690 2387.510 1312.870 ;
        RECT 2387.930 1311.690 2389.110 1312.870 ;
        RECT 2386.330 1133.290 2387.510 1134.470 ;
        RECT 2387.930 1133.290 2389.110 1134.470 ;
        RECT 2386.330 1131.690 2387.510 1132.870 ;
        RECT 2387.930 1131.690 2389.110 1132.870 ;
        RECT 2386.330 953.290 2387.510 954.470 ;
        RECT 2387.930 953.290 2389.110 954.470 ;
        RECT 2386.330 951.690 2387.510 952.870 ;
        RECT 2387.930 951.690 2389.110 952.870 ;
        RECT 2386.330 773.290 2387.510 774.470 ;
        RECT 2387.930 773.290 2389.110 774.470 ;
        RECT 2386.330 771.690 2387.510 772.870 ;
        RECT 2387.930 771.690 2389.110 772.870 ;
        RECT 2386.330 593.290 2387.510 594.470 ;
        RECT 2387.930 593.290 2389.110 594.470 ;
        RECT 2386.330 591.690 2387.510 592.870 ;
        RECT 2387.930 591.690 2389.110 592.870 ;
        RECT 2386.330 413.290 2387.510 414.470 ;
        RECT 2387.930 413.290 2389.110 414.470 ;
        RECT 2386.330 411.690 2387.510 412.870 ;
        RECT 2387.930 411.690 2389.110 412.870 ;
        RECT 2386.330 233.290 2387.510 234.470 ;
        RECT 2387.930 233.290 2389.110 234.470 ;
        RECT 2386.330 231.690 2387.510 232.870 ;
        RECT 2387.930 231.690 2389.110 232.870 ;
        RECT 2386.330 53.290 2387.510 54.470 ;
        RECT 2387.930 53.290 2389.110 54.470 ;
        RECT 2386.330 51.690 2387.510 52.870 ;
        RECT 2387.930 51.690 2389.110 52.870 ;
        RECT 2386.330 -22.110 2387.510 -20.930 ;
        RECT 2387.930 -22.110 2389.110 -20.930 ;
        RECT 2386.330 -23.710 2387.510 -22.530 ;
        RECT 2387.930 -23.710 2389.110 -22.530 ;
        RECT 2566.330 3542.210 2567.510 3543.390 ;
        RECT 2567.930 3542.210 2569.110 3543.390 ;
        RECT 2566.330 3540.610 2567.510 3541.790 ;
        RECT 2567.930 3540.610 2569.110 3541.790 ;
        RECT 2566.330 3473.290 2567.510 3474.470 ;
        RECT 2567.930 3473.290 2569.110 3474.470 ;
        RECT 2566.330 3471.690 2567.510 3472.870 ;
        RECT 2567.930 3471.690 2569.110 3472.870 ;
        RECT 2566.330 3293.290 2567.510 3294.470 ;
        RECT 2567.930 3293.290 2569.110 3294.470 ;
        RECT 2566.330 3291.690 2567.510 3292.870 ;
        RECT 2567.930 3291.690 2569.110 3292.870 ;
        RECT 2566.330 3113.290 2567.510 3114.470 ;
        RECT 2567.930 3113.290 2569.110 3114.470 ;
        RECT 2566.330 3111.690 2567.510 3112.870 ;
        RECT 2567.930 3111.690 2569.110 3112.870 ;
        RECT 2566.330 2933.290 2567.510 2934.470 ;
        RECT 2567.930 2933.290 2569.110 2934.470 ;
        RECT 2566.330 2931.690 2567.510 2932.870 ;
        RECT 2567.930 2931.690 2569.110 2932.870 ;
        RECT 2566.330 2753.290 2567.510 2754.470 ;
        RECT 2567.930 2753.290 2569.110 2754.470 ;
        RECT 2566.330 2751.690 2567.510 2752.870 ;
        RECT 2567.930 2751.690 2569.110 2752.870 ;
        RECT 2566.330 2573.290 2567.510 2574.470 ;
        RECT 2567.930 2573.290 2569.110 2574.470 ;
        RECT 2566.330 2571.690 2567.510 2572.870 ;
        RECT 2567.930 2571.690 2569.110 2572.870 ;
        RECT 2566.330 2393.290 2567.510 2394.470 ;
        RECT 2567.930 2393.290 2569.110 2394.470 ;
        RECT 2566.330 2391.690 2567.510 2392.870 ;
        RECT 2567.930 2391.690 2569.110 2392.870 ;
        RECT 2566.330 2213.290 2567.510 2214.470 ;
        RECT 2567.930 2213.290 2569.110 2214.470 ;
        RECT 2566.330 2211.690 2567.510 2212.870 ;
        RECT 2567.930 2211.690 2569.110 2212.870 ;
        RECT 2566.330 2033.290 2567.510 2034.470 ;
        RECT 2567.930 2033.290 2569.110 2034.470 ;
        RECT 2566.330 2031.690 2567.510 2032.870 ;
        RECT 2567.930 2031.690 2569.110 2032.870 ;
        RECT 2566.330 1853.290 2567.510 1854.470 ;
        RECT 2567.930 1853.290 2569.110 1854.470 ;
        RECT 2566.330 1851.690 2567.510 1852.870 ;
        RECT 2567.930 1851.690 2569.110 1852.870 ;
        RECT 2566.330 1673.290 2567.510 1674.470 ;
        RECT 2567.930 1673.290 2569.110 1674.470 ;
        RECT 2566.330 1671.690 2567.510 1672.870 ;
        RECT 2567.930 1671.690 2569.110 1672.870 ;
        RECT 2566.330 1493.290 2567.510 1494.470 ;
        RECT 2567.930 1493.290 2569.110 1494.470 ;
        RECT 2566.330 1491.690 2567.510 1492.870 ;
        RECT 2567.930 1491.690 2569.110 1492.870 ;
        RECT 2566.330 1313.290 2567.510 1314.470 ;
        RECT 2567.930 1313.290 2569.110 1314.470 ;
        RECT 2566.330 1311.690 2567.510 1312.870 ;
        RECT 2567.930 1311.690 2569.110 1312.870 ;
        RECT 2566.330 1133.290 2567.510 1134.470 ;
        RECT 2567.930 1133.290 2569.110 1134.470 ;
        RECT 2566.330 1131.690 2567.510 1132.870 ;
        RECT 2567.930 1131.690 2569.110 1132.870 ;
        RECT 2566.330 953.290 2567.510 954.470 ;
        RECT 2567.930 953.290 2569.110 954.470 ;
        RECT 2566.330 951.690 2567.510 952.870 ;
        RECT 2567.930 951.690 2569.110 952.870 ;
        RECT 2566.330 773.290 2567.510 774.470 ;
        RECT 2567.930 773.290 2569.110 774.470 ;
        RECT 2566.330 771.690 2567.510 772.870 ;
        RECT 2567.930 771.690 2569.110 772.870 ;
        RECT 2566.330 593.290 2567.510 594.470 ;
        RECT 2567.930 593.290 2569.110 594.470 ;
        RECT 2566.330 591.690 2567.510 592.870 ;
        RECT 2567.930 591.690 2569.110 592.870 ;
        RECT 2566.330 413.290 2567.510 414.470 ;
        RECT 2567.930 413.290 2569.110 414.470 ;
        RECT 2566.330 411.690 2567.510 412.870 ;
        RECT 2567.930 411.690 2569.110 412.870 ;
        RECT 2566.330 233.290 2567.510 234.470 ;
        RECT 2567.930 233.290 2569.110 234.470 ;
        RECT 2566.330 231.690 2567.510 232.870 ;
        RECT 2567.930 231.690 2569.110 232.870 ;
        RECT 2566.330 53.290 2567.510 54.470 ;
        RECT 2567.930 53.290 2569.110 54.470 ;
        RECT 2566.330 51.690 2567.510 52.870 ;
        RECT 2567.930 51.690 2569.110 52.870 ;
        RECT 2566.330 -22.110 2567.510 -20.930 ;
        RECT 2567.930 -22.110 2569.110 -20.930 ;
        RECT 2566.330 -23.710 2567.510 -22.530 ;
        RECT 2567.930 -23.710 2569.110 -22.530 ;
        RECT 2746.330 3542.210 2747.510 3543.390 ;
        RECT 2747.930 3542.210 2749.110 3543.390 ;
        RECT 2746.330 3540.610 2747.510 3541.790 ;
        RECT 2747.930 3540.610 2749.110 3541.790 ;
        RECT 2746.330 3473.290 2747.510 3474.470 ;
        RECT 2747.930 3473.290 2749.110 3474.470 ;
        RECT 2746.330 3471.690 2747.510 3472.870 ;
        RECT 2747.930 3471.690 2749.110 3472.870 ;
        RECT 2746.330 3293.290 2747.510 3294.470 ;
        RECT 2747.930 3293.290 2749.110 3294.470 ;
        RECT 2746.330 3291.690 2747.510 3292.870 ;
        RECT 2747.930 3291.690 2749.110 3292.870 ;
        RECT 2746.330 3113.290 2747.510 3114.470 ;
        RECT 2747.930 3113.290 2749.110 3114.470 ;
        RECT 2746.330 3111.690 2747.510 3112.870 ;
        RECT 2747.930 3111.690 2749.110 3112.870 ;
        RECT 2746.330 2933.290 2747.510 2934.470 ;
        RECT 2747.930 2933.290 2749.110 2934.470 ;
        RECT 2746.330 2931.690 2747.510 2932.870 ;
        RECT 2747.930 2931.690 2749.110 2932.870 ;
        RECT 2746.330 2753.290 2747.510 2754.470 ;
        RECT 2747.930 2753.290 2749.110 2754.470 ;
        RECT 2746.330 2751.690 2747.510 2752.870 ;
        RECT 2747.930 2751.690 2749.110 2752.870 ;
        RECT 2746.330 2573.290 2747.510 2574.470 ;
        RECT 2747.930 2573.290 2749.110 2574.470 ;
        RECT 2746.330 2571.690 2747.510 2572.870 ;
        RECT 2747.930 2571.690 2749.110 2572.870 ;
        RECT 2746.330 2393.290 2747.510 2394.470 ;
        RECT 2747.930 2393.290 2749.110 2394.470 ;
        RECT 2746.330 2391.690 2747.510 2392.870 ;
        RECT 2747.930 2391.690 2749.110 2392.870 ;
        RECT 2746.330 2213.290 2747.510 2214.470 ;
        RECT 2747.930 2213.290 2749.110 2214.470 ;
        RECT 2746.330 2211.690 2747.510 2212.870 ;
        RECT 2747.930 2211.690 2749.110 2212.870 ;
        RECT 2746.330 2033.290 2747.510 2034.470 ;
        RECT 2747.930 2033.290 2749.110 2034.470 ;
        RECT 2746.330 2031.690 2747.510 2032.870 ;
        RECT 2747.930 2031.690 2749.110 2032.870 ;
        RECT 2746.330 1853.290 2747.510 1854.470 ;
        RECT 2747.930 1853.290 2749.110 1854.470 ;
        RECT 2746.330 1851.690 2747.510 1852.870 ;
        RECT 2747.930 1851.690 2749.110 1852.870 ;
        RECT 2746.330 1673.290 2747.510 1674.470 ;
        RECT 2747.930 1673.290 2749.110 1674.470 ;
        RECT 2746.330 1671.690 2747.510 1672.870 ;
        RECT 2747.930 1671.690 2749.110 1672.870 ;
        RECT 2746.330 1493.290 2747.510 1494.470 ;
        RECT 2747.930 1493.290 2749.110 1494.470 ;
        RECT 2746.330 1491.690 2747.510 1492.870 ;
        RECT 2747.930 1491.690 2749.110 1492.870 ;
        RECT 2746.330 1313.290 2747.510 1314.470 ;
        RECT 2747.930 1313.290 2749.110 1314.470 ;
        RECT 2746.330 1311.690 2747.510 1312.870 ;
        RECT 2747.930 1311.690 2749.110 1312.870 ;
        RECT 2746.330 1133.290 2747.510 1134.470 ;
        RECT 2747.930 1133.290 2749.110 1134.470 ;
        RECT 2746.330 1131.690 2747.510 1132.870 ;
        RECT 2747.930 1131.690 2749.110 1132.870 ;
        RECT 2746.330 953.290 2747.510 954.470 ;
        RECT 2747.930 953.290 2749.110 954.470 ;
        RECT 2746.330 951.690 2747.510 952.870 ;
        RECT 2747.930 951.690 2749.110 952.870 ;
        RECT 2746.330 773.290 2747.510 774.470 ;
        RECT 2747.930 773.290 2749.110 774.470 ;
        RECT 2746.330 771.690 2747.510 772.870 ;
        RECT 2747.930 771.690 2749.110 772.870 ;
        RECT 2746.330 593.290 2747.510 594.470 ;
        RECT 2747.930 593.290 2749.110 594.470 ;
        RECT 2746.330 591.690 2747.510 592.870 ;
        RECT 2747.930 591.690 2749.110 592.870 ;
        RECT 2746.330 413.290 2747.510 414.470 ;
        RECT 2747.930 413.290 2749.110 414.470 ;
        RECT 2746.330 411.690 2747.510 412.870 ;
        RECT 2747.930 411.690 2749.110 412.870 ;
        RECT 2746.330 233.290 2747.510 234.470 ;
        RECT 2747.930 233.290 2749.110 234.470 ;
        RECT 2746.330 231.690 2747.510 232.870 ;
        RECT 2747.930 231.690 2749.110 232.870 ;
        RECT 2746.330 53.290 2747.510 54.470 ;
        RECT 2747.930 53.290 2749.110 54.470 ;
        RECT 2746.330 51.690 2747.510 52.870 ;
        RECT 2747.930 51.690 2749.110 52.870 ;
        RECT 2746.330 -22.110 2747.510 -20.930 ;
        RECT 2747.930 -22.110 2749.110 -20.930 ;
        RECT 2746.330 -23.710 2747.510 -22.530 ;
        RECT 2747.930 -23.710 2749.110 -22.530 ;
        RECT 2945.910 3542.210 2947.090 3543.390 ;
        RECT 2947.510 3542.210 2948.690 3543.390 ;
        RECT 2945.910 3540.610 2947.090 3541.790 ;
        RECT 2947.510 3540.610 2948.690 3541.790 ;
        RECT 2945.910 3473.290 2947.090 3474.470 ;
        RECT 2947.510 3473.290 2948.690 3474.470 ;
        RECT 2945.910 3471.690 2947.090 3472.870 ;
        RECT 2947.510 3471.690 2948.690 3472.870 ;
        RECT 2945.910 3293.290 2947.090 3294.470 ;
        RECT 2947.510 3293.290 2948.690 3294.470 ;
        RECT 2945.910 3291.690 2947.090 3292.870 ;
        RECT 2947.510 3291.690 2948.690 3292.870 ;
        RECT 2945.910 3113.290 2947.090 3114.470 ;
        RECT 2947.510 3113.290 2948.690 3114.470 ;
        RECT 2945.910 3111.690 2947.090 3112.870 ;
        RECT 2947.510 3111.690 2948.690 3112.870 ;
        RECT 2945.910 2933.290 2947.090 2934.470 ;
        RECT 2947.510 2933.290 2948.690 2934.470 ;
        RECT 2945.910 2931.690 2947.090 2932.870 ;
        RECT 2947.510 2931.690 2948.690 2932.870 ;
        RECT 2945.910 2753.290 2947.090 2754.470 ;
        RECT 2947.510 2753.290 2948.690 2754.470 ;
        RECT 2945.910 2751.690 2947.090 2752.870 ;
        RECT 2947.510 2751.690 2948.690 2752.870 ;
        RECT 2945.910 2573.290 2947.090 2574.470 ;
        RECT 2947.510 2573.290 2948.690 2574.470 ;
        RECT 2945.910 2571.690 2947.090 2572.870 ;
        RECT 2947.510 2571.690 2948.690 2572.870 ;
        RECT 2945.910 2393.290 2947.090 2394.470 ;
        RECT 2947.510 2393.290 2948.690 2394.470 ;
        RECT 2945.910 2391.690 2947.090 2392.870 ;
        RECT 2947.510 2391.690 2948.690 2392.870 ;
        RECT 2945.910 2213.290 2947.090 2214.470 ;
        RECT 2947.510 2213.290 2948.690 2214.470 ;
        RECT 2945.910 2211.690 2947.090 2212.870 ;
        RECT 2947.510 2211.690 2948.690 2212.870 ;
        RECT 2945.910 2033.290 2947.090 2034.470 ;
        RECT 2947.510 2033.290 2948.690 2034.470 ;
        RECT 2945.910 2031.690 2947.090 2032.870 ;
        RECT 2947.510 2031.690 2948.690 2032.870 ;
        RECT 2945.910 1853.290 2947.090 1854.470 ;
        RECT 2947.510 1853.290 2948.690 1854.470 ;
        RECT 2945.910 1851.690 2947.090 1852.870 ;
        RECT 2947.510 1851.690 2948.690 1852.870 ;
        RECT 2945.910 1673.290 2947.090 1674.470 ;
        RECT 2947.510 1673.290 2948.690 1674.470 ;
        RECT 2945.910 1671.690 2947.090 1672.870 ;
        RECT 2947.510 1671.690 2948.690 1672.870 ;
        RECT 2945.910 1493.290 2947.090 1494.470 ;
        RECT 2947.510 1493.290 2948.690 1494.470 ;
        RECT 2945.910 1491.690 2947.090 1492.870 ;
        RECT 2947.510 1491.690 2948.690 1492.870 ;
        RECT 2945.910 1313.290 2947.090 1314.470 ;
        RECT 2947.510 1313.290 2948.690 1314.470 ;
        RECT 2945.910 1311.690 2947.090 1312.870 ;
        RECT 2947.510 1311.690 2948.690 1312.870 ;
        RECT 2945.910 1133.290 2947.090 1134.470 ;
        RECT 2947.510 1133.290 2948.690 1134.470 ;
        RECT 2945.910 1131.690 2947.090 1132.870 ;
        RECT 2947.510 1131.690 2948.690 1132.870 ;
        RECT 2945.910 953.290 2947.090 954.470 ;
        RECT 2947.510 953.290 2948.690 954.470 ;
        RECT 2945.910 951.690 2947.090 952.870 ;
        RECT 2947.510 951.690 2948.690 952.870 ;
        RECT 2945.910 773.290 2947.090 774.470 ;
        RECT 2947.510 773.290 2948.690 774.470 ;
        RECT 2945.910 771.690 2947.090 772.870 ;
        RECT 2947.510 771.690 2948.690 772.870 ;
        RECT 2945.910 593.290 2947.090 594.470 ;
        RECT 2947.510 593.290 2948.690 594.470 ;
        RECT 2945.910 591.690 2947.090 592.870 ;
        RECT 2947.510 591.690 2948.690 592.870 ;
        RECT 2945.910 413.290 2947.090 414.470 ;
        RECT 2947.510 413.290 2948.690 414.470 ;
        RECT 2945.910 411.690 2947.090 412.870 ;
        RECT 2947.510 411.690 2948.690 412.870 ;
        RECT 2945.910 233.290 2947.090 234.470 ;
        RECT 2947.510 233.290 2948.690 234.470 ;
        RECT 2945.910 231.690 2947.090 232.870 ;
        RECT 2947.510 231.690 2948.690 232.870 ;
        RECT 2945.910 53.290 2947.090 54.470 ;
        RECT 2947.510 53.290 2948.690 54.470 ;
        RECT 2945.910 51.690 2947.090 52.870 ;
        RECT 2947.510 51.690 2948.690 52.870 ;
        RECT 2945.910 -22.110 2947.090 -20.930 ;
        RECT 2947.510 -22.110 2948.690 -20.930 ;
        RECT 2945.910 -23.710 2947.090 -22.530 ;
        RECT 2947.510 -23.710 2948.690 -22.530 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
        RECT -34.030 951.530 2953.650 954.630 ;
        RECT -34.030 771.530 2953.650 774.630 ;
        RECT -34.030 591.530 2953.650 594.630 ;
        RECT -34.030 411.530 2953.650 414.630 ;
        RECT -34.030 231.530 2953.650 234.630 ;
        RECT -34.030 51.530 2953.650 54.630 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
        RECT 244.770 1010.000 247.870 3557.950 ;
        RECT 424.770 1010.000 427.870 3557.950 ;
        RECT 604.770 1010.000 607.870 3557.950 ;
        RECT 784.770 1010.000 787.870 3557.950 ;
        RECT 964.770 1010.000 967.870 3557.950 ;
        RECT 244.770 -38.270 247.870 390.000 ;
        RECT 424.770 -38.270 427.870 390.000 ;
        RECT 604.770 -38.270 607.870 390.000 ;
        RECT 784.770 -38.270 787.870 390.000 ;
        RECT 964.770 -38.270 967.870 390.000 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER via4 ;
        RECT -38.670 3551.810 -37.490 3552.990 ;
        RECT -37.070 3551.810 -35.890 3552.990 ;
        RECT -38.670 3550.210 -37.490 3551.390 ;
        RECT -37.070 3550.210 -35.890 3551.390 ;
        RECT -38.670 3491.890 -37.490 3493.070 ;
        RECT -37.070 3491.890 -35.890 3493.070 ;
        RECT -38.670 3490.290 -37.490 3491.470 ;
        RECT -37.070 3490.290 -35.890 3491.470 ;
        RECT -38.670 3311.890 -37.490 3313.070 ;
        RECT -37.070 3311.890 -35.890 3313.070 ;
        RECT -38.670 3310.290 -37.490 3311.470 ;
        RECT -37.070 3310.290 -35.890 3311.470 ;
        RECT -38.670 3131.890 -37.490 3133.070 ;
        RECT -37.070 3131.890 -35.890 3133.070 ;
        RECT -38.670 3130.290 -37.490 3131.470 ;
        RECT -37.070 3130.290 -35.890 3131.470 ;
        RECT -38.670 2951.890 -37.490 2953.070 ;
        RECT -37.070 2951.890 -35.890 2953.070 ;
        RECT -38.670 2950.290 -37.490 2951.470 ;
        RECT -37.070 2950.290 -35.890 2951.470 ;
        RECT -38.670 2771.890 -37.490 2773.070 ;
        RECT -37.070 2771.890 -35.890 2773.070 ;
        RECT -38.670 2770.290 -37.490 2771.470 ;
        RECT -37.070 2770.290 -35.890 2771.470 ;
        RECT -38.670 2591.890 -37.490 2593.070 ;
        RECT -37.070 2591.890 -35.890 2593.070 ;
        RECT -38.670 2590.290 -37.490 2591.470 ;
        RECT -37.070 2590.290 -35.890 2591.470 ;
        RECT -38.670 2411.890 -37.490 2413.070 ;
        RECT -37.070 2411.890 -35.890 2413.070 ;
        RECT -38.670 2410.290 -37.490 2411.470 ;
        RECT -37.070 2410.290 -35.890 2411.470 ;
        RECT -38.670 2231.890 -37.490 2233.070 ;
        RECT -37.070 2231.890 -35.890 2233.070 ;
        RECT -38.670 2230.290 -37.490 2231.470 ;
        RECT -37.070 2230.290 -35.890 2231.470 ;
        RECT -38.670 2051.890 -37.490 2053.070 ;
        RECT -37.070 2051.890 -35.890 2053.070 ;
        RECT -38.670 2050.290 -37.490 2051.470 ;
        RECT -37.070 2050.290 -35.890 2051.470 ;
        RECT -38.670 1871.890 -37.490 1873.070 ;
        RECT -37.070 1871.890 -35.890 1873.070 ;
        RECT -38.670 1870.290 -37.490 1871.470 ;
        RECT -37.070 1870.290 -35.890 1871.470 ;
        RECT -38.670 1691.890 -37.490 1693.070 ;
        RECT -37.070 1691.890 -35.890 1693.070 ;
        RECT -38.670 1690.290 -37.490 1691.470 ;
        RECT -37.070 1690.290 -35.890 1691.470 ;
        RECT -38.670 1511.890 -37.490 1513.070 ;
        RECT -37.070 1511.890 -35.890 1513.070 ;
        RECT -38.670 1510.290 -37.490 1511.470 ;
        RECT -37.070 1510.290 -35.890 1511.470 ;
        RECT -38.670 1331.890 -37.490 1333.070 ;
        RECT -37.070 1331.890 -35.890 1333.070 ;
        RECT -38.670 1330.290 -37.490 1331.470 ;
        RECT -37.070 1330.290 -35.890 1331.470 ;
        RECT -38.670 1151.890 -37.490 1153.070 ;
        RECT -37.070 1151.890 -35.890 1153.070 ;
        RECT -38.670 1150.290 -37.490 1151.470 ;
        RECT -37.070 1150.290 -35.890 1151.470 ;
        RECT -38.670 971.890 -37.490 973.070 ;
        RECT -37.070 971.890 -35.890 973.070 ;
        RECT -38.670 970.290 -37.490 971.470 ;
        RECT -37.070 970.290 -35.890 971.470 ;
        RECT -38.670 791.890 -37.490 793.070 ;
        RECT -37.070 791.890 -35.890 793.070 ;
        RECT -38.670 790.290 -37.490 791.470 ;
        RECT -37.070 790.290 -35.890 791.470 ;
        RECT -38.670 611.890 -37.490 613.070 ;
        RECT -37.070 611.890 -35.890 613.070 ;
        RECT -38.670 610.290 -37.490 611.470 ;
        RECT -37.070 610.290 -35.890 611.470 ;
        RECT -38.670 431.890 -37.490 433.070 ;
        RECT -37.070 431.890 -35.890 433.070 ;
        RECT -38.670 430.290 -37.490 431.470 ;
        RECT -37.070 430.290 -35.890 431.470 ;
        RECT -38.670 251.890 -37.490 253.070 ;
        RECT -37.070 251.890 -35.890 253.070 ;
        RECT -38.670 250.290 -37.490 251.470 ;
        RECT -37.070 250.290 -35.890 251.470 ;
        RECT -38.670 71.890 -37.490 73.070 ;
        RECT -37.070 71.890 -35.890 73.070 ;
        RECT -38.670 70.290 -37.490 71.470 ;
        RECT -37.070 70.290 -35.890 71.470 ;
        RECT -38.670 -31.710 -37.490 -30.530 ;
        RECT -37.070 -31.710 -35.890 -30.530 ;
        RECT -38.670 -33.310 -37.490 -32.130 ;
        RECT -37.070 -33.310 -35.890 -32.130 ;
        RECT 64.930 3551.810 66.110 3552.990 ;
        RECT 66.530 3551.810 67.710 3552.990 ;
        RECT 64.930 3550.210 66.110 3551.390 ;
        RECT 66.530 3550.210 67.710 3551.390 ;
        RECT 64.930 3491.890 66.110 3493.070 ;
        RECT 66.530 3491.890 67.710 3493.070 ;
        RECT 64.930 3490.290 66.110 3491.470 ;
        RECT 66.530 3490.290 67.710 3491.470 ;
        RECT 64.930 3311.890 66.110 3313.070 ;
        RECT 66.530 3311.890 67.710 3313.070 ;
        RECT 64.930 3310.290 66.110 3311.470 ;
        RECT 66.530 3310.290 67.710 3311.470 ;
        RECT 64.930 3131.890 66.110 3133.070 ;
        RECT 66.530 3131.890 67.710 3133.070 ;
        RECT 64.930 3130.290 66.110 3131.470 ;
        RECT 66.530 3130.290 67.710 3131.470 ;
        RECT 64.930 2951.890 66.110 2953.070 ;
        RECT 66.530 2951.890 67.710 2953.070 ;
        RECT 64.930 2950.290 66.110 2951.470 ;
        RECT 66.530 2950.290 67.710 2951.470 ;
        RECT 64.930 2771.890 66.110 2773.070 ;
        RECT 66.530 2771.890 67.710 2773.070 ;
        RECT 64.930 2770.290 66.110 2771.470 ;
        RECT 66.530 2770.290 67.710 2771.470 ;
        RECT 64.930 2591.890 66.110 2593.070 ;
        RECT 66.530 2591.890 67.710 2593.070 ;
        RECT 64.930 2590.290 66.110 2591.470 ;
        RECT 66.530 2590.290 67.710 2591.470 ;
        RECT 64.930 2411.890 66.110 2413.070 ;
        RECT 66.530 2411.890 67.710 2413.070 ;
        RECT 64.930 2410.290 66.110 2411.470 ;
        RECT 66.530 2410.290 67.710 2411.470 ;
        RECT 64.930 2231.890 66.110 2233.070 ;
        RECT 66.530 2231.890 67.710 2233.070 ;
        RECT 64.930 2230.290 66.110 2231.470 ;
        RECT 66.530 2230.290 67.710 2231.470 ;
        RECT 64.930 2051.890 66.110 2053.070 ;
        RECT 66.530 2051.890 67.710 2053.070 ;
        RECT 64.930 2050.290 66.110 2051.470 ;
        RECT 66.530 2050.290 67.710 2051.470 ;
        RECT 64.930 1871.890 66.110 1873.070 ;
        RECT 66.530 1871.890 67.710 1873.070 ;
        RECT 64.930 1870.290 66.110 1871.470 ;
        RECT 66.530 1870.290 67.710 1871.470 ;
        RECT 64.930 1691.890 66.110 1693.070 ;
        RECT 66.530 1691.890 67.710 1693.070 ;
        RECT 64.930 1690.290 66.110 1691.470 ;
        RECT 66.530 1690.290 67.710 1691.470 ;
        RECT 64.930 1511.890 66.110 1513.070 ;
        RECT 66.530 1511.890 67.710 1513.070 ;
        RECT 64.930 1510.290 66.110 1511.470 ;
        RECT 66.530 1510.290 67.710 1511.470 ;
        RECT 64.930 1331.890 66.110 1333.070 ;
        RECT 66.530 1331.890 67.710 1333.070 ;
        RECT 64.930 1330.290 66.110 1331.470 ;
        RECT 66.530 1330.290 67.710 1331.470 ;
        RECT 64.930 1151.890 66.110 1153.070 ;
        RECT 66.530 1151.890 67.710 1153.070 ;
        RECT 64.930 1150.290 66.110 1151.470 ;
        RECT 66.530 1150.290 67.710 1151.470 ;
        RECT 244.930 3551.810 246.110 3552.990 ;
        RECT 246.530 3551.810 247.710 3552.990 ;
        RECT 244.930 3550.210 246.110 3551.390 ;
        RECT 246.530 3550.210 247.710 3551.390 ;
        RECT 244.930 3491.890 246.110 3493.070 ;
        RECT 246.530 3491.890 247.710 3493.070 ;
        RECT 244.930 3490.290 246.110 3491.470 ;
        RECT 246.530 3490.290 247.710 3491.470 ;
        RECT 244.930 3311.890 246.110 3313.070 ;
        RECT 246.530 3311.890 247.710 3313.070 ;
        RECT 244.930 3310.290 246.110 3311.470 ;
        RECT 246.530 3310.290 247.710 3311.470 ;
        RECT 244.930 3131.890 246.110 3133.070 ;
        RECT 246.530 3131.890 247.710 3133.070 ;
        RECT 244.930 3130.290 246.110 3131.470 ;
        RECT 246.530 3130.290 247.710 3131.470 ;
        RECT 244.930 2951.890 246.110 2953.070 ;
        RECT 246.530 2951.890 247.710 2953.070 ;
        RECT 244.930 2950.290 246.110 2951.470 ;
        RECT 246.530 2950.290 247.710 2951.470 ;
        RECT 244.930 2771.890 246.110 2773.070 ;
        RECT 246.530 2771.890 247.710 2773.070 ;
        RECT 244.930 2770.290 246.110 2771.470 ;
        RECT 246.530 2770.290 247.710 2771.470 ;
        RECT 244.930 2591.890 246.110 2593.070 ;
        RECT 246.530 2591.890 247.710 2593.070 ;
        RECT 244.930 2590.290 246.110 2591.470 ;
        RECT 246.530 2590.290 247.710 2591.470 ;
        RECT 244.930 2411.890 246.110 2413.070 ;
        RECT 246.530 2411.890 247.710 2413.070 ;
        RECT 244.930 2410.290 246.110 2411.470 ;
        RECT 246.530 2410.290 247.710 2411.470 ;
        RECT 244.930 2231.890 246.110 2233.070 ;
        RECT 246.530 2231.890 247.710 2233.070 ;
        RECT 244.930 2230.290 246.110 2231.470 ;
        RECT 246.530 2230.290 247.710 2231.470 ;
        RECT 244.930 2051.890 246.110 2053.070 ;
        RECT 246.530 2051.890 247.710 2053.070 ;
        RECT 244.930 2050.290 246.110 2051.470 ;
        RECT 246.530 2050.290 247.710 2051.470 ;
        RECT 244.930 1871.890 246.110 1873.070 ;
        RECT 246.530 1871.890 247.710 1873.070 ;
        RECT 244.930 1870.290 246.110 1871.470 ;
        RECT 246.530 1870.290 247.710 1871.470 ;
        RECT 244.930 1691.890 246.110 1693.070 ;
        RECT 246.530 1691.890 247.710 1693.070 ;
        RECT 244.930 1690.290 246.110 1691.470 ;
        RECT 246.530 1690.290 247.710 1691.470 ;
        RECT 244.930 1511.890 246.110 1513.070 ;
        RECT 246.530 1511.890 247.710 1513.070 ;
        RECT 244.930 1510.290 246.110 1511.470 ;
        RECT 246.530 1510.290 247.710 1511.470 ;
        RECT 244.930 1331.890 246.110 1333.070 ;
        RECT 246.530 1331.890 247.710 1333.070 ;
        RECT 244.930 1330.290 246.110 1331.470 ;
        RECT 246.530 1330.290 247.710 1331.470 ;
        RECT 244.930 1151.890 246.110 1153.070 ;
        RECT 246.530 1151.890 247.710 1153.070 ;
        RECT 244.930 1150.290 246.110 1151.470 ;
        RECT 246.530 1150.290 247.710 1151.470 ;
        RECT 424.930 3551.810 426.110 3552.990 ;
        RECT 426.530 3551.810 427.710 3552.990 ;
        RECT 424.930 3550.210 426.110 3551.390 ;
        RECT 426.530 3550.210 427.710 3551.390 ;
        RECT 424.930 3491.890 426.110 3493.070 ;
        RECT 426.530 3491.890 427.710 3493.070 ;
        RECT 424.930 3490.290 426.110 3491.470 ;
        RECT 426.530 3490.290 427.710 3491.470 ;
        RECT 424.930 3311.890 426.110 3313.070 ;
        RECT 426.530 3311.890 427.710 3313.070 ;
        RECT 424.930 3310.290 426.110 3311.470 ;
        RECT 426.530 3310.290 427.710 3311.470 ;
        RECT 424.930 3131.890 426.110 3133.070 ;
        RECT 426.530 3131.890 427.710 3133.070 ;
        RECT 424.930 3130.290 426.110 3131.470 ;
        RECT 426.530 3130.290 427.710 3131.470 ;
        RECT 424.930 2951.890 426.110 2953.070 ;
        RECT 426.530 2951.890 427.710 2953.070 ;
        RECT 424.930 2950.290 426.110 2951.470 ;
        RECT 426.530 2950.290 427.710 2951.470 ;
        RECT 424.930 2771.890 426.110 2773.070 ;
        RECT 426.530 2771.890 427.710 2773.070 ;
        RECT 424.930 2770.290 426.110 2771.470 ;
        RECT 426.530 2770.290 427.710 2771.470 ;
        RECT 424.930 2591.890 426.110 2593.070 ;
        RECT 426.530 2591.890 427.710 2593.070 ;
        RECT 424.930 2590.290 426.110 2591.470 ;
        RECT 426.530 2590.290 427.710 2591.470 ;
        RECT 424.930 2411.890 426.110 2413.070 ;
        RECT 426.530 2411.890 427.710 2413.070 ;
        RECT 424.930 2410.290 426.110 2411.470 ;
        RECT 426.530 2410.290 427.710 2411.470 ;
        RECT 424.930 2231.890 426.110 2233.070 ;
        RECT 426.530 2231.890 427.710 2233.070 ;
        RECT 424.930 2230.290 426.110 2231.470 ;
        RECT 426.530 2230.290 427.710 2231.470 ;
        RECT 424.930 2051.890 426.110 2053.070 ;
        RECT 426.530 2051.890 427.710 2053.070 ;
        RECT 424.930 2050.290 426.110 2051.470 ;
        RECT 426.530 2050.290 427.710 2051.470 ;
        RECT 424.930 1871.890 426.110 1873.070 ;
        RECT 426.530 1871.890 427.710 1873.070 ;
        RECT 424.930 1870.290 426.110 1871.470 ;
        RECT 426.530 1870.290 427.710 1871.470 ;
        RECT 424.930 1691.890 426.110 1693.070 ;
        RECT 426.530 1691.890 427.710 1693.070 ;
        RECT 424.930 1690.290 426.110 1691.470 ;
        RECT 426.530 1690.290 427.710 1691.470 ;
        RECT 424.930 1511.890 426.110 1513.070 ;
        RECT 426.530 1511.890 427.710 1513.070 ;
        RECT 424.930 1510.290 426.110 1511.470 ;
        RECT 426.530 1510.290 427.710 1511.470 ;
        RECT 424.930 1331.890 426.110 1333.070 ;
        RECT 426.530 1331.890 427.710 1333.070 ;
        RECT 424.930 1330.290 426.110 1331.470 ;
        RECT 426.530 1330.290 427.710 1331.470 ;
        RECT 424.930 1151.890 426.110 1153.070 ;
        RECT 426.530 1151.890 427.710 1153.070 ;
        RECT 424.930 1150.290 426.110 1151.470 ;
        RECT 426.530 1150.290 427.710 1151.470 ;
        RECT 604.930 3551.810 606.110 3552.990 ;
        RECT 606.530 3551.810 607.710 3552.990 ;
        RECT 604.930 3550.210 606.110 3551.390 ;
        RECT 606.530 3550.210 607.710 3551.390 ;
        RECT 604.930 3491.890 606.110 3493.070 ;
        RECT 606.530 3491.890 607.710 3493.070 ;
        RECT 604.930 3490.290 606.110 3491.470 ;
        RECT 606.530 3490.290 607.710 3491.470 ;
        RECT 604.930 3311.890 606.110 3313.070 ;
        RECT 606.530 3311.890 607.710 3313.070 ;
        RECT 604.930 3310.290 606.110 3311.470 ;
        RECT 606.530 3310.290 607.710 3311.470 ;
        RECT 604.930 3131.890 606.110 3133.070 ;
        RECT 606.530 3131.890 607.710 3133.070 ;
        RECT 604.930 3130.290 606.110 3131.470 ;
        RECT 606.530 3130.290 607.710 3131.470 ;
        RECT 604.930 2951.890 606.110 2953.070 ;
        RECT 606.530 2951.890 607.710 2953.070 ;
        RECT 604.930 2950.290 606.110 2951.470 ;
        RECT 606.530 2950.290 607.710 2951.470 ;
        RECT 604.930 2771.890 606.110 2773.070 ;
        RECT 606.530 2771.890 607.710 2773.070 ;
        RECT 604.930 2770.290 606.110 2771.470 ;
        RECT 606.530 2770.290 607.710 2771.470 ;
        RECT 604.930 2591.890 606.110 2593.070 ;
        RECT 606.530 2591.890 607.710 2593.070 ;
        RECT 604.930 2590.290 606.110 2591.470 ;
        RECT 606.530 2590.290 607.710 2591.470 ;
        RECT 604.930 2411.890 606.110 2413.070 ;
        RECT 606.530 2411.890 607.710 2413.070 ;
        RECT 604.930 2410.290 606.110 2411.470 ;
        RECT 606.530 2410.290 607.710 2411.470 ;
        RECT 604.930 2231.890 606.110 2233.070 ;
        RECT 606.530 2231.890 607.710 2233.070 ;
        RECT 604.930 2230.290 606.110 2231.470 ;
        RECT 606.530 2230.290 607.710 2231.470 ;
        RECT 604.930 2051.890 606.110 2053.070 ;
        RECT 606.530 2051.890 607.710 2053.070 ;
        RECT 604.930 2050.290 606.110 2051.470 ;
        RECT 606.530 2050.290 607.710 2051.470 ;
        RECT 604.930 1871.890 606.110 1873.070 ;
        RECT 606.530 1871.890 607.710 1873.070 ;
        RECT 604.930 1870.290 606.110 1871.470 ;
        RECT 606.530 1870.290 607.710 1871.470 ;
        RECT 604.930 1691.890 606.110 1693.070 ;
        RECT 606.530 1691.890 607.710 1693.070 ;
        RECT 604.930 1690.290 606.110 1691.470 ;
        RECT 606.530 1690.290 607.710 1691.470 ;
        RECT 604.930 1511.890 606.110 1513.070 ;
        RECT 606.530 1511.890 607.710 1513.070 ;
        RECT 604.930 1510.290 606.110 1511.470 ;
        RECT 606.530 1510.290 607.710 1511.470 ;
        RECT 604.930 1331.890 606.110 1333.070 ;
        RECT 606.530 1331.890 607.710 1333.070 ;
        RECT 604.930 1330.290 606.110 1331.470 ;
        RECT 606.530 1330.290 607.710 1331.470 ;
        RECT 604.930 1151.890 606.110 1153.070 ;
        RECT 606.530 1151.890 607.710 1153.070 ;
        RECT 604.930 1150.290 606.110 1151.470 ;
        RECT 606.530 1150.290 607.710 1151.470 ;
        RECT 784.930 3551.810 786.110 3552.990 ;
        RECT 786.530 3551.810 787.710 3552.990 ;
        RECT 784.930 3550.210 786.110 3551.390 ;
        RECT 786.530 3550.210 787.710 3551.390 ;
        RECT 784.930 3491.890 786.110 3493.070 ;
        RECT 786.530 3491.890 787.710 3493.070 ;
        RECT 784.930 3490.290 786.110 3491.470 ;
        RECT 786.530 3490.290 787.710 3491.470 ;
        RECT 784.930 3311.890 786.110 3313.070 ;
        RECT 786.530 3311.890 787.710 3313.070 ;
        RECT 784.930 3310.290 786.110 3311.470 ;
        RECT 786.530 3310.290 787.710 3311.470 ;
        RECT 784.930 3131.890 786.110 3133.070 ;
        RECT 786.530 3131.890 787.710 3133.070 ;
        RECT 784.930 3130.290 786.110 3131.470 ;
        RECT 786.530 3130.290 787.710 3131.470 ;
        RECT 784.930 2951.890 786.110 2953.070 ;
        RECT 786.530 2951.890 787.710 2953.070 ;
        RECT 784.930 2950.290 786.110 2951.470 ;
        RECT 786.530 2950.290 787.710 2951.470 ;
        RECT 784.930 2771.890 786.110 2773.070 ;
        RECT 786.530 2771.890 787.710 2773.070 ;
        RECT 784.930 2770.290 786.110 2771.470 ;
        RECT 786.530 2770.290 787.710 2771.470 ;
        RECT 784.930 2591.890 786.110 2593.070 ;
        RECT 786.530 2591.890 787.710 2593.070 ;
        RECT 784.930 2590.290 786.110 2591.470 ;
        RECT 786.530 2590.290 787.710 2591.470 ;
        RECT 784.930 2411.890 786.110 2413.070 ;
        RECT 786.530 2411.890 787.710 2413.070 ;
        RECT 784.930 2410.290 786.110 2411.470 ;
        RECT 786.530 2410.290 787.710 2411.470 ;
        RECT 784.930 2231.890 786.110 2233.070 ;
        RECT 786.530 2231.890 787.710 2233.070 ;
        RECT 784.930 2230.290 786.110 2231.470 ;
        RECT 786.530 2230.290 787.710 2231.470 ;
        RECT 784.930 2051.890 786.110 2053.070 ;
        RECT 786.530 2051.890 787.710 2053.070 ;
        RECT 784.930 2050.290 786.110 2051.470 ;
        RECT 786.530 2050.290 787.710 2051.470 ;
        RECT 784.930 1871.890 786.110 1873.070 ;
        RECT 786.530 1871.890 787.710 1873.070 ;
        RECT 784.930 1870.290 786.110 1871.470 ;
        RECT 786.530 1870.290 787.710 1871.470 ;
        RECT 784.930 1691.890 786.110 1693.070 ;
        RECT 786.530 1691.890 787.710 1693.070 ;
        RECT 784.930 1690.290 786.110 1691.470 ;
        RECT 786.530 1690.290 787.710 1691.470 ;
        RECT 784.930 1511.890 786.110 1513.070 ;
        RECT 786.530 1511.890 787.710 1513.070 ;
        RECT 784.930 1510.290 786.110 1511.470 ;
        RECT 786.530 1510.290 787.710 1511.470 ;
        RECT 784.930 1331.890 786.110 1333.070 ;
        RECT 786.530 1331.890 787.710 1333.070 ;
        RECT 784.930 1330.290 786.110 1331.470 ;
        RECT 786.530 1330.290 787.710 1331.470 ;
        RECT 784.930 1151.890 786.110 1153.070 ;
        RECT 786.530 1151.890 787.710 1153.070 ;
        RECT 784.930 1150.290 786.110 1151.470 ;
        RECT 786.530 1150.290 787.710 1151.470 ;
        RECT 964.930 3551.810 966.110 3552.990 ;
        RECT 966.530 3551.810 967.710 3552.990 ;
        RECT 964.930 3550.210 966.110 3551.390 ;
        RECT 966.530 3550.210 967.710 3551.390 ;
        RECT 964.930 3491.890 966.110 3493.070 ;
        RECT 966.530 3491.890 967.710 3493.070 ;
        RECT 964.930 3490.290 966.110 3491.470 ;
        RECT 966.530 3490.290 967.710 3491.470 ;
        RECT 964.930 3311.890 966.110 3313.070 ;
        RECT 966.530 3311.890 967.710 3313.070 ;
        RECT 964.930 3310.290 966.110 3311.470 ;
        RECT 966.530 3310.290 967.710 3311.470 ;
        RECT 964.930 3131.890 966.110 3133.070 ;
        RECT 966.530 3131.890 967.710 3133.070 ;
        RECT 964.930 3130.290 966.110 3131.470 ;
        RECT 966.530 3130.290 967.710 3131.470 ;
        RECT 964.930 2951.890 966.110 2953.070 ;
        RECT 966.530 2951.890 967.710 2953.070 ;
        RECT 964.930 2950.290 966.110 2951.470 ;
        RECT 966.530 2950.290 967.710 2951.470 ;
        RECT 964.930 2771.890 966.110 2773.070 ;
        RECT 966.530 2771.890 967.710 2773.070 ;
        RECT 964.930 2770.290 966.110 2771.470 ;
        RECT 966.530 2770.290 967.710 2771.470 ;
        RECT 964.930 2591.890 966.110 2593.070 ;
        RECT 966.530 2591.890 967.710 2593.070 ;
        RECT 964.930 2590.290 966.110 2591.470 ;
        RECT 966.530 2590.290 967.710 2591.470 ;
        RECT 964.930 2411.890 966.110 2413.070 ;
        RECT 966.530 2411.890 967.710 2413.070 ;
        RECT 964.930 2410.290 966.110 2411.470 ;
        RECT 966.530 2410.290 967.710 2411.470 ;
        RECT 964.930 2231.890 966.110 2233.070 ;
        RECT 966.530 2231.890 967.710 2233.070 ;
        RECT 964.930 2230.290 966.110 2231.470 ;
        RECT 966.530 2230.290 967.710 2231.470 ;
        RECT 964.930 2051.890 966.110 2053.070 ;
        RECT 966.530 2051.890 967.710 2053.070 ;
        RECT 964.930 2050.290 966.110 2051.470 ;
        RECT 966.530 2050.290 967.710 2051.470 ;
        RECT 964.930 1871.890 966.110 1873.070 ;
        RECT 966.530 1871.890 967.710 1873.070 ;
        RECT 964.930 1870.290 966.110 1871.470 ;
        RECT 966.530 1870.290 967.710 1871.470 ;
        RECT 964.930 1691.890 966.110 1693.070 ;
        RECT 966.530 1691.890 967.710 1693.070 ;
        RECT 964.930 1690.290 966.110 1691.470 ;
        RECT 966.530 1690.290 967.710 1691.470 ;
        RECT 964.930 1511.890 966.110 1513.070 ;
        RECT 966.530 1511.890 967.710 1513.070 ;
        RECT 964.930 1510.290 966.110 1511.470 ;
        RECT 966.530 1510.290 967.710 1511.470 ;
        RECT 964.930 1331.890 966.110 1333.070 ;
        RECT 966.530 1331.890 967.710 1333.070 ;
        RECT 964.930 1330.290 966.110 1331.470 ;
        RECT 966.530 1330.290 967.710 1331.470 ;
        RECT 964.930 1151.890 966.110 1153.070 ;
        RECT 966.530 1151.890 967.710 1153.070 ;
        RECT 964.930 1150.290 966.110 1151.470 ;
        RECT 966.530 1150.290 967.710 1151.470 ;
        RECT 1144.930 3551.810 1146.110 3552.990 ;
        RECT 1146.530 3551.810 1147.710 3552.990 ;
        RECT 1144.930 3550.210 1146.110 3551.390 ;
        RECT 1146.530 3550.210 1147.710 3551.390 ;
        RECT 1144.930 3491.890 1146.110 3493.070 ;
        RECT 1146.530 3491.890 1147.710 3493.070 ;
        RECT 1144.930 3490.290 1146.110 3491.470 ;
        RECT 1146.530 3490.290 1147.710 3491.470 ;
        RECT 1144.930 3311.890 1146.110 3313.070 ;
        RECT 1146.530 3311.890 1147.710 3313.070 ;
        RECT 1144.930 3310.290 1146.110 3311.470 ;
        RECT 1146.530 3310.290 1147.710 3311.470 ;
        RECT 1144.930 3131.890 1146.110 3133.070 ;
        RECT 1146.530 3131.890 1147.710 3133.070 ;
        RECT 1144.930 3130.290 1146.110 3131.470 ;
        RECT 1146.530 3130.290 1147.710 3131.470 ;
        RECT 1144.930 2951.890 1146.110 2953.070 ;
        RECT 1146.530 2951.890 1147.710 2953.070 ;
        RECT 1144.930 2950.290 1146.110 2951.470 ;
        RECT 1146.530 2950.290 1147.710 2951.470 ;
        RECT 1144.930 2771.890 1146.110 2773.070 ;
        RECT 1146.530 2771.890 1147.710 2773.070 ;
        RECT 1144.930 2770.290 1146.110 2771.470 ;
        RECT 1146.530 2770.290 1147.710 2771.470 ;
        RECT 1144.930 2591.890 1146.110 2593.070 ;
        RECT 1146.530 2591.890 1147.710 2593.070 ;
        RECT 1144.930 2590.290 1146.110 2591.470 ;
        RECT 1146.530 2590.290 1147.710 2591.470 ;
        RECT 1144.930 2411.890 1146.110 2413.070 ;
        RECT 1146.530 2411.890 1147.710 2413.070 ;
        RECT 1144.930 2410.290 1146.110 2411.470 ;
        RECT 1146.530 2410.290 1147.710 2411.470 ;
        RECT 1144.930 2231.890 1146.110 2233.070 ;
        RECT 1146.530 2231.890 1147.710 2233.070 ;
        RECT 1144.930 2230.290 1146.110 2231.470 ;
        RECT 1146.530 2230.290 1147.710 2231.470 ;
        RECT 1144.930 2051.890 1146.110 2053.070 ;
        RECT 1146.530 2051.890 1147.710 2053.070 ;
        RECT 1144.930 2050.290 1146.110 2051.470 ;
        RECT 1146.530 2050.290 1147.710 2051.470 ;
        RECT 1144.930 1871.890 1146.110 1873.070 ;
        RECT 1146.530 1871.890 1147.710 1873.070 ;
        RECT 1144.930 1870.290 1146.110 1871.470 ;
        RECT 1146.530 1870.290 1147.710 1871.470 ;
        RECT 1144.930 1691.890 1146.110 1693.070 ;
        RECT 1146.530 1691.890 1147.710 1693.070 ;
        RECT 1144.930 1690.290 1146.110 1691.470 ;
        RECT 1146.530 1690.290 1147.710 1691.470 ;
        RECT 1144.930 1511.890 1146.110 1513.070 ;
        RECT 1146.530 1511.890 1147.710 1513.070 ;
        RECT 1144.930 1510.290 1146.110 1511.470 ;
        RECT 1146.530 1510.290 1147.710 1511.470 ;
        RECT 1144.930 1331.890 1146.110 1333.070 ;
        RECT 1146.530 1331.890 1147.710 1333.070 ;
        RECT 1144.930 1330.290 1146.110 1331.470 ;
        RECT 1146.530 1330.290 1147.710 1331.470 ;
        RECT 1144.930 1151.890 1146.110 1153.070 ;
        RECT 1146.530 1151.890 1147.710 1153.070 ;
        RECT 1144.930 1150.290 1146.110 1151.470 ;
        RECT 1146.530 1150.290 1147.710 1151.470 ;
        RECT 64.930 971.890 66.110 973.070 ;
        RECT 66.530 971.890 67.710 973.070 ;
        RECT 64.930 970.290 66.110 971.470 ;
        RECT 66.530 970.290 67.710 971.470 ;
        RECT 64.930 791.890 66.110 793.070 ;
        RECT 66.530 791.890 67.710 793.070 ;
        RECT 64.930 790.290 66.110 791.470 ;
        RECT 66.530 790.290 67.710 791.470 ;
        RECT 64.930 611.890 66.110 613.070 ;
        RECT 66.530 611.890 67.710 613.070 ;
        RECT 64.930 610.290 66.110 611.470 ;
        RECT 66.530 610.290 67.710 611.470 ;
        RECT 64.930 431.890 66.110 433.070 ;
        RECT 66.530 431.890 67.710 433.070 ;
        RECT 64.930 430.290 66.110 431.470 ;
        RECT 66.530 430.290 67.710 431.470 ;
        RECT 1144.930 971.890 1146.110 973.070 ;
        RECT 1146.530 971.890 1147.710 973.070 ;
        RECT 1144.930 970.290 1146.110 971.470 ;
        RECT 1146.530 970.290 1147.710 971.470 ;
        RECT 1144.930 791.890 1146.110 793.070 ;
        RECT 1146.530 791.890 1147.710 793.070 ;
        RECT 1144.930 790.290 1146.110 791.470 ;
        RECT 1146.530 790.290 1147.710 791.470 ;
        RECT 1144.930 611.890 1146.110 613.070 ;
        RECT 1146.530 611.890 1147.710 613.070 ;
        RECT 1144.930 610.290 1146.110 611.470 ;
        RECT 1146.530 610.290 1147.710 611.470 ;
        RECT 1144.930 431.890 1146.110 433.070 ;
        RECT 1146.530 431.890 1147.710 433.070 ;
        RECT 1144.930 430.290 1146.110 431.470 ;
        RECT 1146.530 430.290 1147.710 431.470 ;
        RECT 64.930 251.890 66.110 253.070 ;
        RECT 66.530 251.890 67.710 253.070 ;
        RECT 64.930 250.290 66.110 251.470 ;
        RECT 66.530 250.290 67.710 251.470 ;
        RECT 64.930 71.890 66.110 73.070 ;
        RECT 66.530 71.890 67.710 73.070 ;
        RECT 64.930 70.290 66.110 71.470 ;
        RECT 66.530 70.290 67.710 71.470 ;
        RECT 64.930 -31.710 66.110 -30.530 ;
        RECT 66.530 -31.710 67.710 -30.530 ;
        RECT 64.930 -33.310 66.110 -32.130 ;
        RECT 66.530 -33.310 67.710 -32.130 ;
        RECT 244.930 251.890 246.110 253.070 ;
        RECT 246.530 251.890 247.710 253.070 ;
        RECT 244.930 250.290 246.110 251.470 ;
        RECT 246.530 250.290 247.710 251.470 ;
        RECT 244.930 71.890 246.110 73.070 ;
        RECT 246.530 71.890 247.710 73.070 ;
        RECT 244.930 70.290 246.110 71.470 ;
        RECT 246.530 70.290 247.710 71.470 ;
        RECT 244.930 -31.710 246.110 -30.530 ;
        RECT 246.530 -31.710 247.710 -30.530 ;
        RECT 244.930 -33.310 246.110 -32.130 ;
        RECT 246.530 -33.310 247.710 -32.130 ;
        RECT 424.930 251.890 426.110 253.070 ;
        RECT 426.530 251.890 427.710 253.070 ;
        RECT 424.930 250.290 426.110 251.470 ;
        RECT 426.530 250.290 427.710 251.470 ;
        RECT 424.930 71.890 426.110 73.070 ;
        RECT 426.530 71.890 427.710 73.070 ;
        RECT 424.930 70.290 426.110 71.470 ;
        RECT 426.530 70.290 427.710 71.470 ;
        RECT 424.930 -31.710 426.110 -30.530 ;
        RECT 426.530 -31.710 427.710 -30.530 ;
        RECT 424.930 -33.310 426.110 -32.130 ;
        RECT 426.530 -33.310 427.710 -32.130 ;
        RECT 604.930 251.890 606.110 253.070 ;
        RECT 606.530 251.890 607.710 253.070 ;
        RECT 604.930 250.290 606.110 251.470 ;
        RECT 606.530 250.290 607.710 251.470 ;
        RECT 604.930 71.890 606.110 73.070 ;
        RECT 606.530 71.890 607.710 73.070 ;
        RECT 604.930 70.290 606.110 71.470 ;
        RECT 606.530 70.290 607.710 71.470 ;
        RECT 604.930 -31.710 606.110 -30.530 ;
        RECT 606.530 -31.710 607.710 -30.530 ;
        RECT 604.930 -33.310 606.110 -32.130 ;
        RECT 606.530 -33.310 607.710 -32.130 ;
        RECT 784.930 251.890 786.110 253.070 ;
        RECT 786.530 251.890 787.710 253.070 ;
        RECT 784.930 250.290 786.110 251.470 ;
        RECT 786.530 250.290 787.710 251.470 ;
        RECT 784.930 71.890 786.110 73.070 ;
        RECT 786.530 71.890 787.710 73.070 ;
        RECT 784.930 70.290 786.110 71.470 ;
        RECT 786.530 70.290 787.710 71.470 ;
        RECT 784.930 -31.710 786.110 -30.530 ;
        RECT 786.530 -31.710 787.710 -30.530 ;
        RECT 784.930 -33.310 786.110 -32.130 ;
        RECT 786.530 -33.310 787.710 -32.130 ;
        RECT 964.930 251.890 966.110 253.070 ;
        RECT 966.530 251.890 967.710 253.070 ;
        RECT 964.930 250.290 966.110 251.470 ;
        RECT 966.530 250.290 967.710 251.470 ;
        RECT 964.930 71.890 966.110 73.070 ;
        RECT 966.530 71.890 967.710 73.070 ;
        RECT 964.930 70.290 966.110 71.470 ;
        RECT 966.530 70.290 967.710 71.470 ;
        RECT 964.930 -31.710 966.110 -30.530 ;
        RECT 966.530 -31.710 967.710 -30.530 ;
        RECT 964.930 -33.310 966.110 -32.130 ;
        RECT 966.530 -33.310 967.710 -32.130 ;
        RECT 1144.930 251.890 1146.110 253.070 ;
        RECT 1146.530 251.890 1147.710 253.070 ;
        RECT 1144.930 250.290 1146.110 251.470 ;
        RECT 1146.530 250.290 1147.710 251.470 ;
        RECT 1144.930 71.890 1146.110 73.070 ;
        RECT 1146.530 71.890 1147.710 73.070 ;
        RECT 1144.930 70.290 1146.110 71.470 ;
        RECT 1146.530 70.290 1147.710 71.470 ;
        RECT 1144.930 -31.710 1146.110 -30.530 ;
        RECT 1146.530 -31.710 1147.710 -30.530 ;
        RECT 1144.930 -33.310 1146.110 -32.130 ;
        RECT 1146.530 -33.310 1147.710 -32.130 ;
        RECT 1324.930 3551.810 1326.110 3552.990 ;
        RECT 1326.530 3551.810 1327.710 3552.990 ;
        RECT 1324.930 3550.210 1326.110 3551.390 ;
        RECT 1326.530 3550.210 1327.710 3551.390 ;
        RECT 1324.930 3491.890 1326.110 3493.070 ;
        RECT 1326.530 3491.890 1327.710 3493.070 ;
        RECT 1324.930 3490.290 1326.110 3491.470 ;
        RECT 1326.530 3490.290 1327.710 3491.470 ;
        RECT 1324.930 3311.890 1326.110 3313.070 ;
        RECT 1326.530 3311.890 1327.710 3313.070 ;
        RECT 1324.930 3310.290 1326.110 3311.470 ;
        RECT 1326.530 3310.290 1327.710 3311.470 ;
        RECT 1324.930 3131.890 1326.110 3133.070 ;
        RECT 1326.530 3131.890 1327.710 3133.070 ;
        RECT 1324.930 3130.290 1326.110 3131.470 ;
        RECT 1326.530 3130.290 1327.710 3131.470 ;
        RECT 1324.930 2951.890 1326.110 2953.070 ;
        RECT 1326.530 2951.890 1327.710 2953.070 ;
        RECT 1324.930 2950.290 1326.110 2951.470 ;
        RECT 1326.530 2950.290 1327.710 2951.470 ;
        RECT 1324.930 2771.890 1326.110 2773.070 ;
        RECT 1326.530 2771.890 1327.710 2773.070 ;
        RECT 1324.930 2770.290 1326.110 2771.470 ;
        RECT 1326.530 2770.290 1327.710 2771.470 ;
        RECT 1324.930 2591.890 1326.110 2593.070 ;
        RECT 1326.530 2591.890 1327.710 2593.070 ;
        RECT 1324.930 2590.290 1326.110 2591.470 ;
        RECT 1326.530 2590.290 1327.710 2591.470 ;
        RECT 1324.930 2411.890 1326.110 2413.070 ;
        RECT 1326.530 2411.890 1327.710 2413.070 ;
        RECT 1324.930 2410.290 1326.110 2411.470 ;
        RECT 1326.530 2410.290 1327.710 2411.470 ;
        RECT 1324.930 2231.890 1326.110 2233.070 ;
        RECT 1326.530 2231.890 1327.710 2233.070 ;
        RECT 1324.930 2230.290 1326.110 2231.470 ;
        RECT 1326.530 2230.290 1327.710 2231.470 ;
        RECT 1324.930 2051.890 1326.110 2053.070 ;
        RECT 1326.530 2051.890 1327.710 2053.070 ;
        RECT 1324.930 2050.290 1326.110 2051.470 ;
        RECT 1326.530 2050.290 1327.710 2051.470 ;
        RECT 1324.930 1871.890 1326.110 1873.070 ;
        RECT 1326.530 1871.890 1327.710 1873.070 ;
        RECT 1324.930 1870.290 1326.110 1871.470 ;
        RECT 1326.530 1870.290 1327.710 1871.470 ;
        RECT 1324.930 1691.890 1326.110 1693.070 ;
        RECT 1326.530 1691.890 1327.710 1693.070 ;
        RECT 1324.930 1690.290 1326.110 1691.470 ;
        RECT 1326.530 1690.290 1327.710 1691.470 ;
        RECT 1324.930 1511.890 1326.110 1513.070 ;
        RECT 1326.530 1511.890 1327.710 1513.070 ;
        RECT 1324.930 1510.290 1326.110 1511.470 ;
        RECT 1326.530 1510.290 1327.710 1511.470 ;
        RECT 1324.930 1331.890 1326.110 1333.070 ;
        RECT 1326.530 1331.890 1327.710 1333.070 ;
        RECT 1324.930 1330.290 1326.110 1331.470 ;
        RECT 1326.530 1330.290 1327.710 1331.470 ;
        RECT 1324.930 1151.890 1326.110 1153.070 ;
        RECT 1326.530 1151.890 1327.710 1153.070 ;
        RECT 1324.930 1150.290 1326.110 1151.470 ;
        RECT 1326.530 1150.290 1327.710 1151.470 ;
        RECT 1324.930 971.890 1326.110 973.070 ;
        RECT 1326.530 971.890 1327.710 973.070 ;
        RECT 1324.930 970.290 1326.110 971.470 ;
        RECT 1326.530 970.290 1327.710 971.470 ;
        RECT 1324.930 791.890 1326.110 793.070 ;
        RECT 1326.530 791.890 1327.710 793.070 ;
        RECT 1324.930 790.290 1326.110 791.470 ;
        RECT 1326.530 790.290 1327.710 791.470 ;
        RECT 1324.930 611.890 1326.110 613.070 ;
        RECT 1326.530 611.890 1327.710 613.070 ;
        RECT 1324.930 610.290 1326.110 611.470 ;
        RECT 1326.530 610.290 1327.710 611.470 ;
        RECT 1324.930 431.890 1326.110 433.070 ;
        RECT 1326.530 431.890 1327.710 433.070 ;
        RECT 1324.930 430.290 1326.110 431.470 ;
        RECT 1326.530 430.290 1327.710 431.470 ;
        RECT 1324.930 251.890 1326.110 253.070 ;
        RECT 1326.530 251.890 1327.710 253.070 ;
        RECT 1324.930 250.290 1326.110 251.470 ;
        RECT 1326.530 250.290 1327.710 251.470 ;
        RECT 1324.930 71.890 1326.110 73.070 ;
        RECT 1326.530 71.890 1327.710 73.070 ;
        RECT 1324.930 70.290 1326.110 71.470 ;
        RECT 1326.530 70.290 1327.710 71.470 ;
        RECT 1324.930 -31.710 1326.110 -30.530 ;
        RECT 1326.530 -31.710 1327.710 -30.530 ;
        RECT 1324.930 -33.310 1326.110 -32.130 ;
        RECT 1326.530 -33.310 1327.710 -32.130 ;
        RECT 1504.930 3551.810 1506.110 3552.990 ;
        RECT 1506.530 3551.810 1507.710 3552.990 ;
        RECT 1504.930 3550.210 1506.110 3551.390 ;
        RECT 1506.530 3550.210 1507.710 3551.390 ;
        RECT 1504.930 3491.890 1506.110 3493.070 ;
        RECT 1506.530 3491.890 1507.710 3493.070 ;
        RECT 1504.930 3490.290 1506.110 3491.470 ;
        RECT 1506.530 3490.290 1507.710 3491.470 ;
        RECT 1504.930 3311.890 1506.110 3313.070 ;
        RECT 1506.530 3311.890 1507.710 3313.070 ;
        RECT 1504.930 3310.290 1506.110 3311.470 ;
        RECT 1506.530 3310.290 1507.710 3311.470 ;
        RECT 1504.930 3131.890 1506.110 3133.070 ;
        RECT 1506.530 3131.890 1507.710 3133.070 ;
        RECT 1504.930 3130.290 1506.110 3131.470 ;
        RECT 1506.530 3130.290 1507.710 3131.470 ;
        RECT 1504.930 2951.890 1506.110 2953.070 ;
        RECT 1506.530 2951.890 1507.710 2953.070 ;
        RECT 1504.930 2950.290 1506.110 2951.470 ;
        RECT 1506.530 2950.290 1507.710 2951.470 ;
        RECT 1504.930 2771.890 1506.110 2773.070 ;
        RECT 1506.530 2771.890 1507.710 2773.070 ;
        RECT 1504.930 2770.290 1506.110 2771.470 ;
        RECT 1506.530 2770.290 1507.710 2771.470 ;
        RECT 1504.930 2591.890 1506.110 2593.070 ;
        RECT 1506.530 2591.890 1507.710 2593.070 ;
        RECT 1504.930 2590.290 1506.110 2591.470 ;
        RECT 1506.530 2590.290 1507.710 2591.470 ;
        RECT 1504.930 2411.890 1506.110 2413.070 ;
        RECT 1506.530 2411.890 1507.710 2413.070 ;
        RECT 1504.930 2410.290 1506.110 2411.470 ;
        RECT 1506.530 2410.290 1507.710 2411.470 ;
        RECT 1504.930 2231.890 1506.110 2233.070 ;
        RECT 1506.530 2231.890 1507.710 2233.070 ;
        RECT 1504.930 2230.290 1506.110 2231.470 ;
        RECT 1506.530 2230.290 1507.710 2231.470 ;
        RECT 1504.930 2051.890 1506.110 2053.070 ;
        RECT 1506.530 2051.890 1507.710 2053.070 ;
        RECT 1504.930 2050.290 1506.110 2051.470 ;
        RECT 1506.530 2050.290 1507.710 2051.470 ;
        RECT 1504.930 1871.890 1506.110 1873.070 ;
        RECT 1506.530 1871.890 1507.710 1873.070 ;
        RECT 1504.930 1870.290 1506.110 1871.470 ;
        RECT 1506.530 1870.290 1507.710 1871.470 ;
        RECT 1504.930 1691.890 1506.110 1693.070 ;
        RECT 1506.530 1691.890 1507.710 1693.070 ;
        RECT 1504.930 1690.290 1506.110 1691.470 ;
        RECT 1506.530 1690.290 1507.710 1691.470 ;
        RECT 1504.930 1511.890 1506.110 1513.070 ;
        RECT 1506.530 1511.890 1507.710 1513.070 ;
        RECT 1504.930 1510.290 1506.110 1511.470 ;
        RECT 1506.530 1510.290 1507.710 1511.470 ;
        RECT 1504.930 1331.890 1506.110 1333.070 ;
        RECT 1506.530 1331.890 1507.710 1333.070 ;
        RECT 1504.930 1330.290 1506.110 1331.470 ;
        RECT 1506.530 1330.290 1507.710 1331.470 ;
        RECT 1504.930 1151.890 1506.110 1153.070 ;
        RECT 1506.530 1151.890 1507.710 1153.070 ;
        RECT 1504.930 1150.290 1506.110 1151.470 ;
        RECT 1506.530 1150.290 1507.710 1151.470 ;
        RECT 1504.930 971.890 1506.110 973.070 ;
        RECT 1506.530 971.890 1507.710 973.070 ;
        RECT 1504.930 970.290 1506.110 971.470 ;
        RECT 1506.530 970.290 1507.710 971.470 ;
        RECT 1504.930 791.890 1506.110 793.070 ;
        RECT 1506.530 791.890 1507.710 793.070 ;
        RECT 1504.930 790.290 1506.110 791.470 ;
        RECT 1506.530 790.290 1507.710 791.470 ;
        RECT 1504.930 611.890 1506.110 613.070 ;
        RECT 1506.530 611.890 1507.710 613.070 ;
        RECT 1504.930 610.290 1506.110 611.470 ;
        RECT 1506.530 610.290 1507.710 611.470 ;
        RECT 1504.930 431.890 1506.110 433.070 ;
        RECT 1506.530 431.890 1507.710 433.070 ;
        RECT 1504.930 430.290 1506.110 431.470 ;
        RECT 1506.530 430.290 1507.710 431.470 ;
        RECT 1504.930 251.890 1506.110 253.070 ;
        RECT 1506.530 251.890 1507.710 253.070 ;
        RECT 1504.930 250.290 1506.110 251.470 ;
        RECT 1506.530 250.290 1507.710 251.470 ;
        RECT 1504.930 71.890 1506.110 73.070 ;
        RECT 1506.530 71.890 1507.710 73.070 ;
        RECT 1504.930 70.290 1506.110 71.470 ;
        RECT 1506.530 70.290 1507.710 71.470 ;
        RECT 1504.930 -31.710 1506.110 -30.530 ;
        RECT 1506.530 -31.710 1507.710 -30.530 ;
        RECT 1504.930 -33.310 1506.110 -32.130 ;
        RECT 1506.530 -33.310 1507.710 -32.130 ;
        RECT 1684.930 3551.810 1686.110 3552.990 ;
        RECT 1686.530 3551.810 1687.710 3552.990 ;
        RECT 1684.930 3550.210 1686.110 3551.390 ;
        RECT 1686.530 3550.210 1687.710 3551.390 ;
        RECT 1684.930 3491.890 1686.110 3493.070 ;
        RECT 1686.530 3491.890 1687.710 3493.070 ;
        RECT 1684.930 3490.290 1686.110 3491.470 ;
        RECT 1686.530 3490.290 1687.710 3491.470 ;
        RECT 1684.930 3311.890 1686.110 3313.070 ;
        RECT 1686.530 3311.890 1687.710 3313.070 ;
        RECT 1684.930 3310.290 1686.110 3311.470 ;
        RECT 1686.530 3310.290 1687.710 3311.470 ;
        RECT 1684.930 3131.890 1686.110 3133.070 ;
        RECT 1686.530 3131.890 1687.710 3133.070 ;
        RECT 1684.930 3130.290 1686.110 3131.470 ;
        RECT 1686.530 3130.290 1687.710 3131.470 ;
        RECT 1684.930 2951.890 1686.110 2953.070 ;
        RECT 1686.530 2951.890 1687.710 2953.070 ;
        RECT 1684.930 2950.290 1686.110 2951.470 ;
        RECT 1686.530 2950.290 1687.710 2951.470 ;
        RECT 1684.930 2771.890 1686.110 2773.070 ;
        RECT 1686.530 2771.890 1687.710 2773.070 ;
        RECT 1684.930 2770.290 1686.110 2771.470 ;
        RECT 1686.530 2770.290 1687.710 2771.470 ;
        RECT 1684.930 2591.890 1686.110 2593.070 ;
        RECT 1686.530 2591.890 1687.710 2593.070 ;
        RECT 1684.930 2590.290 1686.110 2591.470 ;
        RECT 1686.530 2590.290 1687.710 2591.470 ;
        RECT 1684.930 2411.890 1686.110 2413.070 ;
        RECT 1686.530 2411.890 1687.710 2413.070 ;
        RECT 1684.930 2410.290 1686.110 2411.470 ;
        RECT 1686.530 2410.290 1687.710 2411.470 ;
        RECT 1684.930 2231.890 1686.110 2233.070 ;
        RECT 1686.530 2231.890 1687.710 2233.070 ;
        RECT 1684.930 2230.290 1686.110 2231.470 ;
        RECT 1686.530 2230.290 1687.710 2231.470 ;
        RECT 1684.930 2051.890 1686.110 2053.070 ;
        RECT 1686.530 2051.890 1687.710 2053.070 ;
        RECT 1684.930 2050.290 1686.110 2051.470 ;
        RECT 1686.530 2050.290 1687.710 2051.470 ;
        RECT 1684.930 1871.890 1686.110 1873.070 ;
        RECT 1686.530 1871.890 1687.710 1873.070 ;
        RECT 1684.930 1870.290 1686.110 1871.470 ;
        RECT 1686.530 1870.290 1687.710 1871.470 ;
        RECT 1684.930 1691.890 1686.110 1693.070 ;
        RECT 1686.530 1691.890 1687.710 1693.070 ;
        RECT 1684.930 1690.290 1686.110 1691.470 ;
        RECT 1686.530 1690.290 1687.710 1691.470 ;
        RECT 1684.930 1511.890 1686.110 1513.070 ;
        RECT 1686.530 1511.890 1687.710 1513.070 ;
        RECT 1684.930 1510.290 1686.110 1511.470 ;
        RECT 1686.530 1510.290 1687.710 1511.470 ;
        RECT 1684.930 1331.890 1686.110 1333.070 ;
        RECT 1686.530 1331.890 1687.710 1333.070 ;
        RECT 1684.930 1330.290 1686.110 1331.470 ;
        RECT 1686.530 1330.290 1687.710 1331.470 ;
        RECT 1684.930 1151.890 1686.110 1153.070 ;
        RECT 1686.530 1151.890 1687.710 1153.070 ;
        RECT 1684.930 1150.290 1686.110 1151.470 ;
        RECT 1686.530 1150.290 1687.710 1151.470 ;
        RECT 1684.930 971.890 1686.110 973.070 ;
        RECT 1686.530 971.890 1687.710 973.070 ;
        RECT 1684.930 970.290 1686.110 971.470 ;
        RECT 1686.530 970.290 1687.710 971.470 ;
        RECT 1684.930 791.890 1686.110 793.070 ;
        RECT 1686.530 791.890 1687.710 793.070 ;
        RECT 1684.930 790.290 1686.110 791.470 ;
        RECT 1686.530 790.290 1687.710 791.470 ;
        RECT 1684.930 611.890 1686.110 613.070 ;
        RECT 1686.530 611.890 1687.710 613.070 ;
        RECT 1684.930 610.290 1686.110 611.470 ;
        RECT 1686.530 610.290 1687.710 611.470 ;
        RECT 1684.930 431.890 1686.110 433.070 ;
        RECT 1686.530 431.890 1687.710 433.070 ;
        RECT 1684.930 430.290 1686.110 431.470 ;
        RECT 1686.530 430.290 1687.710 431.470 ;
        RECT 1684.930 251.890 1686.110 253.070 ;
        RECT 1686.530 251.890 1687.710 253.070 ;
        RECT 1684.930 250.290 1686.110 251.470 ;
        RECT 1686.530 250.290 1687.710 251.470 ;
        RECT 1684.930 71.890 1686.110 73.070 ;
        RECT 1686.530 71.890 1687.710 73.070 ;
        RECT 1684.930 70.290 1686.110 71.470 ;
        RECT 1686.530 70.290 1687.710 71.470 ;
        RECT 1684.930 -31.710 1686.110 -30.530 ;
        RECT 1686.530 -31.710 1687.710 -30.530 ;
        RECT 1684.930 -33.310 1686.110 -32.130 ;
        RECT 1686.530 -33.310 1687.710 -32.130 ;
        RECT 1864.930 3551.810 1866.110 3552.990 ;
        RECT 1866.530 3551.810 1867.710 3552.990 ;
        RECT 1864.930 3550.210 1866.110 3551.390 ;
        RECT 1866.530 3550.210 1867.710 3551.390 ;
        RECT 1864.930 3491.890 1866.110 3493.070 ;
        RECT 1866.530 3491.890 1867.710 3493.070 ;
        RECT 1864.930 3490.290 1866.110 3491.470 ;
        RECT 1866.530 3490.290 1867.710 3491.470 ;
        RECT 1864.930 3311.890 1866.110 3313.070 ;
        RECT 1866.530 3311.890 1867.710 3313.070 ;
        RECT 1864.930 3310.290 1866.110 3311.470 ;
        RECT 1866.530 3310.290 1867.710 3311.470 ;
        RECT 1864.930 3131.890 1866.110 3133.070 ;
        RECT 1866.530 3131.890 1867.710 3133.070 ;
        RECT 1864.930 3130.290 1866.110 3131.470 ;
        RECT 1866.530 3130.290 1867.710 3131.470 ;
        RECT 1864.930 2951.890 1866.110 2953.070 ;
        RECT 1866.530 2951.890 1867.710 2953.070 ;
        RECT 1864.930 2950.290 1866.110 2951.470 ;
        RECT 1866.530 2950.290 1867.710 2951.470 ;
        RECT 1864.930 2771.890 1866.110 2773.070 ;
        RECT 1866.530 2771.890 1867.710 2773.070 ;
        RECT 1864.930 2770.290 1866.110 2771.470 ;
        RECT 1866.530 2770.290 1867.710 2771.470 ;
        RECT 1864.930 2591.890 1866.110 2593.070 ;
        RECT 1866.530 2591.890 1867.710 2593.070 ;
        RECT 1864.930 2590.290 1866.110 2591.470 ;
        RECT 1866.530 2590.290 1867.710 2591.470 ;
        RECT 1864.930 2411.890 1866.110 2413.070 ;
        RECT 1866.530 2411.890 1867.710 2413.070 ;
        RECT 1864.930 2410.290 1866.110 2411.470 ;
        RECT 1866.530 2410.290 1867.710 2411.470 ;
        RECT 1864.930 2231.890 1866.110 2233.070 ;
        RECT 1866.530 2231.890 1867.710 2233.070 ;
        RECT 1864.930 2230.290 1866.110 2231.470 ;
        RECT 1866.530 2230.290 1867.710 2231.470 ;
        RECT 1864.930 2051.890 1866.110 2053.070 ;
        RECT 1866.530 2051.890 1867.710 2053.070 ;
        RECT 1864.930 2050.290 1866.110 2051.470 ;
        RECT 1866.530 2050.290 1867.710 2051.470 ;
        RECT 1864.930 1871.890 1866.110 1873.070 ;
        RECT 1866.530 1871.890 1867.710 1873.070 ;
        RECT 1864.930 1870.290 1866.110 1871.470 ;
        RECT 1866.530 1870.290 1867.710 1871.470 ;
        RECT 1864.930 1691.890 1866.110 1693.070 ;
        RECT 1866.530 1691.890 1867.710 1693.070 ;
        RECT 1864.930 1690.290 1866.110 1691.470 ;
        RECT 1866.530 1690.290 1867.710 1691.470 ;
        RECT 1864.930 1511.890 1866.110 1513.070 ;
        RECT 1866.530 1511.890 1867.710 1513.070 ;
        RECT 1864.930 1510.290 1866.110 1511.470 ;
        RECT 1866.530 1510.290 1867.710 1511.470 ;
        RECT 1864.930 1331.890 1866.110 1333.070 ;
        RECT 1866.530 1331.890 1867.710 1333.070 ;
        RECT 1864.930 1330.290 1866.110 1331.470 ;
        RECT 1866.530 1330.290 1867.710 1331.470 ;
        RECT 1864.930 1151.890 1866.110 1153.070 ;
        RECT 1866.530 1151.890 1867.710 1153.070 ;
        RECT 1864.930 1150.290 1866.110 1151.470 ;
        RECT 1866.530 1150.290 1867.710 1151.470 ;
        RECT 1864.930 971.890 1866.110 973.070 ;
        RECT 1866.530 971.890 1867.710 973.070 ;
        RECT 1864.930 970.290 1866.110 971.470 ;
        RECT 1866.530 970.290 1867.710 971.470 ;
        RECT 1864.930 791.890 1866.110 793.070 ;
        RECT 1866.530 791.890 1867.710 793.070 ;
        RECT 1864.930 790.290 1866.110 791.470 ;
        RECT 1866.530 790.290 1867.710 791.470 ;
        RECT 1864.930 611.890 1866.110 613.070 ;
        RECT 1866.530 611.890 1867.710 613.070 ;
        RECT 1864.930 610.290 1866.110 611.470 ;
        RECT 1866.530 610.290 1867.710 611.470 ;
        RECT 1864.930 431.890 1866.110 433.070 ;
        RECT 1866.530 431.890 1867.710 433.070 ;
        RECT 1864.930 430.290 1866.110 431.470 ;
        RECT 1866.530 430.290 1867.710 431.470 ;
        RECT 1864.930 251.890 1866.110 253.070 ;
        RECT 1866.530 251.890 1867.710 253.070 ;
        RECT 1864.930 250.290 1866.110 251.470 ;
        RECT 1866.530 250.290 1867.710 251.470 ;
        RECT 1864.930 71.890 1866.110 73.070 ;
        RECT 1866.530 71.890 1867.710 73.070 ;
        RECT 1864.930 70.290 1866.110 71.470 ;
        RECT 1866.530 70.290 1867.710 71.470 ;
        RECT 1864.930 -31.710 1866.110 -30.530 ;
        RECT 1866.530 -31.710 1867.710 -30.530 ;
        RECT 1864.930 -33.310 1866.110 -32.130 ;
        RECT 1866.530 -33.310 1867.710 -32.130 ;
        RECT 2044.930 3551.810 2046.110 3552.990 ;
        RECT 2046.530 3551.810 2047.710 3552.990 ;
        RECT 2044.930 3550.210 2046.110 3551.390 ;
        RECT 2046.530 3550.210 2047.710 3551.390 ;
        RECT 2044.930 3491.890 2046.110 3493.070 ;
        RECT 2046.530 3491.890 2047.710 3493.070 ;
        RECT 2044.930 3490.290 2046.110 3491.470 ;
        RECT 2046.530 3490.290 2047.710 3491.470 ;
        RECT 2044.930 3311.890 2046.110 3313.070 ;
        RECT 2046.530 3311.890 2047.710 3313.070 ;
        RECT 2044.930 3310.290 2046.110 3311.470 ;
        RECT 2046.530 3310.290 2047.710 3311.470 ;
        RECT 2044.930 3131.890 2046.110 3133.070 ;
        RECT 2046.530 3131.890 2047.710 3133.070 ;
        RECT 2044.930 3130.290 2046.110 3131.470 ;
        RECT 2046.530 3130.290 2047.710 3131.470 ;
        RECT 2044.930 2951.890 2046.110 2953.070 ;
        RECT 2046.530 2951.890 2047.710 2953.070 ;
        RECT 2044.930 2950.290 2046.110 2951.470 ;
        RECT 2046.530 2950.290 2047.710 2951.470 ;
        RECT 2044.930 2771.890 2046.110 2773.070 ;
        RECT 2046.530 2771.890 2047.710 2773.070 ;
        RECT 2044.930 2770.290 2046.110 2771.470 ;
        RECT 2046.530 2770.290 2047.710 2771.470 ;
        RECT 2044.930 2591.890 2046.110 2593.070 ;
        RECT 2046.530 2591.890 2047.710 2593.070 ;
        RECT 2044.930 2590.290 2046.110 2591.470 ;
        RECT 2046.530 2590.290 2047.710 2591.470 ;
        RECT 2044.930 2411.890 2046.110 2413.070 ;
        RECT 2046.530 2411.890 2047.710 2413.070 ;
        RECT 2044.930 2410.290 2046.110 2411.470 ;
        RECT 2046.530 2410.290 2047.710 2411.470 ;
        RECT 2044.930 2231.890 2046.110 2233.070 ;
        RECT 2046.530 2231.890 2047.710 2233.070 ;
        RECT 2044.930 2230.290 2046.110 2231.470 ;
        RECT 2046.530 2230.290 2047.710 2231.470 ;
        RECT 2044.930 2051.890 2046.110 2053.070 ;
        RECT 2046.530 2051.890 2047.710 2053.070 ;
        RECT 2044.930 2050.290 2046.110 2051.470 ;
        RECT 2046.530 2050.290 2047.710 2051.470 ;
        RECT 2044.930 1871.890 2046.110 1873.070 ;
        RECT 2046.530 1871.890 2047.710 1873.070 ;
        RECT 2044.930 1870.290 2046.110 1871.470 ;
        RECT 2046.530 1870.290 2047.710 1871.470 ;
        RECT 2044.930 1691.890 2046.110 1693.070 ;
        RECT 2046.530 1691.890 2047.710 1693.070 ;
        RECT 2044.930 1690.290 2046.110 1691.470 ;
        RECT 2046.530 1690.290 2047.710 1691.470 ;
        RECT 2044.930 1511.890 2046.110 1513.070 ;
        RECT 2046.530 1511.890 2047.710 1513.070 ;
        RECT 2044.930 1510.290 2046.110 1511.470 ;
        RECT 2046.530 1510.290 2047.710 1511.470 ;
        RECT 2044.930 1331.890 2046.110 1333.070 ;
        RECT 2046.530 1331.890 2047.710 1333.070 ;
        RECT 2044.930 1330.290 2046.110 1331.470 ;
        RECT 2046.530 1330.290 2047.710 1331.470 ;
        RECT 2044.930 1151.890 2046.110 1153.070 ;
        RECT 2046.530 1151.890 2047.710 1153.070 ;
        RECT 2044.930 1150.290 2046.110 1151.470 ;
        RECT 2046.530 1150.290 2047.710 1151.470 ;
        RECT 2044.930 971.890 2046.110 973.070 ;
        RECT 2046.530 971.890 2047.710 973.070 ;
        RECT 2044.930 970.290 2046.110 971.470 ;
        RECT 2046.530 970.290 2047.710 971.470 ;
        RECT 2044.930 791.890 2046.110 793.070 ;
        RECT 2046.530 791.890 2047.710 793.070 ;
        RECT 2044.930 790.290 2046.110 791.470 ;
        RECT 2046.530 790.290 2047.710 791.470 ;
        RECT 2044.930 611.890 2046.110 613.070 ;
        RECT 2046.530 611.890 2047.710 613.070 ;
        RECT 2044.930 610.290 2046.110 611.470 ;
        RECT 2046.530 610.290 2047.710 611.470 ;
        RECT 2044.930 431.890 2046.110 433.070 ;
        RECT 2046.530 431.890 2047.710 433.070 ;
        RECT 2044.930 430.290 2046.110 431.470 ;
        RECT 2046.530 430.290 2047.710 431.470 ;
        RECT 2044.930 251.890 2046.110 253.070 ;
        RECT 2046.530 251.890 2047.710 253.070 ;
        RECT 2044.930 250.290 2046.110 251.470 ;
        RECT 2046.530 250.290 2047.710 251.470 ;
        RECT 2044.930 71.890 2046.110 73.070 ;
        RECT 2046.530 71.890 2047.710 73.070 ;
        RECT 2044.930 70.290 2046.110 71.470 ;
        RECT 2046.530 70.290 2047.710 71.470 ;
        RECT 2044.930 -31.710 2046.110 -30.530 ;
        RECT 2046.530 -31.710 2047.710 -30.530 ;
        RECT 2044.930 -33.310 2046.110 -32.130 ;
        RECT 2046.530 -33.310 2047.710 -32.130 ;
        RECT 2224.930 3551.810 2226.110 3552.990 ;
        RECT 2226.530 3551.810 2227.710 3552.990 ;
        RECT 2224.930 3550.210 2226.110 3551.390 ;
        RECT 2226.530 3550.210 2227.710 3551.390 ;
        RECT 2224.930 3491.890 2226.110 3493.070 ;
        RECT 2226.530 3491.890 2227.710 3493.070 ;
        RECT 2224.930 3490.290 2226.110 3491.470 ;
        RECT 2226.530 3490.290 2227.710 3491.470 ;
        RECT 2224.930 3311.890 2226.110 3313.070 ;
        RECT 2226.530 3311.890 2227.710 3313.070 ;
        RECT 2224.930 3310.290 2226.110 3311.470 ;
        RECT 2226.530 3310.290 2227.710 3311.470 ;
        RECT 2224.930 3131.890 2226.110 3133.070 ;
        RECT 2226.530 3131.890 2227.710 3133.070 ;
        RECT 2224.930 3130.290 2226.110 3131.470 ;
        RECT 2226.530 3130.290 2227.710 3131.470 ;
        RECT 2224.930 2951.890 2226.110 2953.070 ;
        RECT 2226.530 2951.890 2227.710 2953.070 ;
        RECT 2224.930 2950.290 2226.110 2951.470 ;
        RECT 2226.530 2950.290 2227.710 2951.470 ;
        RECT 2224.930 2771.890 2226.110 2773.070 ;
        RECT 2226.530 2771.890 2227.710 2773.070 ;
        RECT 2224.930 2770.290 2226.110 2771.470 ;
        RECT 2226.530 2770.290 2227.710 2771.470 ;
        RECT 2224.930 2591.890 2226.110 2593.070 ;
        RECT 2226.530 2591.890 2227.710 2593.070 ;
        RECT 2224.930 2590.290 2226.110 2591.470 ;
        RECT 2226.530 2590.290 2227.710 2591.470 ;
        RECT 2224.930 2411.890 2226.110 2413.070 ;
        RECT 2226.530 2411.890 2227.710 2413.070 ;
        RECT 2224.930 2410.290 2226.110 2411.470 ;
        RECT 2226.530 2410.290 2227.710 2411.470 ;
        RECT 2224.930 2231.890 2226.110 2233.070 ;
        RECT 2226.530 2231.890 2227.710 2233.070 ;
        RECT 2224.930 2230.290 2226.110 2231.470 ;
        RECT 2226.530 2230.290 2227.710 2231.470 ;
        RECT 2224.930 2051.890 2226.110 2053.070 ;
        RECT 2226.530 2051.890 2227.710 2053.070 ;
        RECT 2224.930 2050.290 2226.110 2051.470 ;
        RECT 2226.530 2050.290 2227.710 2051.470 ;
        RECT 2224.930 1871.890 2226.110 1873.070 ;
        RECT 2226.530 1871.890 2227.710 1873.070 ;
        RECT 2224.930 1870.290 2226.110 1871.470 ;
        RECT 2226.530 1870.290 2227.710 1871.470 ;
        RECT 2224.930 1691.890 2226.110 1693.070 ;
        RECT 2226.530 1691.890 2227.710 1693.070 ;
        RECT 2224.930 1690.290 2226.110 1691.470 ;
        RECT 2226.530 1690.290 2227.710 1691.470 ;
        RECT 2224.930 1511.890 2226.110 1513.070 ;
        RECT 2226.530 1511.890 2227.710 1513.070 ;
        RECT 2224.930 1510.290 2226.110 1511.470 ;
        RECT 2226.530 1510.290 2227.710 1511.470 ;
        RECT 2224.930 1331.890 2226.110 1333.070 ;
        RECT 2226.530 1331.890 2227.710 1333.070 ;
        RECT 2224.930 1330.290 2226.110 1331.470 ;
        RECT 2226.530 1330.290 2227.710 1331.470 ;
        RECT 2224.930 1151.890 2226.110 1153.070 ;
        RECT 2226.530 1151.890 2227.710 1153.070 ;
        RECT 2224.930 1150.290 2226.110 1151.470 ;
        RECT 2226.530 1150.290 2227.710 1151.470 ;
        RECT 2224.930 971.890 2226.110 973.070 ;
        RECT 2226.530 971.890 2227.710 973.070 ;
        RECT 2224.930 970.290 2226.110 971.470 ;
        RECT 2226.530 970.290 2227.710 971.470 ;
        RECT 2224.930 791.890 2226.110 793.070 ;
        RECT 2226.530 791.890 2227.710 793.070 ;
        RECT 2224.930 790.290 2226.110 791.470 ;
        RECT 2226.530 790.290 2227.710 791.470 ;
        RECT 2224.930 611.890 2226.110 613.070 ;
        RECT 2226.530 611.890 2227.710 613.070 ;
        RECT 2224.930 610.290 2226.110 611.470 ;
        RECT 2226.530 610.290 2227.710 611.470 ;
        RECT 2224.930 431.890 2226.110 433.070 ;
        RECT 2226.530 431.890 2227.710 433.070 ;
        RECT 2224.930 430.290 2226.110 431.470 ;
        RECT 2226.530 430.290 2227.710 431.470 ;
        RECT 2224.930 251.890 2226.110 253.070 ;
        RECT 2226.530 251.890 2227.710 253.070 ;
        RECT 2224.930 250.290 2226.110 251.470 ;
        RECT 2226.530 250.290 2227.710 251.470 ;
        RECT 2224.930 71.890 2226.110 73.070 ;
        RECT 2226.530 71.890 2227.710 73.070 ;
        RECT 2224.930 70.290 2226.110 71.470 ;
        RECT 2226.530 70.290 2227.710 71.470 ;
        RECT 2224.930 -31.710 2226.110 -30.530 ;
        RECT 2226.530 -31.710 2227.710 -30.530 ;
        RECT 2224.930 -33.310 2226.110 -32.130 ;
        RECT 2226.530 -33.310 2227.710 -32.130 ;
        RECT 2404.930 3551.810 2406.110 3552.990 ;
        RECT 2406.530 3551.810 2407.710 3552.990 ;
        RECT 2404.930 3550.210 2406.110 3551.390 ;
        RECT 2406.530 3550.210 2407.710 3551.390 ;
        RECT 2404.930 3491.890 2406.110 3493.070 ;
        RECT 2406.530 3491.890 2407.710 3493.070 ;
        RECT 2404.930 3490.290 2406.110 3491.470 ;
        RECT 2406.530 3490.290 2407.710 3491.470 ;
        RECT 2404.930 3311.890 2406.110 3313.070 ;
        RECT 2406.530 3311.890 2407.710 3313.070 ;
        RECT 2404.930 3310.290 2406.110 3311.470 ;
        RECT 2406.530 3310.290 2407.710 3311.470 ;
        RECT 2404.930 3131.890 2406.110 3133.070 ;
        RECT 2406.530 3131.890 2407.710 3133.070 ;
        RECT 2404.930 3130.290 2406.110 3131.470 ;
        RECT 2406.530 3130.290 2407.710 3131.470 ;
        RECT 2404.930 2951.890 2406.110 2953.070 ;
        RECT 2406.530 2951.890 2407.710 2953.070 ;
        RECT 2404.930 2950.290 2406.110 2951.470 ;
        RECT 2406.530 2950.290 2407.710 2951.470 ;
        RECT 2404.930 2771.890 2406.110 2773.070 ;
        RECT 2406.530 2771.890 2407.710 2773.070 ;
        RECT 2404.930 2770.290 2406.110 2771.470 ;
        RECT 2406.530 2770.290 2407.710 2771.470 ;
        RECT 2404.930 2591.890 2406.110 2593.070 ;
        RECT 2406.530 2591.890 2407.710 2593.070 ;
        RECT 2404.930 2590.290 2406.110 2591.470 ;
        RECT 2406.530 2590.290 2407.710 2591.470 ;
        RECT 2404.930 2411.890 2406.110 2413.070 ;
        RECT 2406.530 2411.890 2407.710 2413.070 ;
        RECT 2404.930 2410.290 2406.110 2411.470 ;
        RECT 2406.530 2410.290 2407.710 2411.470 ;
        RECT 2404.930 2231.890 2406.110 2233.070 ;
        RECT 2406.530 2231.890 2407.710 2233.070 ;
        RECT 2404.930 2230.290 2406.110 2231.470 ;
        RECT 2406.530 2230.290 2407.710 2231.470 ;
        RECT 2404.930 2051.890 2406.110 2053.070 ;
        RECT 2406.530 2051.890 2407.710 2053.070 ;
        RECT 2404.930 2050.290 2406.110 2051.470 ;
        RECT 2406.530 2050.290 2407.710 2051.470 ;
        RECT 2404.930 1871.890 2406.110 1873.070 ;
        RECT 2406.530 1871.890 2407.710 1873.070 ;
        RECT 2404.930 1870.290 2406.110 1871.470 ;
        RECT 2406.530 1870.290 2407.710 1871.470 ;
        RECT 2404.930 1691.890 2406.110 1693.070 ;
        RECT 2406.530 1691.890 2407.710 1693.070 ;
        RECT 2404.930 1690.290 2406.110 1691.470 ;
        RECT 2406.530 1690.290 2407.710 1691.470 ;
        RECT 2404.930 1511.890 2406.110 1513.070 ;
        RECT 2406.530 1511.890 2407.710 1513.070 ;
        RECT 2404.930 1510.290 2406.110 1511.470 ;
        RECT 2406.530 1510.290 2407.710 1511.470 ;
        RECT 2404.930 1331.890 2406.110 1333.070 ;
        RECT 2406.530 1331.890 2407.710 1333.070 ;
        RECT 2404.930 1330.290 2406.110 1331.470 ;
        RECT 2406.530 1330.290 2407.710 1331.470 ;
        RECT 2404.930 1151.890 2406.110 1153.070 ;
        RECT 2406.530 1151.890 2407.710 1153.070 ;
        RECT 2404.930 1150.290 2406.110 1151.470 ;
        RECT 2406.530 1150.290 2407.710 1151.470 ;
        RECT 2404.930 971.890 2406.110 973.070 ;
        RECT 2406.530 971.890 2407.710 973.070 ;
        RECT 2404.930 970.290 2406.110 971.470 ;
        RECT 2406.530 970.290 2407.710 971.470 ;
        RECT 2404.930 791.890 2406.110 793.070 ;
        RECT 2406.530 791.890 2407.710 793.070 ;
        RECT 2404.930 790.290 2406.110 791.470 ;
        RECT 2406.530 790.290 2407.710 791.470 ;
        RECT 2404.930 611.890 2406.110 613.070 ;
        RECT 2406.530 611.890 2407.710 613.070 ;
        RECT 2404.930 610.290 2406.110 611.470 ;
        RECT 2406.530 610.290 2407.710 611.470 ;
        RECT 2404.930 431.890 2406.110 433.070 ;
        RECT 2406.530 431.890 2407.710 433.070 ;
        RECT 2404.930 430.290 2406.110 431.470 ;
        RECT 2406.530 430.290 2407.710 431.470 ;
        RECT 2404.930 251.890 2406.110 253.070 ;
        RECT 2406.530 251.890 2407.710 253.070 ;
        RECT 2404.930 250.290 2406.110 251.470 ;
        RECT 2406.530 250.290 2407.710 251.470 ;
        RECT 2404.930 71.890 2406.110 73.070 ;
        RECT 2406.530 71.890 2407.710 73.070 ;
        RECT 2404.930 70.290 2406.110 71.470 ;
        RECT 2406.530 70.290 2407.710 71.470 ;
        RECT 2404.930 -31.710 2406.110 -30.530 ;
        RECT 2406.530 -31.710 2407.710 -30.530 ;
        RECT 2404.930 -33.310 2406.110 -32.130 ;
        RECT 2406.530 -33.310 2407.710 -32.130 ;
        RECT 2584.930 3551.810 2586.110 3552.990 ;
        RECT 2586.530 3551.810 2587.710 3552.990 ;
        RECT 2584.930 3550.210 2586.110 3551.390 ;
        RECT 2586.530 3550.210 2587.710 3551.390 ;
        RECT 2584.930 3491.890 2586.110 3493.070 ;
        RECT 2586.530 3491.890 2587.710 3493.070 ;
        RECT 2584.930 3490.290 2586.110 3491.470 ;
        RECT 2586.530 3490.290 2587.710 3491.470 ;
        RECT 2584.930 3311.890 2586.110 3313.070 ;
        RECT 2586.530 3311.890 2587.710 3313.070 ;
        RECT 2584.930 3310.290 2586.110 3311.470 ;
        RECT 2586.530 3310.290 2587.710 3311.470 ;
        RECT 2584.930 3131.890 2586.110 3133.070 ;
        RECT 2586.530 3131.890 2587.710 3133.070 ;
        RECT 2584.930 3130.290 2586.110 3131.470 ;
        RECT 2586.530 3130.290 2587.710 3131.470 ;
        RECT 2584.930 2951.890 2586.110 2953.070 ;
        RECT 2586.530 2951.890 2587.710 2953.070 ;
        RECT 2584.930 2950.290 2586.110 2951.470 ;
        RECT 2586.530 2950.290 2587.710 2951.470 ;
        RECT 2584.930 2771.890 2586.110 2773.070 ;
        RECT 2586.530 2771.890 2587.710 2773.070 ;
        RECT 2584.930 2770.290 2586.110 2771.470 ;
        RECT 2586.530 2770.290 2587.710 2771.470 ;
        RECT 2584.930 2591.890 2586.110 2593.070 ;
        RECT 2586.530 2591.890 2587.710 2593.070 ;
        RECT 2584.930 2590.290 2586.110 2591.470 ;
        RECT 2586.530 2590.290 2587.710 2591.470 ;
        RECT 2584.930 2411.890 2586.110 2413.070 ;
        RECT 2586.530 2411.890 2587.710 2413.070 ;
        RECT 2584.930 2410.290 2586.110 2411.470 ;
        RECT 2586.530 2410.290 2587.710 2411.470 ;
        RECT 2584.930 2231.890 2586.110 2233.070 ;
        RECT 2586.530 2231.890 2587.710 2233.070 ;
        RECT 2584.930 2230.290 2586.110 2231.470 ;
        RECT 2586.530 2230.290 2587.710 2231.470 ;
        RECT 2584.930 2051.890 2586.110 2053.070 ;
        RECT 2586.530 2051.890 2587.710 2053.070 ;
        RECT 2584.930 2050.290 2586.110 2051.470 ;
        RECT 2586.530 2050.290 2587.710 2051.470 ;
        RECT 2584.930 1871.890 2586.110 1873.070 ;
        RECT 2586.530 1871.890 2587.710 1873.070 ;
        RECT 2584.930 1870.290 2586.110 1871.470 ;
        RECT 2586.530 1870.290 2587.710 1871.470 ;
        RECT 2584.930 1691.890 2586.110 1693.070 ;
        RECT 2586.530 1691.890 2587.710 1693.070 ;
        RECT 2584.930 1690.290 2586.110 1691.470 ;
        RECT 2586.530 1690.290 2587.710 1691.470 ;
        RECT 2584.930 1511.890 2586.110 1513.070 ;
        RECT 2586.530 1511.890 2587.710 1513.070 ;
        RECT 2584.930 1510.290 2586.110 1511.470 ;
        RECT 2586.530 1510.290 2587.710 1511.470 ;
        RECT 2584.930 1331.890 2586.110 1333.070 ;
        RECT 2586.530 1331.890 2587.710 1333.070 ;
        RECT 2584.930 1330.290 2586.110 1331.470 ;
        RECT 2586.530 1330.290 2587.710 1331.470 ;
        RECT 2584.930 1151.890 2586.110 1153.070 ;
        RECT 2586.530 1151.890 2587.710 1153.070 ;
        RECT 2584.930 1150.290 2586.110 1151.470 ;
        RECT 2586.530 1150.290 2587.710 1151.470 ;
        RECT 2584.930 971.890 2586.110 973.070 ;
        RECT 2586.530 971.890 2587.710 973.070 ;
        RECT 2584.930 970.290 2586.110 971.470 ;
        RECT 2586.530 970.290 2587.710 971.470 ;
        RECT 2584.930 791.890 2586.110 793.070 ;
        RECT 2586.530 791.890 2587.710 793.070 ;
        RECT 2584.930 790.290 2586.110 791.470 ;
        RECT 2586.530 790.290 2587.710 791.470 ;
        RECT 2584.930 611.890 2586.110 613.070 ;
        RECT 2586.530 611.890 2587.710 613.070 ;
        RECT 2584.930 610.290 2586.110 611.470 ;
        RECT 2586.530 610.290 2587.710 611.470 ;
        RECT 2584.930 431.890 2586.110 433.070 ;
        RECT 2586.530 431.890 2587.710 433.070 ;
        RECT 2584.930 430.290 2586.110 431.470 ;
        RECT 2586.530 430.290 2587.710 431.470 ;
        RECT 2584.930 251.890 2586.110 253.070 ;
        RECT 2586.530 251.890 2587.710 253.070 ;
        RECT 2584.930 250.290 2586.110 251.470 ;
        RECT 2586.530 250.290 2587.710 251.470 ;
        RECT 2584.930 71.890 2586.110 73.070 ;
        RECT 2586.530 71.890 2587.710 73.070 ;
        RECT 2584.930 70.290 2586.110 71.470 ;
        RECT 2586.530 70.290 2587.710 71.470 ;
        RECT 2584.930 -31.710 2586.110 -30.530 ;
        RECT 2586.530 -31.710 2587.710 -30.530 ;
        RECT 2584.930 -33.310 2586.110 -32.130 ;
        RECT 2586.530 -33.310 2587.710 -32.130 ;
        RECT 2764.930 3551.810 2766.110 3552.990 ;
        RECT 2766.530 3551.810 2767.710 3552.990 ;
        RECT 2764.930 3550.210 2766.110 3551.390 ;
        RECT 2766.530 3550.210 2767.710 3551.390 ;
        RECT 2764.930 3491.890 2766.110 3493.070 ;
        RECT 2766.530 3491.890 2767.710 3493.070 ;
        RECT 2764.930 3490.290 2766.110 3491.470 ;
        RECT 2766.530 3490.290 2767.710 3491.470 ;
        RECT 2764.930 3311.890 2766.110 3313.070 ;
        RECT 2766.530 3311.890 2767.710 3313.070 ;
        RECT 2764.930 3310.290 2766.110 3311.470 ;
        RECT 2766.530 3310.290 2767.710 3311.470 ;
        RECT 2764.930 3131.890 2766.110 3133.070 ;
        RECT 2766.530 3131.890 2767.710 3133.070 ;
        RECT 2764.930 3130.290 2766.110 3131.470 ;
        RECT 2766.530 3130.290 2767.710 3131.470 ;
        RECT 2764.930 2951.890 2766.110 2953.070 ;
        RECT 2766.530 2951.890 2767.710 2953.070 ;
        RECT 2764.930 2950.290 2766.110 2951.470 ;
        RECT 2766.530 2950.290 2767.710 2951.470 ;
        RECT 2764.930 2771.890 2766.110 2773.070 ;
        RECT 2766.530 2771.890 2767.710 2773.070 ;
        RECT 2764.930 2770.290 2766.110 2771.470 ;
        RECT 2766.530 2770.290 2767.710 2771.470 ;
        RECT 2764.930 2591.890 2766.110 2593.070 ;
        RECT 2766.530 2591.890 2767.710 2593.070 ;
        RECT 2764.930 2590.290 2766.110 2591.470 ;
        RECT 2766.530 2590.290 2767.710 2591.470 ;
        RECT 2764.930 2411.890 2766.110 2413.070 ;
        RECT 2766.530 2411.890 2767.710 2413.070 ;
        RECT 2764.930 2410.290 2766.110 2411.470 ;
        RECT 2766.530 2410.290 2767.710 2411.470 ;
        RECT 2764.930 2231.890 2766.110 2233.070 ;
        RECT 2766.530 2231.890 2767.710 2233.070 ;
        RECT 2764.930 2230.290 2766.110 2231.470 ;
        RECT 2766.530 2230.290 2767.710 2231.470 ;
        RECT 2764.930 2051.890 2766.110 2053.070 ;
        RECT 2766.530 2051.890 2767.710 2053.070 ;
        RECT 2764.930 2050.290 2766.110 2051.470 ;
        RECT 2766.530 2050.290 2767.710 2051.470 ;
        RECT 2764.930 1871.890 2766.110 1873.070 ;
        RECT 2766.530 1871.890 2767.710 1873.070 ;
        RECT 2764.930 1870.290 2766.110 1871.470 ;
        RECT 2766.530 1870.290 2767.710 1871.470 ;
        RECT 2764.930 1691.890 2766.110 1693.070 ;
        RECT 2766.530 1691.890 2767.710 1693.070 ;
        RECT 2764.930 1690.290 2766.110 1691.470 ;
        RECT 2766.530 1690.290 2767.710 1691.470 ;
        RECT 2764.930 1511.890 2766.110 1513.070 ;
        RECT 2766.530 1511.890 2767.710 1513.070 ;
        RECT 2764.930 1510.290 2766.110 1511.470 ;
        RECT 2766.530 1510.290 2767.710 1511.470 ;
        RECT 2764.930 1331.890 2766.110 1333.070 ;
        RECT 2766.530 1331.890 2767.710 1333.070 ;
        RECT 2764.930 1330.290 2766.110 1331.470 ;
        RECT 2766.530 1330.290 2767.710 1331.470 ;
        RECT 2764.930 1151.890 2766.110 1153.070 ;
        RECT 2766.530 1151.890 2767.710 1153.070 ;
        RECT 2764.930 1150.290 2766.110 1151.470 ;
        RECT 2766.530 1150.290 2767.710 1151.470 ;
        RECT 2764.930 971.890 2766.110 973.070 ;
        RECT 2766.530 971.890 2767.710 973.070 ;
        RECT 2764.930 970.290 2766.110 971.470 ;
        RECT 2766.530 970.290 2767.710 971.470 ;
        RECT 2764.930 791.890 2766.110 793.070 ;
        RECT 2766.530 791.890 2767.710 793.070 ;
        RECT 2764.930 790.290 2766.110 791.470 ;
        RECT 2766.530 790.290 2767.710 791.470 ;
        RECT 2764.930 611.890 2766.110 613.070 ;
        RECT 2766.530 611.890 2767.710 613.070 ;
        RECT 2764.930 610.290 2766.110 611.470 ;
        RECT 2766.530 610.290 2767.710 611.470 ;
        RECT 2764.930 431.890 2766.110 433.070 ;
        RECT 2766.530 431.890 2767.710 433.070 ;
        RECT 2764.930 430.290 2766.110 431.470 ;
        RECT 2766.530 430.290 2767.710 431.470 ;
        RECT 2764.930 251.890 2766.110 253.070 ;
        RECT 2766.530 251.890 2767.710 253.070 ;
        RECT 2764.930 250.290 2766.110 251.470 ;
        RECT 2766.530 250.290 2767.710 251.470 ;
        RECT 2764.930 71.890 2766.110 73.070 ;
        RECT 2766.530 71.890 2767.710 73.070 ;
        RECT 2764.930 70.290 2766.110 71.470 ;
        RECT 2766.530 70.290 2767.710 71.470 ;
        RECT 2764.930 -31.710 2766.110 -30.530 ;
        RECT 2766.530 -31.710 2767.710 -30.530 ;
        RECT 2764.930 -33.310 2766.110 -32.130 ;
        RECT 2766.530 -33.310 2767.710 -32.130 ;
        RECT 2955.510 3551.810 2956.690 3552.990 ;
        RECT 2957.110 3551.810 2958.290 3552.990 ;
        RECT 2955.510 3550.210 2956.690 3551.390 ;
        RECT 2957.110 3550.210 2958.290 3551.390 ;
        RECT 2955.510 3491.890 2956.690 3493.070 ;
        RECT 2957.110 3491.890 2958.290 3493.070 ;
        RECT 2955.510 3490.290 2956.690 3491.470 ;
        RECT 2957.110 3490.290 2958.290 3491.470 ;
        RECT 2955.510 3311.890 2956.690 3313.070 ;
        RECT 2957.110 3311.890 2958.290 3313.070 ;
        RECT 2955.510 3310.290 2956.690 3311.470 ;
        RECT 2957.110 3310.290 2958.290 3311.470 ;
        RECT 2955.510 3131.890 2956.690 3133.070 ;
        RECT 2957.110 3131.890 2958.290 3133.070 ;
        RECT 2955.510 3130.290 2956.690 3131.470 ;
        RECT 2957.110 3130.290 2958.290 3131.470 ;
        RECT 2955.510 2951.890 2956.690 2953.070 ;
        RECT 2957.110 2951.890 2958.290 2953.070 ;
        RECT 2955.510 2950.290 2956.690 2951.470 ;
        RECT 2957.110 2950.290 2958.290 2951.470 ;
        RECT 2955.510 2771.890 2956.690 2773.070 ;
        RECT 2957.110 2771.890 2958.290 2773.070 ;
        RECT 2955.510 2770.290 2956.690 2771.470 ;
        RECT 2957.110 2770.290 2958.290 2771.470 ;
        RECT 2955.510 2591.890 2956.690 2593.070 ;
        RECT 2957.110 2591.890 2958.290 2593.070 ;
        RECT 2955.510 2590.290 2956.690 2591.470 ;
        RECT 2957.110 2590.290 2958.290 2591.470 ;
        RECT 2955.510 2411.890 2956.690 2413.070 ;
        RECT 2957.110 2411.890 2958.290 2413.070 ;
        RECT 2955.510 2410.290 2956.690 2411.470 ;
        RECT 2957.110 2410.290 2958.290 2411.470 ;
        RECT 2955.510 2231.890 2956.690 2233.070 ;
        RECT 2957.110 2231.890 2958.290 2233.070 ;
        RECT 2955.510 2230.290 2956.690 2231.470 ;
        RECT 2957.110 2230.290 2958.290 2231.470 ;
        RECT 2955.510 2051.890 2956.690 2053.070 ;
        RECT 2957.110 2051.890 2958.290 2053.070 ;
        RECT 2955.510 2050.290 2956.690 2051.470 ;
        RECT 2957.110 2050.290 2958.290 2051.470 ;
        RECT 2955.510 1871.890 2956.690 1873.070 ;
        RECT 2957.110 1871.890 2958.290 1873.070 ;
        RECT 2955.510 1870.290 2956.690 1871.470 ;
        RECT 2957.110 1870.290 2958.290 1871.470 ;
        RECT 2955.510 1691.890 2956.690 1693.070 ;
        RECT 2957.110 1691.890 2958.290 1693.070 ;
        RECT 2955.510 1690.290 2956.690 1691.470 ;
        RECT 2957.110 1690.290 2958.290 1691.470 ;
        RECT 2955.510 1511.890 2956.690 1513.070 ;
        RECT 2957.110 1511.890 2958.290 1513.070 ;
        RECT 2955.510 1510.290 2956.690 1511.470 ;
        RECT 2957.110 1510.290 2958.290 1511.470 ;
        RECT 2955.510 1331.890 2956.690 1333.070 ;
        RECT 2957.110 1331.890 2958.290 1333.070 ;
        RECT 2955.510 1330.290 2956.690 1331.470 ;
        RECT 2957.110 1330.290 2958.290 1331.470 ;
        RECT 2955.510 1151.890 2956.690 1153.070 ;
        RECT 2957.110 1151.890 2958.290 1153.070 ;
        RECT 2955.510 1150.290 2956.690 1151.470 ;
        RECT 2957.110 1150.290 2958.290 1151.470 ;
        RECT 2955.510 971.890 2956.690 973.070 ;
        RECT 2957.110 971.890 2958.290 973.070 ;
        RECT 2955.510 970.290 2956.690 971.470 ;
        RECT 2957.110 970.290 2958.290 971.470 ;
        RECT 2955.510 791.890 2956.690 793.070 ;
        RECT 2957.110 791.890 2958.290 793.070 ;
        RECT 2955.510 790.290 2956.690 791.470 ;
        RECT 2957.110 790.290 2958.290 791.470 ;
        RECT 2955.510 611.890 2956.690 613.070 ;
        RECT 2957.110 611.890 2958.290 613.070 ;
        RECT 2955.510 610.290 2956.690 611.470 ;
        RECT 2957.110 610.290 2958.290 611.470 ;
        RECT 2955.510 431.890 2956.690 433.070 ;
        RECT 2957.110 431.890 2958.290 433.070 ;
        RECT 2955.510 430.290 2956.690 431.470 ;
        RECT 2957.110 430.290 2958.290 431.470 ;
        RECT 2955.510 251.890 2956.690 253.070 ;
        RECT 2957.110 251.890 2958.290 253.070 ;
        RECT 2955.510 250.290 2956.690 251.470 ;
        RECT 2957.110 250.290 2958.290 251.470 ;
        RECT 2955.510 71.890 2956.690 73.070 ;
        RECT 2957.110 71.890 2958.290 73.070 ;
        RECT 2955.510 70.290 2956.690 71.470 ;
        RECT 2957.110 70.290 2958.290 71.470 ;
        RECT 2955.510 -31.710 2956.690 -30.530 ;
        RECT 2957.110 -31.710 2958.290 -30.530 ;
        RECT 2955.510 -33.310 2956.690 -32.130 ;
        RECT 2957.110 -33.310 2958.290 -32.130 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
        RECT -43.630 970.130 2963.250 973.230 ;
        RECT -43.630 790.130 2963.250 793.230 ;
        RECT -43.630 610.130 2963.250 613.230 ;
        RECT -43.630 430.130 2963.250 433.230 ;
        RECT -43.630 250.130 2963.250 253.230 ;
        RECT -43.630 70.130 2963.250 73.230 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
        RECT 316.170 1010.000 319.270 3548.350 ;
        RECT 496.170 1010.000 499.270 3548.350 ;
        RECT 676.170 1010.000 679.270 3548.350 ;
        RECT 856.170 1010.000 859.270 3548.350 ;
        RECT 1036.170 1010.000 1039.270 3548.350 ;
        RECT 316.170 -28.670 319.270 390.000 ;
        RECT 496.170 -28.670 499.270 390.000 ;
        RECT 676.170 -28.670 679.270 390.000 ;
        RECT 856.170 -28.670 859.270 390.000 ;
        RECT 1036.170 -28.670 1039.270 390.000 ;
        RECT 1216.170 -28.670 1219.270 3548.350 ;
        RECT 1396.170 -28.670 1399.270 3548.350 ;
        RECT 1576.170 -28.670 1579.270 3548.350 ;
        RECT 1756.170 -28.670 1759.270 3548.350 ;
        RECT 1936.170 -28.670 1939.270 3548.350 ;
        RECT 2116.170 -28.670 2119.270 3548.350 ;
        RECT 2296.170 -28.670 2299.270 3548.350 ;
        RECT 2476.170 -28.670 2479.270 3548.350 ;
        RECT 2656.170 -28.670 2659.270 3548.350 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER via4 ;
        RECT -33.870 3547.010 -32.690 3548.190 ;
        RECT -32.270 3547.010 -31.090 3548.190 ;
        RECT -33.870 3545.410 -32.690 3546.590 ;
        RECT -32.270 3545.410 -31.090 3546.590 ;
        RECT -33.870 3383.290 -32.690 3384.470 ;
        RECT -32.270 3383.290 -31.090 3384.470 ;
        RECT -33.870 3381.690 -32.690 3382.870 ;
        RECT -32.270 3381.690 -31.090 3382.870 ;
        RECT -33.870 3203.290 -32.690 3204.470 ;
        RECT -32.270 3203.290 -31.090 3204.470 ;
        RECT -33.870 3201.690 -32.690 3202.870 ;
        RECT -32.270 3201.690 -31.090 3202.870 ;
        RECT -33.870 3023.290 -32.690 3024.470 ;
        RECT -32.270 3023.290 -31.090 3024.470 ;
        RECT -33.870 3021.690 -32.690 3022.870 ;
        RECT -32.270 3021.690 -31.090 3022.870 ;
        RECT -33.870 2843.290 -32.690 2844.470 ;
        RECT -32.270 2843.290 -31.090 2844.470 ;
        RECT -33.870 2841.690 -32.690 2842.870 ;
        RECT -32.270 2841.690 -31.090 2842.870 ;
        RECT -33.870 2663.290 -32.690 2664.470 ;
        RECT -32.270 2663.290 -31.090 2664.470 ;
        RECT -33.870 2661.690 -32.690 2662.870 ;
        RECT -32.270 2661.690 -31.090 2662.870 ;
        RECT -33.870 2483.290 -32.690 2484.470 ;
        RECT -32.270 2483.290 -31.090 2484.470 ;
        RECT -33.870 2481.690 -32.690 2482.870 ;
        RECT -32.270 2481.690 -31.090 2482.870 ;
        RECT -33.870 2303.290 -32.690 2304.470 ;
        RECT -32.270 2303.290 -31.090 2304.470 ;
        RECT -33.870 2301.690 -32.690 2302.870 ;
        RECT -32.270 2301.690 -31.090 2302.870 ;
        RECT -33.870 2123.290 -32.690 2124.470 ;
        RECT -32.270 2123.290 -31.090 2124.470 ;
        RECT -33.870 2121.690 -32.690 2122.870 ;
        RECT -32.270 2121.690 -31.090 2122.870 ;
        RECT -33.870 1943.290 -32.690 1944.470 ;
        RECT -32.270 1943.290 -31.090 1944.470 ;
        RECT -33.870 1941.690 -32.690 1942.870 ;
        RECT -32.270 1941.690 -31.090 1942.870 ;
        RECT -33.870 1763.290 -32.690 1764.470 ;
        RECT -32.270 1763.290 -31.090 1764.470 ;
        RECT -33.870 1761.690 -32.690 1762.870 ;
        RECT -32.270 1761.690 -31.090 1762.870 ;
        RECT -33.870 1583.290 -32.690 1584.470 ;
        RECT -32.270 1583.290 -31.090 1584.470 ;
        RECT -33.870 1581.690 -32.690 1582.870 ;
        RECT -32.270 1581.690 -31.090 1582.870 ;
        RECT -33.870 1403.290 -32.690 1404.470 ;
        RECT -32.270 1403.290 -31.090 1404.470 ;
        RECT -33.870 1401.690 -32.690 1402.870 ;
        RECT -32.270 1401.690 -31.090 1402.870 ;
        RECT -33.870 1223.290 -32.690 1224.470 ;
        RECT -32.270 1223.290 -31.090 1224.470 ;
        RECT -33.870 1221.690 -32.690 1222.870 ;
        RECT -32.270 1221.690 -31.090 1222.870 ;
        RECT -33.870 1043.290 -32.690 1044.470 ;
        RECT -32.270 1043.290 -31.090 1044.470 ;
        RECT -33.870 1041.690 -32.690 1042.870 ;
        RECT -32.270 1041.690 -31.090 1042.870 ;
        RECT -33.870 863.290 -32.690 864.470 ;
        RECT -32.270 863.290 -31.090 864.470 ;
        RECT -33.870 861.690 -32.690 862.870 ;
        RECT -32.270 861.690 -31.090 862.870 ;
        RECT -33.870 683.290 -32.690 684.470 ;
        RECT -32.270 683.290 -31.090 684.470 ;
        RECT -33.870 681.690 -32.690 682.870 ;
        RECT -32.270 681.690 -31.090 682.870 ;
        RECT -33.870 503.290 -32.690 504.470 ;
        RECT -32.270 503.290 -31.090 504.470 ;
        RECT -33.870 501.690 -32.690 502.870 ;
        RECT -32.270 501.690 -31.090 502.870 ;
        RECT -33.870 323.290 -32.690 324.470 ;
        RECT -32.270 323.290 -31.090 324.470 ;
        RECT -33.870 321.690 -32.690 322.870 ;
        RECT -32.270 321.690 -31.090 322.870 ;
        RECT -33.870 143.290 -32.690 144.470 ;
        RECT -32.270 143.290 -31.090 144.470 ;
        RECT -33.870 141.690 -32.690 142.870 ;
        RECT -32.270 141.690 -31.090 142.870 ;
        RECT -33.870 -26.910 -32.690 -25.730 ;
        RECT -32.270 -26.910 -31.090 -25.730 ;
        RECT -33.870 -28.510 -32.690 -27.330 ;
        RECT -32.270 -28.510 -31.090 -27.330 ;
        RECT 136.330 3547.010 137.510 3548.190 ;
        RECT 137.930 3547.010 139.110 3548.190 ;
        RECT 136.330 3545.410 137.510 3546.590 ;
        RECT 137.930 3545.410 139.110 3546.590 ;
        RECT 136.330 3383.290 137.510 3384.470 ;
        RECT 137.930 3383.290 139.110 3384.470 ;
        RECT 136.330 3381.690 137.510 3382.870 ;
        RECT 137.930 3381.690 139.110 3382.870 ;
        RECT 136.330 3203.290 137.510 3204.470 ;
        RECT 137.930 3203.290 139.110 3204.470 ;
        RECT 136.330 3201.690 137.510 3202.870 ;
        RECT 137.930 3201.690 139.110 3202.870 ;
        RECT 136.330 3023.290 137.510 3024.470 ;
        RECT 137.930 3023.290 139.110 3024.470 ;
        RECT 136.330 3021.690 137.510 3022.870 ;
        RECT 137.930 3021.690 139.110 3022.870 ;
        RECT 136.330 2843.290 137.510 2844.470 ;
        RECT 137.930 2843.290 139.110 2844.470 ;
        RECT 136.330 2841.690 137.510 2842.870 ;
        RECT 137.930 2841.690 139.110 2842.870 ;
        RECT 136.330 2663.290 137.510 2664.470 ;
        RECT 137.930 2663.290 139.110 2664.470 ;
        RECT 136.330 2661.690 137.510 2662.870 ;
        RECT 137.930 2661.690 139.110 2662.870 ;
        RECT 136.330 2483.290 137.510 2484.470 ;
        RECT 137.930 2483.290 139.110 2484.470 ;
        RECT 136.330 2481.690 137.510 2482.870 ;
        RECT 137.930 2481.690 139.110 2482.870 ;
        RECT 136.330 2303.290 137.510 2304.470 ;
        RECT 137.930 2303.290 139.110 2304.470 ;
        RECT 136.330 2301.690 137.510 2302.870 ;
        RECT 137.930 2301.690 139.110 2302.870 ;
        RECT 136.330 2123.290 137.510 2124.470 ;
        RECT 137.930 2123.290 139.110 2124.470 ;
        RECT 136.330 2121.690 137.510 2122.870 ;
        RECT 137.930 2121.690 139.110 2122.870 ;
        RECT 136.330 1943.290 137.510 1944.470 ;
        RECT 137.930 1943.290 139.110 1944.470 ;
        RECT 136.330 1941.690 137.510 1942.870 ;
        RECT 137.930 1941.690 139.110 1942.870 ;
        RECT 136.330 1763.290 137.510 1764.470 ;
        RECT 137.930 1763.290 139.110 1764.470 ;
        RECT 136.330 1761.690 137.510 1762.870 ;
        RECT 137.930 1761.690 139.110 1762.870 ;
        RECT 136.330 1583.290 137.510 1584.470 ;
        RECT 137.930 1583.290 139.110 1584.470 ;
        RECT 136.330 1581.690 137.510 1582.870 ;
        RECT 137.930 1581.690 139.110 1582.870 ;
        RECT 136.330 1403.290 137.510 1404.470 ;
        RECT 137.930 1403.290 139.110 1404.470 ;
        RECT 136.330 1401.690 137.510 1402.870 ;
        RECT 137.930 1401.690 139.110 1402.870 ;
        RECT 136.330 1223.290 137.510 1224.470 ;
        RECT 137.930 1223.290 139.110 1224.470 ;
        RECT 136.330 1221.690 137.510 1222.870 ;
        RECT 137.930 1221.690 139.110 1222.870 ;
        RECT 136.330 1043.290 137.510 1044.470 ;
        RECT 137.930 1043.290 139.110 1044.470 ;
        RECT 136.330 1041.690 137.510 1042.870 ;
        RECT 137.930 1041.690 139.110 1042.870 ;
        RECT 316.330 3547.010 317.510 3548.190 ;
        RECT 317.930 3547.010 319.110 3548.190 ;
        RECT 316.330 3545.410 317.510 3546.590 ;
        RECT 317.930 3545.410 319.110 3546.590 ;
        RECT 316.330 3383.290 317.510 3384.470 ;
        RECT 317.930 3383.290 319.110 3384.470 ;
        RECT 316.330 3381.690 317.510 3382.870 ;
        RECT 317.930 3381.690 319.110 3382.870 ;
        RECT 316.330 3203.290 317.510 3204.470 ;
        RECT 317.930 3203.290 319.110 3204.470 ;
        RECT 316.330 3201.690 317.510 3202.870 ;
        RECT 317.930 3201.690 319.110 3202.870 ;
        RECT 316.330 3023.290 317.510 3024.470 ;
        RECT 317.930 3023.290 319.110 3024.470 ;
        RECT 316.330 3021.690 317.510 3022.870 ;
        RECT 317.930 3021.690 319.110 3022.870 ;
        RECT 316.330 2843.290 317.510 2844.470 ;
        RECT 317.930 2843.290 319.110 2844.470 ;
        RECT 316.330 2841.690 317.510 2842.870 ;
        RECT 317.930 2841.690 319.110 2842.870 ;
        RECT 316.330 2663.290 317.510 2664.470 ;
        RECT 317.930 2663.290 319.110 2664.470 ;
        RECT 316.330 2661.690 317.510 2662.870 ;
        RECT 317.930 2661.690 319.110 2662.870 ;
        RECT 316.330 2483.290 317.510 2484.470 ;
        RECT 317.930 2483.290 319.110 2484.470 ;
        RECT 316.330 2481.690 317.510 2482.870 ;
        RECT 317.930 2481.690 319.110 2482.870 ;
        RECT 316.330 2303.290 317.510 2304.470 ;
        RECT 317.930 2303.290 319.110 2304.470 ;
        RECT 316.330 2301.690 317.510 2302.870 ;
        RECT 317.930 2301.690 319.110 2302.870 ;
        RECT 316.330 2123.290 317.510 2124.470 ;
        RECT 317.930 2123.290 319.110 2124.470 ;
        RECT 316.330 2121.690 317.510 2122.870 ;
        RECT 317.930 2121.690 319.110 2122.870 ;
        RECT 316.330 1943.290 317.510 1944.470 ;
        RECT 317.930 1943.290 319.110 1944.470 ;
        RECT 316.330 1941.690 317.510 1942.870 ;
        RECT 317.930 1941.690 319.110 1942.870 ;
        RECT 316.330 1763.290 317.510 1764.470 ;
        RECT 317.930 1763.290 319.110 1764.470 ;
        RECT 316.330 1761.690 317.510 1762.870 ;
        RECT 317.930 1761.690 319.110 1762.870 ;
        RECT 316.330 1583.290 317.510 1584.470 ;
        RECT 317.930 1583.290 319.110 1584.470 ;
        RECT 316.330 1581.690 317.510 1582.870 ;
        RECT 317.930 1581.690 319.110 1582.870 ;
        RECT 316.330 1403.290 317.510 1404.470 ;
        RECT 317.930 1403.290 319.110 1404.470 ;
        RECT 316.330 1401.690 317.510 1402.870 ;
        RECT 317.930 1401.690 319.110 1402.870 ;
        RECT 316.330 1223.290 317.510 1224.470 ;
        RECT 317.930 1223.290 319.110 1224.470 ;
        RECT 316.330 1221.690 317.510 1222.870 ;
        RECT 317.930 1221.690 319.110 1222.870 ;
        RECT 316.330 1043.290 317.510 1044.470 ;
        RECT 317.930 1043.290 319.110 1044.470 ;
        RECT 316.330 1041.690 317.510 1042.870 ;
        RECT 317.930 1041.690 319.110 1042.870 ;
        RECT 496.330 3547.010 497.510 3548.190 ;
        RECT 497.930 3547.010 499.110 3548.190 ;
        RECT 496.330 3545.410 497.510 3546.590 ;
        RECT 497.930 3545.410 499.110 3546.590 ;
        RECT 496.330 3383.290 497.510 3384.470 ;
        RECT 497.930 3383.290 499.110 3384.470 ;
        RECT 496.330 3381.690 497.510 3382.870 ;
        RECT 497.930 3381.690 499.110 3382.870 ;
        RECT 496.330 3203.290 497.510 3204.470 ;
        RECT 497.930 3203.290 499.110 3204.470 ;
        RECT 496.330 3201.690 497.510 3202.870 ;
        RECT 497.930 3201.690 499.110 3202.870 ;
        RECT 496.330 3023.290 497.510 3024.470 ;
        RECT 497.930 3023.290 499.110 3024.470 ;
        RECT 496.330 3021.690 497.510 3022.870 ;
        RECT 497.930 3021.690 499.110 3022.870 ;
        RECT 496.330 2843.290 497.510 2844.470 ;
        RECT 497.930 2843.290 499.110 2844.470 ;
        RECT 496.330 2841.690 497.510 2842.870 ;
        RECT 497.930 2841.690 499.110 2842.870 ;
        RECT 496.330 2663.290 497.510 2664.470 ;
        RECT 497.930 2663.290 499.110 2664.470 ;
        RECT 496.330 2661.690 497.510 2662.870 ;
        RECT 497.930 2661.690 499.110 2662.870 ;
        RECT 496.330 2483.290 497.510 2484.470 ;
        RECT 497.930 2483.290 499.110 2484.470 ;
        RECT 496.330 2481.690 497.510 2482.870 ;
        RECT 497.930 2481.690 499.110 2482.870 ;
        RECT 496.330 2303.290 497.510 2304.470 ;
        RECT 497.930 2303.290 499.110 2304.470 ;
        RECT 496.330 2301.690 497.510 2302.870 ;
        RECT 497.930 2301.690 499.110 2302.870 ;
        RECT 496.330 2123.290 497.510 2124.470 ;
        RECT 497.930 2123.290 499.110 2124.470 ;
        RECT 496.330 2121.690 497.510 2122.870 ;
        RECT 497.930 2121.690 499.110 2122.870 ;
        RECT 496.330 1943.290 497.510 1944.470 ;
        RECT 497.930 1943.290 499.110 1944.470 ;
        RECT 496.330 1941.690 497.510 1942.870 ;
        RECT 497.930 1941.690 499.110 1942.870 ;
        RECT 496.330 1763.290 497.510 1764.470 ;
        RECT 497.930 1763.290 499.110 1764.470 ;
        RECT 496.330 1761.690 497.510 1762.870 ;
        RECT 497.930 1761.690 499.110 1762.870 ;
        RECT 496.330 1583.290 497.510 1584.470 ;
        RECT 497.930 1583.290 499.110 1584.470 ;
        RECT 496.330 1581.690 497.510 1582.870 ;
        RECT 497.930 1581.690 499.110 1582.870 ;
        RECT 496.330 1403.290 497.510 1404.470 ;
        RECT 497.930 1403.290 499.110 1404.470 ;
        RECT 496.330 1401.690 497.510 1402.870 ;
        RECT 497.930 1401.690 499.110 1402.870 ;
        RECT 496.330 1223.290 497.510 1224.470 ;
        RECT 497.930 1223.290 499.110 1224.470 ;
        RECT 496.330 1221.690 497.510 1222.870 ;
        RECT 497.930 1221.690 499.110 1222.870 ;
        RECT 496.330 1043.290 497.510 1044.470 ;
        RECT 497.930 1043.290 499.110 1044.470 ;
        RECT 496.330 1041.690 497.510 1042.870 ;
        RECT 497.930 1041.690 499.110 1042.870 ;
        RECT 676.330 3547.010 677.510 3548.190 ;
        RECT 677.930 3547.010 679.110 3548.190 ;
        RECT 676.330 3545.410 677.510 3546.590 ;
        RECT 677.930 3545.410 679.110 3546.590 ;
        RECT 676.330 3383.290 677.510 3384.470 ;
        RECT 677.930 3383.290 679.110 3384.470 ;
        RECT 676.330 3381.690 677.510 3382.870 ;
        RECT 677.930 3381.690 679.110 3382.870 ;
        RECT 676.330 3203.290 677.510 3204.470 ;
        RECT 677.930 3203.290 679.110 3204.470 ;
        RECT 676.330 3201.690 677.510 3202.870 ;
        RECT 677.930 3201.690 679.110 3202.870 ;
        RECT 676.330 3023.290 677.510 3024.470 ;
        RECT 677.930 3023.290 679.110 3024.470 ;
        RECT 676.330 3021.690 677.510 3022.870 ;
        RECT 677.930 3021.690 679.110 3022.870 ;
        RECT 676.330 2843.290 677.510 2844.470 ;
        RECT 677.930 2843.290 679.110 2844.470 ;
        RECT 676.330 2841.690 677.510 2842.870 ;
        RECT 677.930 2841.690 679.110 2842.870 ;
        RECT 676.330 2663.290 677.510 2664.470 ;
        RECT 677.930 2663.290 679.110 2664.470 ;
        RECT 676.330 2661.690 677.510 2662.870 ;
        RECT 677.930 2661.690 679.110 2662.870 ;
        RECT 676.330 2483.290 677.510 2484.470 ;
        RECT 677.930 2483.290 679.110 2484.470 ;
        RECT 676.330 2481.690 677.510 2482.870 ;
        RECT 677.930 2481.690 679.110 2482.870 ;
        RECT 676.330 2303.290 677.510 2304.470 ;
        RECT 677.930 2303.290 679.110 2304.470 ;
        RECT 676.330 2301.690 677.510 2302.870 ;
        RECT 677.930 2301.690 679.110 2302.870 ;
        RECT 676.330 2123.290 677.510 2124.470 ;
        RECT 677.930 2123.290 679.110 2124.470 ;
        RECT 676.330 2121.690 677.510 2122.870 ;
        RECT 677.930 2121.690 679.110 2122.870 ;
        RECT 676.330 1943.290 677.510 1944.470 ;
        RECT 677.930 1943.290 679.110 1944.470 ;
        RECT 676.330 1941.690 677.510 1942.870 ;
        RECT 677.930 1941.690 679.110 1942.870 ;
        RECT 676.330 1763.290 677.510 1764.470 ;
        RECT 677.930 1763.290 679.110 1764.470 ;
        RECT 676.330 1761.690 677.510 1762.870 ;
        RECT 677.930 1761.690 679.110 1762.870 ;
        RECT 676.330 1583.290 677.510 1584.470 ;
        RECT 677.930 1583.290 679.110 1584.470 ;
        RECT 676.330 1581.690 677.510 1582.870 ;
        RECT 677.930 1581.690 679.110 1582.870 ;
        RECT 676.330 1403.290 677.510 1404.470 ;
        RECT 677.930 1403.290 679.110 1404.470 ;
        RECT 676.330 1401.690 677.510 1402.870 ;
        RECT 677.930 1401.690 679.110 1402.870 ;
        RECT 676.330 1223.290 677.510 1224.470 ;
        RECT 677.930 1223.290 679.110 1224.470 ;
        RECT 676.330 1221.690 677.510 1222.870 ;
        RECT 677.930 1221.690 679.110 1222.870 ;
        RECT 676.330 1043.290 677.510 1044.470 ;
        RECT 677.930 1043.290 679.110 1044.470 ;
        RECT 676.330 1041.690 677.510 1042.870 ;
        RECT 677.930 1041.690 679.110 1042.870 ;
        RECT 856.330 3547.010 857.510 3548.190 ;
        RECT 857.930 3547.010 859.110 3548.190 ;
        RECT 856.330 3545.410 857.510 3546.590 ;
        RECT 857.930 3545.410 859.110 3546.590 ;
        RECT 856.330 3383.290 857.510 3384.470 ;
        RECT 857.930 3383.290 859.110 3384.470 ;
        RECT 856.330 3381.690 857.510 3382.870 ;
        RECT 857.930 3381.690 859.110 3382.870 ;
        RECT 856.330 3203.290 857.510 3204.470 ;
        RECT 857.930 3203.290 859.110 3204.470 ;
        RECT 856.330 3201.690 857.510 3202.870 ;
        RECT 857.930 3201.690 859.110 3202.870 ;
        RECT 856.330 3023.290 857.510 3024.470 ;
        RECT 857.930 3023.290 859.110 3024.470 ;
        RECT 856.330 3021.690 857.510 3022.870 ;
        RECT 857.930 3021.690 859.110 3022.870 ;
        RECT 856.330 2843.290 857.510 2844.470 ;
        RECT 857.930 2843.290 859.110 2844.470 ;
        RECT 856.330 2841.690 857.510 2842.870 ;
        RECT 857.930 2841.690 859.110 2842.870 ;
        RECT 856.330 2663.290 857.510 2664.470 ;
        RECT 857.930 2663.290 859.110 2664.470 ;
        RECT 856.330 2661.690 857.510 2662.870 ;
        RECT 857.930 2661.690 859.110 2662.870 ;
        RECT 856.330 2483.290 857.510 2484.470 ;
        RECT 857.930 2483.290 859.110 2484.470 ;
        RECT 856.330 2481.690 857.510 2482.870 ;
        RECT 857.930 2481.690 859.110 2482.870 ;
        RECT 856.330 2303.290 857.510 2304.470 ;
        RECT 857.930 2303.290 859.110 2304.470 ;
        RECT 856.330 2301.690 857.510 2302.870 ;
        RECT 857.930 2301.690 859.110 2302.870 ;
        RECT 856.330 2123.290 857.510 2124.470 ;
        RECT 857.930 2123.290 859.110 2124.470 ;
        RECT 856.330 2121.690 857.510 2122.870 ;
        RECT 857.930 2121.690 859.110 2122.870 ;
        RECT 856.330 1943.290 857.510 1944.470 ;
        RECT 857.930 1943.290 859.110 1944.470 ;
        RECT 856.330 1941.690 857.510 1942.870 ;
        RECT 857.930 1941.690 859.110 1942.870 ;
        RECT 856.330 1763.290 857.510 1764.470 ;
        RECT 857.930 1763.290 859.110 1764.470 ;
        RECT 856.330 1761.690 857.510 1762.870 ;
        RECT 857.930 1761.690 859.110 1762.870 ;
        RECT 856.330 1583.290 857.510 1584.470 ;
        RECT 857.930 1583.290 859.110 1584.470 ;
        RECT 856.330 1581.690 857.510 1582.870 ;
        RECT 857.930 1581.690 859.110 1582.870 ;
        RECT 856.330 1403.290 857.510 1404.470 ;
        RECT 857.930 1403.290 859.110 1404.470 ;
        RECT 856.330 1401.690 857.510 1402.870 ;
        RECT 857.930 1401.690 859.110 1402.870 ;
        RECT 856.330 1223.290 857.510 1224.470 ;
        RECT 857.930 1223.290 859.110 1224.470 ;
        RECT 856.330 1221.690 857.510 1222.870 ;
        RECT 857.930 1221.690 859.110 1222.870 ;
        RECT 856.330 1043.290 857.510 1044.470 ;
        RECT 857.930 1043.290 859.110 1044.470 ;
        RECT 856.330 1041.690 857.510 1042.870 ;
        RECT 857.930 1041.690 859.110 1042.870 ;
        RECT 1036.330 3547.010 1037.510 3548.190 ;
        RECT 1037.930 3547.010 1039.110 3548.190 ;
        RECT 1036.330 3545.410 1037.510 3546.590 ;
        RECT 1037.930 3545.410 1039.110 3546.590 ;
        RECT 1036.330 3383.290 1037.510 3384.470 ;
        RECT 1037.930 3383.290 1039.110 3384.470 ;
        RECT 1036.330 3381.690 1037.510 3382.870 ;
        RECT 1037.930 3381.690 1039.110 3382.870 ;
        RECT 1036.330 3203.290 1037.510 3204.470 ;
        RECT 1037.930 3203.290 1039.110 3204.470 ;
        RECT 1036.330 3201.690 1037.510 3202.870 ;
        RECT 1037.930 3201.690 1039.110 3202.870 ;
        RECT 1036.330 3023.290 1037.510 3024.470 ;
        RECT 1037.930 3023.290 1039.110 3024.470 ;
        RECT 1036.330 3021.690 1037.510 3022.870 ;
        RECT 1037.930 3021.690 1039.110 3022.870 ;
        RECT 1036.330 2843.290 1037.510 2844.470 ;
        RECT 1037.930 2843.290 1039.110 2844.470 ;
        RECT 1036.330 2841.690 1037.510 2842.870 ;
        RECT 1037.930 2841.690 1039.110 2842.870 ;
        RECT 1036.330 2663.290 1037.510 2664.470 ;
        RECT 1037.930 2663.290 1039.110 2664.470 ;
        RECT 1036.330 2661.690 1037.510 2662.870 ;
        RECT 1037.930 2661.690 1039.110 2662.870 ;
        RECT 1036.330 2483.290 1037.510 2484.470 ;
        RECT 1037.930 2483.290 1039.110 2484.470 ;
        RECT 1036.330 2481.690 1037.510 2482.870 ;
        RECT 1037.930 2481.690 1039.110 2482.870 ;
        RECT 1036.330 2303.290 1037.510 2304.470 ;
        RECT 1037.930 2303.290 1039.110 2304.470 ;
        RECT 1036.330 2301.690 1037.510 2302.870 ;
        RECT 1037.930 2301.690 1039.110 2302.870 ;
        RECT 1036.330 2123.290 1037.510 2124.470 ;
        RECT 1037.930 2123.290 1039.110 2124.470 ;
        RECT 1036.330 2121.690 1037.510 2122.870 ;
        RECT 1037.930 2121.690 1039.110 2122.870 ;
        RECT 1036.330 1943.290 1037.510 1944.470 ;
        RECT 1037.930 1943.290 1039.110 1944.470 ;
        RECT 1036.330 1941.690 1037.510 1942.870 ;
        RECT 1037.930 1941.690 1039.110 1942.870 ;
        RECT 1036.330 1763.290 1037.510 1764.470 ;
        RECT 1037.930 1763.290 1039.110 1764.470 ;
        RECT 1036.330 1761.690 1037.510 1762.870 ;
        RECT 1037.930 1761.690 1039.110 1762.870 ;
        RECT 1036.330 1583.290 1037.510 1584.470 ;
        RECT 1037.930 1583.290 1039.110 1584.470 ;
        RECT 1036.330 1581.690 1037.510 1582.870 ;
        RECT 1037.930 1581.690 1039.110 1582.870 ;
        RECT 1036.330 1403.290 1037.510 1404.470 ;
        RECT 1037.930 1403.290 1039.110 1404.470 ;
        RECT 1036.330 1401.690 1037.510 1402.870 ;
        RECT 1037.930 1401.690 1039.110 1402.870 ;
        RECT 1036.330 1223.290 1037.510 1224.470 ;
        RECT 1037.930 1223.290 1039.110 1224.470 ;
        RECT 1036.330 1221.690 1037.510 1222.870 ;
        RECT 1037.930 1221.690 1039.110 1222.870 ;
        RECT 1036.330 1043.290 1037.510 1044.470 ;
        RECT 1037.930 1043.290 1039.110 1044.470 ;
        RECT 1036.330 1041.690 1037.510 1042.870 ;
        RECT 1037.930 1041.690 1039.110 1042.870 ;
        RECT 1216.330 3547.010 1217.510 3548.190 ;
        RECT 1217.930 3547.010 1219.110 3548.190 ;
        RECT 1216.330 3545.410 1217.510 3546.590 ;
        RECT 1217.930 3545.410 1219.110 3546.590 ;
        RECT 1216.330 3383.290 1217.510 3384.470 ;
        RECT 1217.930 3383.290 1219.110 3384.470 ;
        RECT 1216.330 3381.690 1217.510 3382.870 ;
        RECT 1217.930 3381.690 1219.110 3382.870 ;
        RECT 1216.330 3203.290 1217.510 3204.470 ;
        RECT 1217.930 3203.290 1219.110 3204.470 ;
        RECT 1216.330 3201.690 1217.510 3202.870 ;
        RECT 1217.930 3201.690 1219.110 3202.870 ;
        RECT 1216.330 3023.290 1217.510 3024.470 ;
        RECT 1217.930 3023.290 1219.110 3024.470 ;
        RECT 1216.330 3021.690 1217.510 3022.870 ;
        RECT 1217.930 3021.690 1219.110 3022.870 ;
        RECT 1216.330 2843.290 1217.510 2844.470 ;
        RECT 1217.930 2843.290 1219.110 2844.470 ;
        RECT 1216.330 2841.690 1217.510 2842.870 ;
        RECT 1217.930 2841.690 1219.110 2842.870 ;
        RECT 1216.330 2663.290 1217.510 2664.470 ;
        RECT 1217.930 2663.290 1219.110 2664.470 ;
        RECT 1216.330 2661.690 1217.510 2662.870 ;
        RECT 1217.930 2661.690 1219.110 2662.870 ;
        RECT 1216.330 2483.290 1217.510 2484.470 ;
        RECT 1217.930 2483.290 1219.110 2484.470 ;
        RECT 1216.330 2481.690 1217.510 2482.870 ;
        RECT 1217.930 2481.690 1219.110 2482.870 ;
        RECT 1216.330 2303.290 1217.510 2304.470 ;
        RECT 1217.930 2303.290 1219.110 2304.470 ;
        RECT 1216.330 2301.690 1217.510 2302.870 ;
        RECT 1217.930 2301.690 1219.110 2302.870 ;
        RECT 1216.330 2123.290 1217.510 2124.470 ;
        RECT 1217.930 2123.290 1219.110 2124.470 ;
        RECT 1216.330 2121.690 1217.510 2122.870 ;
        RECT 1217.930 2121.690 1219.110 2122.870 ;
        RECT 1216.330 1943.290 1217.510 1944.470 ;
        RECT 1217.930 1943.290 1219.110 1944.470 ;
        RECT 1216.330 1941.690 1217.510 1942.870 ;
        RECT 1217.930 1941.690 1219.110 1942.870 ;
        RECT 1216.330 1763.290 1217.510 1764.470 ;
        RECT 1217.930 1763.290 1219.110 1764.470 ;
        RECT 1216.330 1761.690 1217.510 1762.870 ;
        RECT 1217.930 1761.690 1219.110 1762.870 ;
        RECT 1216.330 1583.290 1217.510 1584.470 ;
        RECT 1217.930 1583.290 1219.110 1584.470 ;
        RECT 1216.330 1581.690 1217.510 1582.870 ;
        RECT 1217.930 1581.690 1219.110 1582.870 ;
        RECT 1216.330 1403.290 1217.510 1404.470 ;
        RECT 1217.930 1403.290 1219.110 1404.470 ;
        RECT 1216.330 1401.690 1217.510 1402.870 ;
        RECT 1217.930 1401.690 1219.110 1402.870 ;
        RECT 1216.330 1223.290 1217.510 1224.470 ;
        RECT 1217.930 1223.290 1219.110 1224.470 ;
        RECT 1216.330 1221.690 1217.510 1222.870 ;
        RECT 1217.930 1221.690 1219.110 1222.870 ;
        RECT 1216.330 1043.290 1217.510 1044.470 ;
        RECT 1217.930 1043.290 1219.110 1044.470 ;
        RECT 1216.330 1041.690 1217.510 1042.870 ;
        RECT 1217.930 1041.690 1219.110 1042.870 ;
        RECT 136.330 863.290 137.510 864.470 ;
        RECT 137.930 863.290 139.110 864.470 ;
        RECT 136.330 861.690 137.510 862.870 ;
        RECT 137.930 861.690 139.110 862.870 ;
        RECT 136.330 683.290 137.510 684.470 ;
        RECT 137.930 683.290 139.110 684.470 ;
        RECT 136.330 681.690 137.510 682.870 ;
        RECT 137.930 681.690 139.110 682.870 ;
        RECT 136.330 503.290 137.510 504.470 ;
        RECT 137.930 503.290 139.110 504.470 ;
        RECT 136.330 501.690 137.510 502.870 ;
        RECT 137.930 501.690 139.110 502.870 ;
        RECT 1216.330 863.290 1217.510 864.470 ;
        RECT 1217.930 863.290 1219.110 864.470 ;
        RECT 1216.330 861.690 1217.510 862.870 ;
        RECT 1217.930 861.690 1219.110 862.870 ;
        RECT 1216.330 683.290 1217.510 684.470 ;
        RECT 1217.930 683.290 1219.110 684.470 ;
        RECT 1216.330 681.690 1217.510 682.870 ;
        RECT 1217.930 681.690 1219.110 682.870 ;
        RECT 1216.330 503.290 1217.510 504.470 ;
        RECT 1217.930 503.290 1219.110 504.470 ;
        RECT 1216.330 501.690 1217.510 502.870 ;
        RECT 1217.930 501.690 1219.110 502.870 ;
        RECT 136.330 323.290 137.510 324.470 ;
        RECT 137.930 323.290 139.110 324.470 ;
        RECT 136.330 321.690 137.510 322.870 ;
        RECT 137.930 321.690 139.110 322.870 ;
        RECT 136.330 143.290 137.510 144.470 ;
        RECT 137.930 143.290 139.110 144.470 ;
        RECT 136.330 141.690 137.510 142.870 ;
        RECT 137.930 141.690 139.110 142.870 ;
        RECT 136.330 -26.910 137.510 -25.730 ;
        RECT 137.930 -26.910 139.110 -25.730 ;
        RECT 136.330 -28.510 137.510 -27.330 ;
        RECT 137.930 -28.510 139.110 -27.330 ;
        RECT 316.330 323.290 317.510 324.470 ;
        RECT 317.930 323.290 319.110 324.470 ;
        RECT 316.330 321.690 317.510 322.870 ;
        RECT 317.930 321.690 319.110 322.870 ;
        RECT 316.330 143.290 317.510 144.470 ;
        RECT 317.930 143.290 319.110 144.470 ;
        RECT 316.330 141.690 317.510 142.870 ;
        RECT 317.930 141.690 319.110 142.870 ;
        RECT 316.330 -26.910 317.510 -25.730 ;
        RECT 317.930 -26.910 319.110 -25.730 ;
        RECT 316.330 -28.510 317.510 -27.330 ;
        RECT 317.930 -28.510 319.110 -27.330 ;
        RECT 496.330 323.290 497.510 324.470 ;
        RECT 497.930 323.290 499.110 324.470 ;
        RECT 496.330 321.690 497.510 322.870 ;
        RECT 497.930 321.690 499.110 322.870 ;
        RECT 496.330 143.290 497.510 144.470 ;
        RECT 497.930 143.290 499.110 144.470 ;
        RECT 496.330 141.690 497.510 142.870 ;
        RECT 497.930 141.690 499.110 142.870 ;
        RECT 496.330 -26.910 497.510 -25.730 ;
        RECT 497.930 -26.910 499.110 -25.730 ;
        RECT 496.330 -28.510 497.510 -27.330 ;
        RECT 497.930 -28.510 499.110 -27.330 ;
        RECT 676.330 323.290 677.510 324.470 ;
        RECT 677.930 323.290 679.110 324.470 ;
        RECT 676.330 321.690 677.510 322.870 ;
        RECT 677.930 321.690 679.110 322.870 ;
        RECT 676.330 143.290 677.510 144.470 ;
        RECT 677.930 143.290 679.110 144.470 ;
        RECT 676.330 141.690 677.510 142.870 ;
        RECT 677.930 141.690 679.110 142.870 ;
        RECT 676.330 -26.910 677.510 -25.730 ;
        RECT 677.930 -26.910 679.110 -25.730 ;
        RECT 676.330 -28.510 677.510 -27.330 ;
        RECT 677.930 -28.510 679.110 -27.330 ;
        RECT 856.330 323.290 857.510 324.470 ;
        RECT 857.930 323.290 859.110 324.470 ;
        RECT 856.330 321.690 857.510 322.870 ;
        RECT 857.930 321.690 859.110 322.870 ;
        RECT 856.330 143.290 857.510 144.470 ;
        RECT 857.930 143.290 859.110 144.470 ;
        RECT 856.330 141.690 857.510 142.870 ;
        RECT 857.930 141.690 859.110 142.870 ;
        RECT 856.330 -26.910 857.510 -25.730 ;
        RECT 857.930 -26.910 859.110 -25.730 ;
        RECT 856.330 -28.510 857.510 -27.330 ;
        RECT 857.930 -28.510 859.110 -27.330 ;
        RECT 1036.330 323.290 1037.510 324.470 ;
        RECT 1037.930 323.290 1039.110 324.470 ;
        RECT 1036.330 321.690 1037.510 322.870 ;
        RECT 1037.930 321.690 1039.110 322.870 ;
        RECT 1036.330 143.290 1037.510 144.470 ;
        RECT 1037.930 143.290 1039.110 144.470 ;
        RECT 1036.330 141.690 1037.510 142.870 ;
        RECT 1037.930 141.690 1039.110 142.870 ;
        RECT 1036.330 -26.910 1037.510 -25.730 ;
        RECT 1037.930 -26.910 1039.110 -25.730 ;
        RECT 1036.330 -28.510 1037.510 -27.330 ;
        RECT 1037.930 -28.510 1039.110 -27.330 ;
        RECT 1216.330 323.290 1217.510 324.470 ;
        RECT 1217.930 323.290 1219.110 324.470 ;
        RECT 1216.330 321.690 1217.510 322.870 ;
        RECT 1217.930 321.690 1219.110 322.870 ;
        RECT 1216.330 143.290 1217.510 144.470 ;
        RECT 1217.930 143.290 1219.110 144.470 ;
        RECT 1216.330 141.690 1217.510 142.870 ;
        RECT 1217.930 141.690 1219.110 142.870 ;
        RECT 1216.330 -26.910 1217.510 -25.730 ;
        RECT 1217.930 -26.910 1219.110 -25.730 ;
        RECT 1216.330 -28.510 1217.510 -27.330 ;
        RECT 1217.930 -28.510 1219.110 -27.330 ;
        RECT 1396.330 3547.010 1397.510 3548.190 ;
        RECT 1397.930 3547.010 1399.110 3548.190 ;
        RECT 1396.330 3545.410 1397.510 3546.590 ;
        RECT 1397.930 3545.410 1399.110 3546.590 ;
        RECT 1396.330 3383.290 1397.510 3384.470 ;
        RECT 1397.930 3383.290 1399.110 3384.470 ;
        RECT 1396.330 3381.690 1397.510 3382.870 ;
        RECT 1397.930 3381.690 1399.110 3382.870 ;
        RECT 1396.330 3203.290 1397.510 3204.470 ;
        RECT 1397.930 3203.290 1399.110 3204.470 ;
        RECT 1396.330 3201.690 1397.510 3202.870 ;
        RECT 1397.930 3201.690 1399.110 3202.870 ;
        RECT 1396.330 3023.290 1397.510 3024.470 ;
        RECT 1397.930 3023.290 1399.110 3024.470 ;
        RECT 1396.330 3021.690 1397.510 3022.870 ;
        RECT 1397.930 3021.690 1399.110 3022.870 ;
        RECT 1396.330 2843.290 1397.510 2844.470 ;
        RECT 1397.930 2843.290 1399.110 2844.470 ;
        RECT 1396.330 2841.690 1397.510 2842.870 ;
        RECT 1397.930 2841.690 1399.110 2842.870 ;
        RECT 1396.330 2663.290 1397.510 2664.470 ;
        RECT 1397.930 2663.290 1399.110 2664.470 ;
        RECT 1396.330 2661.690 1397.510 2662.870 ;
        RECT 1397.930 2661.690 1399.110 2662.870 ;
        RECT 1396.330 2483.290 1397.510 2484.470 ;
        RECT 1397.930 2483.290 1399.110 2484.470 ;
        RECT 1396.330 2481.690 1397.510 2482.870 ;
        RECT 1397.930 2481.690 1399.110 2482.870 ;
        RECT 1396.330 2303.290 1397.510 2304.470 ;
        RECT 1397.930 2303.290 1399.110 2304.470 ;
        RECT 1396.330 2301.690 1397.510 2302.870 ;
        RECT 1397.930 2301.690 1399.110 2302.870 ;
        RECT 1396.330 2123.290 1397.510 2124.470 ;
        RECT 1397.930 2123.290 1399.110 2124.470 ;
        RECT 1396.330 2121.690 1397.510 2122.870 ;
        RECT 1397.930 2121.690 1399.110 2122.870 ;
        RECT 1396.330 1943.290 1397.510 1944.470 ;
        RECT 1397.930 1943.290 1399.110 1944.470 ;
        RECT 1396.330 1941.690 1397.510 1942.870 ;
        RECT 1397.930 1941.690 1399.110 1942.870 ;
        RECT 1396.330 1763.290 1397.510 1764.470 ;
        RECT 1397.930 1763.290 1399.110 1764.470 ;
        RECT 1396.330 1761.690 1397.510 1762.870 ;
        RECT 1397.930 1761.690 1399.110 1762.870 ;
        RECT 1396.330 1583.290 1397.510 1584.470 ;
        RECT 1397.930 1583.290 1399.110 1584.470 ;
        RECT 1396.330 1581.690 1397.510 1582.870 ;
        RECT 1397.930 1581.690 1399.110 1582.870 ;
        RECT 1396.330 1403.290 1397.510 1404.470 ;
        RECT 1397.930 1403.290 1399.110 1404.470 ;
        RECT 1396.330 1401.690 1397.510 1402.870 ;
        RECT 1397.930 1401.690 1399.110 1402.870 ;
        RECT 1396.330 1223.290 1397.510 1224.470 ;
        RECT 1397.930 1223.290 1399.110 1224.470 ;
        RECT 1396.330 1221.690 1397.510 1222.870 ;
        RECT 1397.930 1221.690 1399.110 1222.870 ;
        RECT 1396.330 1043.290 1397.510 1044.470 ;
        RECT 1397.930 1043.290 1399.110 1044.470 ;
        RECT 1396.330 1041.690 1397.510 1042.870 ;
        RECT 1397.930 1041.690 1399.110 1042.870 ;
        RECT 1396.330 863.290 1397.510 864.470 ;
        RECT 1397.930 863.290 1399.110 864.470 ;
        RECT 1396.330 861.690 1397.510 862.870 ;
        RECT 1397.930 861.690 1399.110 862.870 ;
        RECT 1396.330 683.290 1397.510 684.470 ;
        RECT 1397.930 683.290 1399.110 684.470 ;
        RECT 1396.330 681.690 1397.510 682.870 ;
        RECT 1397.930 681.690 1399.110 682.870 ;
        RECT 1396.330 503.290 1397.510 504.470 ;
        RECT 1397.930 503.290 1399.110 504.470 ;
        RECT 1396.330 501.690 1397.510 502.870 ;
        RECT 1397.930 501.690 1399.110 502.870 ;
        RECT 1396.330 323.290 1397.510 324.470 ;
        RECT 1397.930 323.290 1399.110 324.470 ;
        RECT 1396.330 321.690 1397.510 322.870 ;
        RECT 1397.930 321.690 1399.110 322.870 ;
        RECT 1396.330 143.290 1397.510 144.470 ;
        RECT 1397.930 143.290 1399.110 144.470 ;
        RECT 1396.330 141.690 1397.510 142.870 ;
        RECT 1397.930 141.690 1399.110 142.870 ;
        RECT 1396.330 -26.910 1397.510 -25.730 ;
        RECT 1397.930 -26.910 1399.110 -25.730 ;
        RECT 1396.330 -28.510 1397.510 -27.330 ;
        RECT 1397.930 -28.510 1399.110 -27.330 ;
        RECT 1576.330 3547.010 1577.510 3548.190 ;
        RECT 1577.930 3547.010 1579.110 3548.190 ;
        RECT 1576.330 3545.410 1577.510 3546.590 ;
        RECT 1577.930 3545.410 1579.110 3546.590 ;
        RECT 1576.330 3383.290 1577.510 3384.470 ;
        RECT 1577.930 3383.290 1579.110 3384.470 ;
        RECT 1576.330 3381.690 1577.510 3382.870 ;
        RECT 1577.930 3381.690 1579.110 3382.870 ;
        RECT 1576.330 3203.290 1577.510 3204.470 ;
        RECT 1577.930 3203.290 1579.110 3204.470 ;
        RECT 1576.330 3201.690 1577.510 3202.870 ;
        RECT 1577.930 3201.690 1579.110 3202.870 ;
        RECT 1576.330 3023.290 1577.510 3024.470 ;
        RECT 1577.930 3023.290 1579.110 3024.470 ;
        RECT 1576.330 3021.690 1577.510 3022.870 ;
        RECT 1577.930 3021.690 1579.110 3022.870 ;
        RECT 1576.330 2843.290 1577.510 2844.470 ;
        RECT 1577.930 2843.290 1579.110 2844.470 ;
        RECT 1576.330 2841.690 1577.510 2842.870 ;
        RECT 1577.930 2841.690 1579.110 2842.870 ;
        RECT 1576.330 2663.290 1577.510 2664.470 ;
        RECT 1577.930 2663.290 1579.110 2664.470 ;
        RECT 1576.330 2661.690 1577.510 2662.870 ;
        RECT 1577.930 2661.690 1579.110 2662.870 ;
        RECT 1576.330 2483.290 1577.510 2484.470 ;
        RECT 1577.930 2483.290 1579.110 2484.470 ;
        RECT 1576.330 2481.690 1577.510 2482.870 ;
        RECT 1577.930 2481.690 1579.110 2482.870 ;
        RECT 1576.330 2303.290 1577.510 2304.470 ;
        RECT 1577.930 2303.290 1579.110 2304.470 ;
        RECT 1576.330 2301.690 1577.510 2302.870 ;
        RECT 1577.930 2301.690 1579.110 2302.870 ;
        RECT 1576.330 2123.290 1577.510 2124.470 ;
        RECT 1577.930 2123.290 1579.110 2124.470 ;
        RECT 1576.330 2121.690 1577.510 2122.870 ;
        RECT 1577.930 2121.690 1579.110 2122.870 ;
        RECT 1576.330 1943.290 1577.510 1944.470 ;
        RECT 1577.930 1943.290 1579.110 1944.470 ;
        RECT 1576.330 1941.690 1577.510 1942.870 ;
        RECT 1577.930 1941.690 1579.110 1942.870 ;
        RECT 1576.330 1763.290 1577.510 1764.470 ;
        RECT 1577.930 1763.290 1579.110 1764.470 ;
        RECT 1576.330 1761.690 1577.510 1762.870 ;
        RECT 1577.930 1761.690 1579.110 1762.870 ;
        RECT 1576.330 1583.290 1577.510 1584.470 ;
        RECT 1577.930 1583.290 1579.110 1584.470 ;
        RECT 1576.330 1581.690 1577.510 1582.870 ;
        RECT 1577.930 1581.690 1579.110 1582.870 ;
        RECT 1576.330 1403.290 1577.510 1404.470 ;
        RECT 1577.930 1403.290 1579.110 1404.470 ;
        RECT 1576.330 1401.690 1577.510 1402.870 ;
        RECT 1577.930 1401.690 1579.110 1402.870 ;
        RECT 1576.330 1223.290 1577.510 1224.470 ;
        RECT 1577.930 1223.290 1579.110 1224.470 ;
        RECT 1576.330 1221.690 1577.510 1222.870 ;
        RECT 1577.930 1221.690 1579.110 1222.870 ;
        RECT 1576.330 1043.290 1577.510 1044.470 ;
        RECT 1577.930 1043.290 1579.110 1044.470 ;
        RECT 1576.330 1041.690 1577.510 1042.870 ;
        RECT 1577.930 1041.690 1579.110 1042.870 ;
        RECT 1576.330 863.290 1577.510 864.470 ;
        RECT 1577.930 863.290 1579.110 864.470 ;
        RECT 1576.330 861.690 1577.510 862.870 ;
        RECT 1577.930 861.690 1579.110 862.870 ;
        RECT 1576.330 683.290 1577.510 684.470 ;
        RECT 1577.930 683.290 1579.110 684.470 ;
        RECT 1576.330 681.690 1577.510 682.870 ;
        RECT 1577.930 681.690 1579.110 682.870 ;
        RECT 1576.330 503.290 1577.510 504.470 ;
        RECT 1577.930 503.290 1579.110 504.470 ;
        RECT 1576.330 501.690 1577.510 502.870 ;
        RECT 1577.930 501.690 1579.110 502.870 ;
        RECT 1576.330 323.290 1577.510 324.470 ;
        RECT 1577.930 323.290 1579.110 324.470 ;
        RECT 1576.330 321.690 1577.510 322.870 ;
        RECT 1577.930 321.690 1579.110 322.870 ;
        RECT 1576.330 143.290 1577.510 144.470 ;
        RECT 1577.930 143.290 1579.110 144.470 ;
        RECT 1576.330 141.690 1577.510 142.870 ;
        RECT 1577.930 141.690 1579.110 142.870 ;
        RECT 1576.330 -26.910 1577.510 -25.730 ;
        RECT 1577.930 -26.910 1579.110 -25.730 ;
        RECT 1576.330 -28.510 1577.510 -27.330 ;
        RECT 1577.930 -28.510 1579.110 -27.330 ;
        RECT 1756.330 3547.010 1757.510 3548.190 ;
        RECT 1757.930 3547.010 1759.110 3548.190 ;
        RECT 1756.330 3545.410 1757.510 3546.590 ;
        RECT 1757.930 3545.410 1759.110 3546.590 ;
        RECT 1756.330 3383.290 1757.510 3384.470 ;
        RECT 1757.930 3383.290 1759.110 3384.470 ;
        RECT 1756.330 3381.690 1757.510 3382.870 ;
        RECT 1757.930 3381.690 1759.110 3382.870 ;
        RECT 1756.330 3203.290 1757.510 3204.470 ;
        RECT 1757.930 3203.290 1759.110 3204.470 ;
        RECT 1756.330 3201.690 1757.510 3202.870 ;
        RECT 1757.930 3201.690 1759.110 3202.870 ;
        RECT 1756.330 3023.290 1757.510 3024.470 ;
        RECT 1757.930 3023.290 1759.110 3024.470 ;
        RECT 1756.330 3021.690 1757.510 3022.870 ;
        RECT 1757.930 3021.690 1759.110 3022.870 ;
        RECT 1756.330 2843.290 1757.510 2844.470 ;
        RECT 1757.930 2843.290 1759.110 2844.470 ;
        RECT 1756.330 2841.690 1757.510 2842.870 ;
        RECT 1757.930 2841.690 1759.110 2842.870 ;
        RECT 1756.330 2663.290 1757.510 2664.470 ;
        RECT 1757.930 2663.290 1759.110 2664.470 ;
        RECT 1756.330 2661.690 1757.510 2662.870 ;
        RECT 1757.930 2661.690 1759.110 2662.870 ;
        RECT 1756.330 2483.290 1757.510 2484.470 ;
        RECT 1757.930 2483.290 1759.110 2484.470 ;
        RECT 1756.330 2481.690 1757.510 2482.870 ;
        RECT 1757.930 2481.690 1759.110 2482.870 ;
        RECT 1756.330 2303.290 1757.510 2304.470 ;
        RECT 1757.930 2303.290 1759.110 2304.470 ;
        RECT 1756.330 2301.690 1757.510 2302.870 ;
        RECT 1757.930 2301.690 1759.110 2302.870 ;
        RECT 1756.330 2123.290 1757.510 2124.470 ;
        RECT 1757.930 2123.290 1759.110 2124.470 ;
        RECT 1756.330 2121.690 1757.510 2122.870 ;
        RECT 1757.930 2121.690 1759.110 2122.870 ;
        RECT 1756.330 1943.290 1757.510 1944.470 ;
        RECT 1757.930 1943.290 1759.110 1944.470 ;
        RECT 1756.330 1941.690 1757.510 1942.870 ;
        RECT 1757.930 1941.690 1759.110 1942.870 ;
        RECT 1756.330 1763.290 1757.510 1764.470 ;
        RECT 1757.930 1763.290 1759.110 1764.470 ;
        RECT 1756.330 1761.690 1757.510 1762.870 ;
        RECT 1757.930 1761.690 1759.110 1762.870 ;
        RECT 1756.330 1583.290 1757.510 1584.470 ;
        RECT 1757.930 1583.290 1759.110 1584.470 ;
        RECT 1756.330 1581.690 1757.510 1582.870 ;
        RECT 1757.930 1581.690 1759.110 1582.870 ;
        RECT 1756.330 1403.290 1757.510 1404.470 ;
        RECT 1757.930 1403.290 1759.110 1404.470 ;
        RECT 1756.330 1401.690 1757.510 1402.870 ;
        RECT 1757.930 1401.690 1759.110 1402.870 ;
        RECT 1756.330 1223.290 1757.510 1224.470 ;
        RECT 1757.930 1223.290 1759.110 1224.470 ;
        RECT 1756.330 1221.690 1757.510 1222.870 ;
        RECT 1757.930 1221.690 1759.110 1222.870 ;
        RECT 1756.330 1043.290 1757.510 1044.470 ;
        RECT 1757.930 1043.290 1759.110 1044.470 ;
        RECT 1756.330 1041.690 1757.510 1042.870 ;
        RECT 1757.930 1041.690 1759.110 1042.870 ;
        RECT 1756.330 863.290 1757.510 864.470 ;
        RECT 1757.930 863.290 1759.110 864.470 ;
        RECT 1756.330 861.690 1757.510 862.870 ;
        RECT 1757.930 861.690 1759.110 862.870 ;
        RECT 1756.330 683.290 1757.510 684.470 ;
        RECT 1757.930 683.290 1759.110 684.470 ;
        RECT 1756.330 681.690 1757.510 682.870 ;
        RECT 1757.930 681.690 1759.110 682.870 ;
        RECT 1756.330 503.290 1757.510 504.470 ;
        RECT 1757.930 503.290 1759.110 504.470 ;
        RECT 1756.330 501.690 1757.510 502.870 ;
        RECT 1757.930 501.690 1759.110 502.870 ;
        RECT 1756.330 323.290 1757.510 324.470 ;
        RECT 1757.930 323.290 1759.110 324.470 ;
        RECT 1756.330 321.690 1757.510 322.870 ;
        RECT 1757.930 321.690 1759.110 322.870 ;
        RECT 1756.330 143.290 1757.510 144.470 ;
        RECT 1757.930 143.290 1759.110 144.470 ;
        RECT 1756.330 141.690 1757.510 142.870 ;
        RECT 1757.930 141.690 1759.110 142.870 ;
        RECT 1756.330 -26.910 1757.510 -25.730 ;
        RECT 1757.930 -26.910 1759.110 -25.730 ;
        RECT 1756.330 -28.510 1757.510 -27.330 ;
        RECT 1757.930 -28.510 1759.110 -27.330 ;
        RECT 1936.330 3547.010 1937.510 3548.190 ;
        RECT 1937.930 3547.010 1939.110 3548.190 ;
        RECT 1936.330 3545.410 1937.510 3546.590 ;
        RECT 1937.930 3545.410 1939.110 3546.590 ;
        RECT 1936.330 3383.290 1937.510 3384.470 ;
        RECT 1937.930 3383.290 1939.110 3384.470 ;
        RECT 1936.330 3381.690 1937.510 3382.870 ;
        RECT 1937.930 3381.690 1939.110 3382.870 ;
        RECT 1936.330 3203.290 1937.510 3204.470 ;
        RECT 1937.930 3203.290 1939.110 3204.470 ;
        RECT 1936.330 3201.690 1937.510 3202.870 ;
        RECT 1937.930 3201.690 1939.110 3202.870 ;
        RECT 1936.330 3023.290 1937.510 3024.470 ;
        RECT 1937.930 3023.290 1939.110 3024.470 ;
        RECT 1936.330 3021.690 1937.510 3022.870 ;
        RECT 1937.930 3021.690 1939.110 3022.870 ;
        RECT 1936.330 2843.290 1937.510 2844.470 ;
        RECT 1937.930 2843.290 1939.110 2844.470 ;
        RECT 1936.330 2841.690 1937.510 2842.870 ;
        RECT 1937.930 2841.690 1939.110 2842.870 ;
        RECT 1936.330 2663.290 1937.510 2664.470 ;
        RECT 1937.930 2663.290 1939.110 2664.470 ;
        RECT 1936.330 2661.690 1937.510 2662.870 ;
        RECT 1937.930 2661.690 1939.110 2662.870 ;
        RECT 1936.330 2483.290 1937.510 2484.470 ;
        RECT 1937.930 2483.290 1939.110 2484.470 ;
        RECT 1936.330 2481.690 1937.510 2482.870 ;
        RECT 1937.930 2481.690 1939.110 2482.870 ;
        RECT 1936.330 2303.290 1937.510 2304.470 ;
        RECT 1937.930 2303.290 1939.110 2304.470 ;
        RECT 1936.330 2301.690 1937.510 2302.870 ;
        RECT 1937.930 2301.690 1939.110 2302.870 ;
        RECT 1936.330 2123.290 1937.510 2124.470 ;
        RECT 1937.930 2123.290 1939.110 2124.470 ;
        RECT 1936.330 2121.690 1937.510 2122.870 ;
        RECT 1937.930 2121.690 1939.110 2122.870 ;
        RECT 1936.330 1943.290 1937.510 1944.470 ;
        RECT 1937.930 1943.290 1939.110 1944.470 ;
        RECT 1936.330 1941.690 1937.510 1942.870 ;
        RECT 1937.930 1941.690 1939.110 1942.870 ;
        RECT 1936.330 1763.290 1937.510 1764.470 ;
        RECT 1937.930 1763.290 1939.110 1764.470 ;
        RECT 1936.330 1761.690 1937.510 1762.870 ;
        RECT 1937.930 1761.690 1939.110 1762.870 ;
        RECT 1936.330 1583.290 1937.510 1584.470 ;
        RECT 1937.930 1583.290 1939.110 1584.470 ;
        RECT 1936.330 1581.690 1937.510 1582.870 ;
        RECT 1937.930 1581.690 1939.110 1582.870 ;
        RECT 1936.330 1403.290 1937.510 1404.470 ;
        RECT 1937.930 1403.290 1939.110 1404.470 ;
        RECT 1936.330 1401.690 1937.510 1402.870 ;
        RECT 1937.930 1401.690 1939.110 1402.870 ;
        RECT 1936.330 1223.290 1937.510 1224.470 ;
        RECT 1937.930 1223.290 1939.110 1224.470 ;
        RECT 1936.330 1221.690 1937.510 1222.870 ;
        RECT 1937.930 1221.690 1939.110 1222.870 ;
        RECT 1936.330 1043.290 1937.510 1044.470 ;
        RECT 1937.930 1043.290 1939.110 1044.470 ;
        RECT 1936.330 1041.690 1937.510 1042.870 ;
        RECT 1937.930 1041.690 1939.110 1042.870 ;
        RECT 1936.330 863.290 1937.510 864.470 ;
        RECT 1937.930 863.290 1939.110 864.470 ;
        RECT 1936.330 861.690 1937.510 862.870 ;
        RECT 1937.930 861.690 1939.110 862.870 ;
        RECT 1936.330 683.290 1937.510 684.470 ;
        RECT 1937.930 683.290 1939.110 684.470 ;
        RECT 1936.330 681.690 1937.510 682.870 ;
        RECT 1937.930 681.690 1939.110 682.870 ;
        RECT 1936.330 503.290 1937.510 504.470 ;
        RECT 1937.930 503.290 1939.110 504.470 ;
        RECT 1936.330 501.690 1937.510 502.870 ;
        RECT 1937.930 501.690 1939.110 502.870 ;
        RECT 1936.330 323.290 1937.510 324.470 ;
        RECT 1937.930 323.290 1939.110 324.470 ;
        RECT 1936.330 321.690 1937.510 322.870 ;
        RECT 1937.930 321.690 1939.110 322.870 ;
        RECT 1936.330 143.290 1937.510 144.470 ;
        RECT 1937.930 143.290 1939.110 144.470 ;
        RECT 1936.330 141.690 1937.510 142.870 ;
        RECT 1937.930 141.690 1939.110 142.870 ;
        RECT 1936.330 -26.910 1937.510 -25.730 ;
        RECT 1937.930 -26.910 1939.110 -25.730 ;
        RECT 1936.330 -28.510 1937.510 -27.330 ;
        RECT 1937.930 -28.510 1939.110 -27.330 ;
        RECT 2116.330 3547.010 2117.510 3548.190 ;
        RECT 2117.930 3547.010 2119.110 3548.190 ;
        RECT 2116.330 3545.410 2117.510 3546.590 ;
        RECT 2117.930 3545.410 2119.110 3546.590 ;
        RECT 2116.330 3383.290 2117.510 3384.470 ;
        RECT 2117.930 3383.290 2119.110 3384.470 ;
        RECT 2116.330 3381.690 2117.510 3382.870 ;
        RECT 2117.930 3381.690 2119.110 3382.870 ;
        RECT 2116.330 3203.290 2117.510 3204.470 ;
        RECT 2117.930 3203.290 2119.110 3204.470 ;
        RECT 2116.330 3201.690 2117.510 3202.870 ;
        RECT 2117.930 3201.690 2119.110 3202.870 ;
        RECT 2116.330 3023.290 2117.510 3024.470 ;
        RECT 2117.930 3023.290 2119.110 3024.470 ;
        RECT 2116.330 3021.690 2117.510 3022.870 ;
        RECT 2117.930 3021.690 2119.110 3022.870 ;
        RECT 2116.330 2843.290 2117.510 2844.470 ;
        RECT 2117.930 2843.290 2119.110 2844.470 ;
        RECT 2116.330 2841.690 2117.510 2842.870 ;
        RECT 2117.930 2841.690 2119.110 2842.870 ;
        RECT 2116.330 2663.290 2117.510 2664.470 ;
        RECT 2117.930 2663.290 2119.110 2664.470 ;
        RECT 2116.330 2661.690 2117.510 2662.870 ;
        RECT 2117.930 2661.690 2119.110 2662.870 ;
        RECT 2116.330 2483.290 2117.510 2484.470 ;
        RECT 2117.930 2483.290 2119.110 2484.470 ;
        RECT 2116.330 2481.690 2117.510 2482.870 ;
        RECT 2117.930 2481.690 2119.110 2482.870 ;
        RECT 2116.330 2303.290 2117.510 2304.470 ;
        RECT 2117.930 2303.290 2119.110 2304.470 ;
        RECT 2116.330 2301.690 2117.510 2302.870 ;
        RECT 2117.930 2301.690 2119.110 2302.870 ;
        RECT 2116.330 2123.290 2117.510 2124.470 ;
        RECT 2117.930 2123.290 2119.110 2124.470 ;
        RECT 2116.330 2121.690 2117.510 2122.870 ;
        RECT 2117.930 2121.690 2119.110 2122.870 ;
        RECT 2116.330 1943.290 2117.510 1944.470 ;
        RECT 2117.930 1943.290 2119.110 1944.470 ;
        RECT 2116.330 1941.690 2117.510 1942.870 ;
        RECT 2117.930 1941.690 2119.110 1942.870 ;
        RECT 2116.330 1763.290 2117.510 1764.470 ;
        RECT 2117.930 1763.290 2119.110 1764.470 ;
        RECT 2116.330 1761.690 2117.510 1762.870 ;
        RECT 2117.930 1761.690 2119.110 1762.870 ;
        RECT 2116.330 1583.290 2117.510 1584.470 ;
        RECT 2117.930 1583.290 2119.110 1584.470 ;
        RECT 2116.330 1581.690 2117.510 1582.870 ;
        RECT 2117.930 1581.690 2119.110 1582.870 ;
        RECT 2116.330 1403.290 2117.510 1404.470 ;
        RECT 2117.930 1403.290 2119.110 1404.470 ;
        RECT 2116.330 1401.690 2117.510 1402.870 ;
        RECT 2117.930 1401.690 2119.110 1402.870 ;
        RECT 2116.330 1223.290 2117.510 1224.470 ;
        RECT 2117.930 1223.290 2119.110 1224.470 ;
        RECT 2116.330 1221.690 2117.510 1222.870 ;
        RECT 2117.930 1221.690 2119.110 1222.870 ;
        RECT 2116.330 1043.290 2117.510 1044.470 ;
        RECT 2117.930 1043.290 2119.110 1044.470 ;
        RECT 2116.330 1041.690 2117.510 1042.870 ;
        RECT 2117.930 1041.690 2119.110 1042.870 ;
        RECT 2116.330 863.290 2117.510 864.470 ;
        RECT 2117.930 863.290 2119.110 864.470 ;
        RECT 2116.330 861.690 2117.510 862.870 ;
        RECT 2117.930 861.690 2119.110 862.870 ;
        RECT 2116.330 683.290 2117.510 684.470 ;
        RECT 2117.930 683.290 2119.110 684.470 ;
        RECT 2116.330 681.690 2117.510 682.870 ;
        RECT 2117.930 681.690 2119.110 682.870 ;
        RECT 2116.330 503.290 2117.510 504.470 ;
        RECT 2117.930 503.290 2119.110 504.470 ;
        RECT 2116.330 501.690 2117.510 502.870 ;
        RECT 2117.930 501.690 2119.110 502.870 ;
        RECT 2116.330 323.290 2117.510 324.470 ;
        RECT 2117.930 323.290 2119.110 324.470 ;
        RECT 2116.330 321.690 2117.510 322.870 ;
        RECT 2117.930 321.690 2119.110 322.870 ;
        RECT 2116.330 143.290 2117.510 144.470 ;
        RECT 2117.930 143.290 2119.110 144.470 ;
        RECT 2116.330 141.690 2117.510 142.870 ;
        RECT 2117.930 141.690 2119.110 142.870 ;
        RECT 2116.330 -26.910 2117.510 -25.730 ;
        RECT 2117.930 -26.910 2119.110 -25.730 ;
        RECT 2116.330 -28.510 2117.510 -27.330 ;
        RECT 2117.930 -28.510 2119.110 -27.330 ;
        RECT 2296.330 3547.010 2297.510 3548.190 ;
        RECT 2297.930 3547.010 2299.110 3548.190 ;
        RECT 2296.330 3545.410 2297.510 3546.590 ;
        RECT 2297.930 3545.410 2299.110 3546.590 ;
        RECT 2296.330 3383.290 2297.510 3384.470 ;
        RECT 2297.930 3383.290 2299.110 3384.470 ;
        RECT 2296.330 3381.690 2297.510 3382.870 ;
        RECT 2297.930 3381.690 2299.110 3382.870 ;
        RECT 2296.330 3203.290 2297.510 3204.470 ;
        RECT 2297.930 3203.290 2299.110 3204.470 ;
        RECT 2296.330 3201.690 2297.510 3202.870 ;
        RECT 2297.930 3201.690 2299.110 3202.870 ;
        RECT 2296.330 3023.290 2297.510 3024.470 ;
        RECT 2297.930 3023.290 2299.110 3024.470 ;
        RECT 2296.330 3021.690 2297.510 3022.870 ;
        RECT 2297.930 3021.690 2299.110 3022.870 ;
        RECT 2296.330 2843.290 2297.510 2844.470 ;
        RECT 2297.930 2843.290 2299.110 2844.470 ;
        RECT 2296.330 2841.690 2297.510 2842.870 ;
        RECT 2297.930 2841.690 2299.110 2842.870 ;
        RECT 2296.330 2663.290 2297.510 2664.470 ;
        RECT 2297.930 2663.290 2299.110 2664.470 ;
        RECT 2296.330 2661.690 2297.510 2662.870 ;
        RECT 2297.930 2661.690 2299.110 2662.870 ;
        RECT 2296.330 2483.290 2297.510 2484.470 ;
        RECT 2297.930 2483.290 2299.110 2484.470 ;
        RECT 2296.330 2481.690 2297.510 2482.870 ;
        RECT 2297.930 2481.690 2299.110 2482.870 ;
        RECT 2296.330 2303.290 2297.510 2304.470 ;
        RECT 2297.930 2303.290 2299.110 2304.470 ;
        RECT 2296.330 2301.690 2297.510 2302.870 ;
        RECT 2297.930 2301.690 2299.110 2302.870 ;
        RECT 2296.330 2123.290 2297.510 2124.470 ;
        RECT 2297.930 2123.290 2299.110 2124.470 ;
        RECT 2296.330 2121.690 2297.510 2122.870 ;
        RECT 2297.930 2121.690 2299.110 2122.870 ;
        RECT 2296.330 1943.290 2297.510 1944.470 ;
        RECT 2297.930 1943.290 2299.110 1944.470 ;
        RECT 2296.330 1941.690 2297.510 1942.870 ;
        RECT 2297.930 1941.690 2299.110 1942.870 ;
        RECT 2296.330 1763.290 2297.510 1764.470 ;
        RECT 2297.930 1763.290 2299.110 1764.470 ;
        RECT 2296.330 1761.690 2297.510 1762.870 ;
        RECT 2297.930 1761.690 2299.110 1762.870 ;
        RECT 2296.330 1583.290 2297.510 1584.470 ;
        RECT 2297.930 1583.290 2299.110 1584.470 ;
        RECT 2296.330 1581.690 2297.510 1582.870 ;
        RECT 2297.930 1581.690 2299.110 1582.870 ;
        RECT 2296.330 1403.290 2297.510 1404.470 ;
        RECT 2297.930 1403.290 2299.110 1404.470 ;
        RECT 2296.330 1401.690 2297.510 1402.870 ;
        RECT 2297.930 1401.690 2299.110 1402.870 ;
        RECT 2296.330 1223.290 2297.510 1224.470 ;
        RECT 2297.930 1223.290 2299.110 1224.470 ;
        RECT 2296.330 1221.690 2297.510 1222.870 ;
        RECT 2297.930 1221.690 2299.110 1222.870 ;
        RECT 2296.330 1043.290 2297.510 1044.470 ;
        RECT 2297.930 1043.290 2299.110 1044.470 ;
        RECT 2296.330 1041.690 2297.510 1042.870 ;
        RECT 2297.930 1041.690 2299.110 1042.870 ;
        RECT 2296.330 863.290 2297.510 864.470 ;
        RECT 2297.930 863.290 2299.110 864.470 ;
        RECT 2296.330 861.690 2297.510 862.870 ;
        RECT 2297.930 861.690 2299.110 862.870 ;
        RECT 2296.330 683.290 2297.510 684.470 ;
        RECT 2297.930 683.290 2299.110 684.470 ;
        RECT 2296.330 681.690 2297.510 682.870 ;
        RECT 2297.930 681.690 2299.110 682.870 ;
        RECT 2296.330 503.290 2297.510 504.470 ;
        RECT 2297.930 503.290 2299.110 504.470 ;
        RECT 2296.330 501.690 2297.510 502.870 ;
        RECT 2297.930 501.690 2299.110 502.870 ;
        RECT 2296.330 323.290 2297.510 324.470 ;
        RECT 2297.930 323.290 2299.110 324.470 ;
        RECT 2296.330 321.690 2297.510 322.870 ;
        RECT 2297.930 321.690 2299.110 322.870 ;
        RECT 2296.330 143.290 2297.510 144.470 ;
        RECT 2297.930 143.290 2299.110 144.470 ;
        RECT 2296.330 141.690 2297.510 142.870 ;
        RECT 2297.930 141.690 2299.110 142.870 ;
        RECT 2296.330 -26.910 2297.510 -25.730 ;
        RECT 2297.930 -26.910 2299.110 -25.730 ;
        RECT 2296.330 -28.510 2297.510 -27.330 ;
        RECT 2297.930 -28.510 2299.110 -27.330 ;
        RECT 2476.330 3547.010 2477.510 3548.190 ;
        RECT 2477.930 3547.010 2479.110 3548.190 ;
        RECT 2476.330 3545.410 2477.510 3546.590 ;
        RECT 2477.930 3545.410 2479.110 3546.590 ;
        RECT 2476.330 3383.290 2477.510 3384.470 ;
        RECT 2477.930 3383.290 2479.110 3384.470 ;
        RECT 2476.330 3381.690 2477.510 3382.870 ;
        RECT 2477.930 3381.690 2479.110 3382.870 ;
        RECT 2476.330 3203.290 2477.510 3204.470 ;
        RECT 2477.930 3203.290 2479.110 3204.470 ;
        RECT 2476.330 3201.690 2477.510 3202.870 ;
        RECT 2477.930 3201.690 2479.110 3202.870 ;
        RECT 2476.330 3023.290 2477.510 3024.470 ;
        RECT 2477.930 3023.290 2479.110 3024.470 ;
        RECT 2476.330 3021.690 2477.510 3022.870 ;
        RECT 2477.930 3021.690 2479.110 3022.870 ;
        RECT 2476.330 2843.290 2477.510 2844.470 ;
        RECT 2477.930 2843.290 2479.110 2844.470 ;
        RECT 2476.330 2841.690 2477.510 2842.870 ;
        RECT 2477.930 2841.690 2479.110 2842.870 ;
        RECT 2476.330 2663.290 2477.510 2664.470 ;
        RECT 2477.930 2663.290 2479.110 2664.470 ;
        RECT 2476.330 2661.690 2477.510 2662.870 ;
        RECT 2477.930 2661.690 2479.110 2662.870 ;
        RECT 2476.330 2483.290 2477.510 2484.470 ;
        RECT 2477.930 2483.290 2479.110 2484.470 ;
        RECT 2476.330 2481.690 2477.510 2482.870 ;
        RECT 2477.930 2481.690 2479.110 2482.870 ;
        RECT 2476.330 2303.290 2477.510 2304.470 ;
        RECT 2477.930 2303.290 2479.110 2304.470 ;
        RECT 2476.330 2301.690 2477.510 2302.870 ;
        RECT 2477.930 2301.690 2479.110 2302.870 ;
        RECT 2476.330 2123.290 2477.510 2124.470 ;
        RECT 2477.930 2123.290 2479.110 2124.470 ;
        RECT 2476.330 2121.690 2477.510 2122.870 ;
        RECT 2477.930 2121.690 2479.110 2122.870 ;
        RECT 2476.330 1943.290 2477.510 1944.470 ;
        RECT 2477.930 1943.290 2479.110 1944.470 ;
        RECT 2476.330 1941.690 2477.510 1942.870 ;
        RECT 2477.930 1941.690 2479.110 1942.870 ;
        RECT 2476.330 1763.290 2477.510 1764.470 ;
        RECT 2477.930 1763.290 2479.110 1764.470 ;
        RECT 2476.330 1761.690 2477.510 1762.870 ;
        RECT 2477.930 1761.690 2479.110 1762.870 ;
        RECT 2476.330 1583.290 2477.510 1584.470 ;
        RECT 2477.930 1583.290 2479.110 1584.470 ;
        RECT 2476.330 1581.690 2477.510 1582.870 ;
        RECT 2477.930 1581.690 2479.110 1582.870 ;
        RECT 2476.330 1403.290 2477.510 1404.470 ;
        RECT 2477.930 1403.290 2479.110 1404.470 ;
        RECT 2476.330 1401.690 2477.510 1402.870 ;
        RECT 2477.930 1401.690 2479.110 1402.870 ;
        RECT 2476.330 1223.290 2477.510 1224.470 ;
        RECT 2477.930 1223.290 2479.110 1224.470 ;
        RECT 2476.330 1221.690 2477.510 1222.870 ;
        RECT 2477.930 1221.690 2479.110 1222.870 ;
        RECT 2476.330 1043.290 2477.510 1044.470 ;
        RECT 2477.930 1043.290 2479.110 1044.470 ;
        RECT 2476.330 1041.690 2477.510 1042.870 ;
        RECT 2477.930 1041.690 2479.110 1042.870 ;
        RECT 2476.330 863.290 2477.510 864.470 ;
        RECT 2477.930 863.290 2479.110 864.470 ;
        RECT 2476.330 861.690 2477.510 862.870 ;
        RECT 2477.930 861.690 2479.110 862.870 ;
        RECT 2476.330 683.290 2477.510 684.470 ;
        RECT 2477.930 683.290 2479.110 684.470 ;
        RECT 2476.330 681.690 2477.510 682.870 ;
        RECT 2477.930 681.690 2479.110 682.870 ;
        RECT 2476.330 503.290 2477.510 504.470 ;
        RECT 2477.930 503.290 2479.110 504.470 ;
        RECT 2476.330 501.690 2477.510 502.870 ;
        RECT 2477.930 501.690 2479.110 502.870 ;
        RECT 2476.330 323.290 2477.510 324.470 ;
        RECT 2477.930 323.290 2479.110 324.470 ;
        RECT 2476.330 321.690 2477.510 322.870 ;
        RECT 2477.930 321.690 2479.110 322.870 ;
        RECT 2476.330 143.290 2477.510 144.470 ;
        RECT 2477.930 143.290 2479.110 144.470 ;
        RECT 2476.330 141.690 2477.510 142.870 ;
        RECT 2477.930 141.690 2479.110 142.870 ;
        RECT 2476.330 -26.910 2477.510 -25.730 ;
        RECT 2477.930 -26.910 2479.110 -25.730 ;
        RECT 2476.330 -28.510 2477.510 -27.330 ;
        RECT 2477.930 -28.510 2479.110 -27.330 ;
        RECT 2656.330 3547.010 2657.510 3548.190 ;
        RECT 2657.930 3547.010 2659.110 3548.190 ;
        RECT 2656.330 3545.410 2657.510 3546.590 ;
        RECT 2657.930 3545.410 2659.110 3546.590 ;
        RECT 2656.330 3383.290 2657.510 3384.470 ;
        RECT 2657.930 3383.290 2659.110 3384.470 ;
        RECT 2656.330 3381.690 2657.510 3382.870 ;
        RECT 2657.930 3381.690 2659.110 3382.870 ;
        RECT 2656.330 3203.290 2657.510 3204.470 ;
        RECT 2657.930 3203.290 2659.110 3204.470 ;
        RECT 2656.330 3201.690 2657.510 3202.870 ;
        RECT 2657.930 3201.690 2659.110 3202.870 ;
        RECT 2656.330 3023.290 2657.510 3024.470 ;
        RECT 2657.930 3023.290 2659.110 3024.470 ;
        RECT 2656.330 3021.690 2657.510 3022.870 ;
        RECT 2657.930 3021.690 2659.110 3022.870 ;
        RECT 2656.330 2843.290 2657.510 2844.470 ;
        RECT 2657.930 2843.290 2659.110 2844.470 ;
        RECT 2656.330 2841.690 2657.510 2842.870 ;
        RECT 2657.930 2841.690 2659.110 2842.870 ;
        RECT 2656.330 2663.290 2657.510 2664.470 ;
        RECT 2657.930 2663.290 2659.110 2664.470 ;
        RECT 2656.330 2661.690 2657.510 2662.870 ;
        RECT 2657.930 2661.690 2659.110 2662.870 ;
        RECT 2656.330 2483.290 2657.510 2484.470 ;
        RECT 2657.930 2483.290 2659.110 2484.470 ;
        RECT 2656.330 2481.690 2657.510 2482.870 ;
        RECT 2657.930 2481.690 2659.110 2482.870 ;
        RECT 2656.330 2303.290 2657.510 2304.470 ;
        RECT 2657.930 2303.290 2659.110 2304.470 ;
        RECT 2656.330 2301.690 2657.510 2302.870 ;
        RECT 2657.930 2301.690 2659.110 2302.870 ;
        RECT 2656.330 2123.290 2657.510 2124.470 ;
        RECT 2657.930 2123.290 2659.110 2124.470 ;
        RECT 2656.330 2121.690 2657.510 2122.870 ;
        RECT 2657.930 2121.690 2659.110 2122.870 ;
        RECT 2656.330 1943.290 2657.510 1944.470 ;
        RECT 2657.930 1943.290 2659.110 1944.470 ;
        RECT 2656.330 1941.690 2657.510 1942.870 ;
        RECT 2657.930 1941.690 2659.110 1942.870 ;
        RECT 2656.330 1763.290 2657.510 1764.470 ;
        RECT 2657.930 1763.290 2659.110 1764.470 ;
        RECT 2656.330 1761.690 2657.510 1762.870 ;
        RECT 2657.930 1761.690 2659.110 1762.870 ;
        RECT 2656.330 1583.290 2657.510 1584.470 ;
        RECT 2657.930 1583.290 2659.110 1584.470 ;
        RECT 2656.330 1581.690 2657.510 1582.870 ;
        RECT 2657.930 1581.690 2659.110 1582.870 ;
        RECT 2656.330 1403.290 2657.510 1404.470 ;
        RECT 2657.930 1403.290 2659.110 1404.470 ;
        RECT 2656.330 1401.690 2657.510 1402.870 ;
        RECT 2657.930 1401.690 2659.110 1402.870 ;
        RECT 2656.330 1223.290 2657.510 1224.470 ;
        RECT 2657.930 1223.290 2659.110 1224.470 ;
        RECT 2656.330 1221.690 2657.510 1222.870 ;
        RECT 2657.930 1221.690 2659.110 1222.870 ;
        RECT 2656.330 1043.290 2657.510 1044.470 ;
        RECT 2657.930 1043.290 2659.110 1044.470 ;
        RECT 2656.330 1041.690 2657.510 1042.870 ;
        RECT 2657.930 1041.690 2659.110 1042.870 ;
        RECT 2656.330 863.290 2657.510 864.470 ;
        RECT 2657.930 863.290 2659.110 864.470 ;
        RECT 2656.330 861.690 2657.510 862.870 ;
        RECT 2657.930 861.690 2659.110 862.870 ;
        RECT 2656.330 683.290 2657.510 684.470 ;
        RECT 2657.930 683.290 2659.110 684.470 ;
        RECT 2656.330 681.690 2657.510 682.870 ;
        RECT 2657.930 681.690 2659.110 682.870 ;
        RECT 2656.330 503.290 2657.510 504.470 ;
        RECT 2657.930 503.290 2659.110 504.470 ;
        RECT 2656.330 501.690 2657.510 502.870 ;
        RECT 2657.930 501.690 2659.110 502.870 ;
        RECT 2656.330 323.290 2657.510 324.470 ;
        RECT 2657.930 323.290 2659.110 324.470 ;
        RECT 2656.330 321.690 2657.510 322.870 ;
        RECT 2657.930 321.690 2659.110 322.870 ;
        RECT 2656.330 143.290 2657.510 144.470 ;
        RECT 2657.930 143.290 2659.110 144.470 ;
        RECT 2656.330 141.690 2657.510 142.870 ;
        RECT 2657.930 141.690 2659.110 142.870 ;
        RECT 2656.330 -26.910 2657.510 -25.730 ;
        RECT 2657.930 -26.910 2659.110 -25.730 ;
        RECT 2656.330 -28.510 2657.510 -27.330 ;
        RECT 2657.930 -28.510 2659.110 -27.330 ;
        RECT 2836.330 3547.010 2837.510 3548.190 ;
        RECT 2837.930 3547.010 2839.110 3548.190 ;
        RECT 2836.330 3545.410 2837.510 3546.590 ;
        RECT 2837.930 3545.410 2839.110 3546.590 ;
        RECT 2836.330 3383.290 2837.510 3384.470 ;
        RECT 2837.930 3383.290 2839.110 3384.470 ;
        RECT 2836.330 3381.690 2837.510 3382.870 ;
        RECT 2837.930 3381.690 2839.110 3382.870 ;
        RECT 2836.330 3203.290 2837.510 3204.470 ;
        RECT 2837.930 3203.290 2839.110 3204.470 ;
        RECT 2836.330 3201.690 2837.510 3202.870 ;
        RECT 2837.930 3201.690 2839.110 3202.870 ;
        RECT 2836.330 3023.290 2837.510 3024.470 ;
        RECT 2837.930 3023.290 2839.110 3024.470 ;
        RECT 2836.330 3021.690 2837.510 3022.870 ;
        RECT 2837.930 3021.690 2839.110 3022.870 ;
        RECT 2836.330 2843.290 2837.510 2844.470 ;
        RECT 2837.930 2843.290 2839.110 2844.470 ;
        RECT 2836.330 2841.690 2837.510 2842.870 ;
        RECT 2837.930 2841.690 2839.110 2842.870 ;
        RECT 2836.330 2663.290 2837.510 2664.470 ;
        RECT 2837.930 2663.290 2839.110 2664.470 ;
        RECT 2836.330 2661.690 2837.510 2662.870 ;
        RECT 2837.930 2661.690 2839.110 2662.870 ;
        RECT 2836.330 2483.290 2837.510 2484.470 ;
        RECT 2837.930 2483.290 2839.110 2484.470 ;
        RECT 2836.330 2481.690 2837.510 2482.870 ;
        RECT 2837.930 2481.690 2839.110 2482.870 ;
        RECT 2836.330 2303.290 2837.510 2304.470 ;
        RECT 2837.930 2303.290 2839.110 2304.470 ;
        RECT 2836.330 2301.690 2837.510 2302.870 ;
        RECT 2837.930 2301.690 2839.110 2302.870 ;
        RECT 2836.330 2123.290 2837.510 2124.470 ;
        RECT 2837.930 2123.290 2839.110 2124.470 ;
        RECT 2836.330 2121.690 2837.510 2122.870 ;
        RECT 2837.930 2121.690 2839.110 2122.870 ;
        RECT 2836.330 1943.290 2837.510 1944.470 ;
        RECT 2837.930 1943.290 2839.110 1944.470 ;
        RECT 2836.330 1941.690 2837.510 1942.870 ;
        RECT 2837.930 1941.690 2839.110 1942.870 ;
        RECT 2836.330 1763.290 2837.510 1764.470 ;
        RECT 2837.930 1763.290 2839.110 1764.470 ;
        RECT 2836.330 1761.690 2837.510 1762.870 ;
        RECT 2837.930 1761.690 2839.110 1762.870 ;
        RECT 2836.330 1583.290 2837.510 1584.470 ;
        RECT 2837.930 1583.290 2839.110 1584.470 ;
        RECT 2836.330 1581.690 2837.510 1582.870 ;
        RECT 2837.930 1581.690 2839.110 1582.870 ;
        RECT 2836.330 1403.290 2837.510 1404.470 ;
        RECT 2837.930 1403.290 2839.110 1404.470 ;
        RECT 2836.330 1401.690 2837.510 1402.870 ;
        RECT 2837.930 1401.690 2839.110 1402.870 ;
        RECT 2836.330 1223.290 2837.510 1224.470 ;
        RECT 2837.930 1223.290 2839.110 1224.470 ;
        RECT 2836.330 1221.690 2837.510 1222.870 ;
        RECT 2837.930 1221.690 2839.110 1222.870 ;
        RECT 2836.330 1043.290 2837.510 1044.470 ;
        RECT 2837.930 1043.290 2839.110 1044.470 ;
        RECT 2836.330 1041.690 2837.510 1042.870 ;
        RECT 2837.930 1041.690 2839.110 1042.870 ;
        RECT 2836.330 863.290 2837.510 864.470 ;
        RECT 2837.930 863.290 2839.110 864.470 ;
        RECT 2836.330 861.690 2837.510 862.870 ;
        RECT 2837.930 861.690 2839.110 862.870 ;
        RECT 2836.330 683.290 2837.510 684.470 ;
        RECT 2837.930 683.290 2839.110 684.470 ;
        RECT 2836.330 681.690 2837.510 682.870 ;
        RECT 2837.930 681.690 2839.110 682.870 ;
        RECT 2836.330 503.290 2837.510 504.470 ;
        RECT 2837.930 503.290 2839.110 504.470 ;
        RECT 2836.330 501.690 2837.510 502.870 ;
        RECT 2837.930 501.690 2839.110 502.870 ;
        RECT 2836.330 323.290 2837.510 324.470 ;
        RECT 2837.930 323.290 2839.110 324.470 ;
        RECT 2836.330 321.690 2837.510 322.870 ;
        RECT 2837.930 321.690 2839.110 322.870 ;
        RECT 2836.330 143.290 2837.510 144.470 ;
        RECT 2837.930 143.290 2839.110 144.470 ;
        RECT 2836.330 141.690 2837.510 142.870 ;
        RECT 2837.930 141.690 2839.110 142.870 ;
        RECT 2836.330 -26.910 2837.510 -25.730 ;
        RECT 2837.930 -26.910 2839.110 -25.730 ;
        RECT 2836.330 -28.510 2837.510 -27.330 ;
        RECT 2837.930 -28.510 2839.110 -27.330 ;
        RECT 2950.710 3547.010 2951.890 3548.190 ;
        RECT 2952.310 3547.010 2953.490 3548.190 ;
        RECT 2950.710 3545.410 2951.890 3546.590 ;
        RECT 2952.310 3545.410 2953.490 3546.590 ;
        RECT 2950.710 3383.290 2951.890 3384.470 ;
        RECT 2952.310 3383.290 2953.490 3384.470 ;
        RECT 2950.710 3381.690 2951.890 3382.870 ;
        RECT 2952.310 3381.690 2953.490 3382.870 ;
        RECT 2950.710 3203.290 2951.890 3204.470 ;
        RECT 2952.310 3203.290 2953.490 3204.470 ;
        RECT 2950.710 3201.690 2951.890 3202.870 ;
        RECT 2952.310 3201.690 2953.490 3202.870 ;
        RECT 2950.710 3023.290 2951.890 3024.470 ;
        RECT 2952.310 3023.290 2953.490 3024.470 ;
        RECT 2950.710 3021.690 2951.890 3022.870 ;
        RECT 2952.310 3021.690 2953.490 3022.870 ;
        RECT 2950.710 2843.290 2951.890 2844.470 ;
        RECT 2952.310 2843.290 2953.490 2844.470 ;
        RECT 2950.710 2841.690 2951.890 2842.870 ;
        RECT 2952.310 2841.690 2953.490 2842.870 ;
        RECT 2950.710 2663.290 2951.890 2664.470 ;
        RECT 2952.310 2663.290 2953.490 2664.470 ;
        RECT 2950.710 2661.690 2951.890 2662.870 ;
        RECT 2952.310 2661.690 2953.490 2662.870 ;
        RECT 2950.710 2483.290 2951.890 2484.470 ;
        RECT 2952.310 2483.290 2953.490 2484.470 ;
        RECT 2950.710 2481.690 2951.890 2482.870 ;
        RECT 2952.310 2481.690 2953.490 2482.870 ;
        RECT 2950.710 2303.290 2951.890 2304.470 ;
        RECT 2952.310 2303.290 2953.490 2304.470 ;
        RECT 2950.710 2301.690 2951.890 2302.870 ;
        RECT 2952.310 2301.690 2953.490 2302.870 ;
        RECT 2950.710 2123.290 2951.890 2124.470 ;
        RECT 2952.310 2123.290 2953.490 2124.470 ;
        RECT 2950.710 2121.690 2951.890 2122.870 ;
        RECT 2952.310 2121.690 2953.490 2122.870 ;
        RECT 2950.710 1943.290 2951.890 1944.470 ;
        RECT 2952.310 1943.290 2953.490 1944.470 ;
        RECT 2950.710 1941.690 2951.890 1942.870 ;
        RECT 2952.310 1941.690 2953.490 1942.870 ;
        RECT 2950.710 1763.290 2951.890 1764.470 ;
        RECT 2952.310 1763.290 2953.490 1764.470 ;
        RECT 2950.710 1761.690 2951.890 1762.870 ;
        RECT 2952.310 1761.690 2953.490 1762.870 ;
        RECT 2950.710 1583.290 2951.890 1584.470 ;
        RECT 2952.310 1583.290 2953.490 1584.470 ;
        RECT 2950.710 1581.690 2951.890 1582.870 ;
        RECT 2952.310 1581.690 2953.490 1582.870 ;
        RECT 2950.710 1403.290 2951.890 1404.470 ;
        RECT 2952.310 1403.290 2953.490 1404.470 ;
        RECT 2950.710 1401.690 2951.890 1402.870 ;
        RECT 2952.310 1401.690 2953.490 1402.870 ;
        RECT 2950.710 1223.290 2951.890 1224.470 ;
        RECT 2952.310 1223.290 2953.490 1224.470 ;
        RECT 2950.710 1221.690 2951.890 1222.870 ;
        RECT 2952.310 1221.690 2953.490 1222.870 ;
        RECT 2950.710 1043.290 2951.890 1044.470 ;
        RECT 2952.310 1043.290 2953.490 1044.470 ;
        RECT 2950.710 1041.690 2951.890 1042.870 ;
        RECT 2952.310 1041.690 2953.490 1042.870 ;
        RECT 2950.710 863.290 2951.890 864.470 ;
        RECT 2952.310 863.290 2953.490 864.470 ;
        RECT 2950.710 861.690 2951.890 862.870 ;
        RECT 2952.310 861.690 2953.490 862.870 ;
        RECT 2950.710 683.290 2951.890 684.470 ;
        RECT 2952.310 683.290 2953.490 684.470 ;
        RECT 2950.710 681.690 2951.890 682.870 ;
        RECT 2952.310 681.690 2953.490 682.870 ;
        RECT 2950.710 503.290 2951.890 504.470 ;
        RECT 2952.310 503.290 2953.490 504.470 ;
        RECT 2950.710 501.690 2951.890 502.870 ;
        RECT 2952.310 501.690 2953.490 502.870 ;
        RECT 2950.710 323.290 2951.890 324.470 ;
        RECT 2952.310 323.290 2953.490 324.470 ;
        RECT 2950.710 321.690 2951.890 322.870 ;
        RECT 2952.310 321.690 2953.490 322.870 ;
        RECT 2950.710 143.290 2951.890 144.470 ;
        RECT 2952.310 143.290 2953.490 144.470 ;
        RECT 2950.710 141.690 2951.890 142.870 ;
        RECT 2952.310 141.690 2953.490 142.870 ;
        RECT 2950.710 -26.910 2951.890 -25.730 ;
        RECT 2952.310 -26.910 2953.490 -25.730 ;
        RECT 2950.710 -28.510 2951.890 -27.330 ;
        RECT 2952.310 -28.510 2953.490 -27.330 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
        RECT -34.030 861.530 2953.650 864.630 ;
        RECT -34.030 681.530 2953.650 684.630 ;
        RECT -34.030 501.530 2953.650 504.630 ;
        RECT -34.030 321.530 2953.650 324.630 ;
        RECT -34.030 141.530 2953.650 144.630 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
        RECT 334.770 1010.000 337.870 3557.950 ;
        RECT 514.770 1010.000 517.870 3557.950 ;
        RECT 694.770 1010.000 697.870 3557.950 ;
        RECT 874.770 1010.000 877.870 3557.950 ;
        RECT 1054.770 1010.000 1057.870 3557.950 ;
        RECT 334.770 -38.270 337.870 390.000 ;
        RECT 514.770 -38.270 517.870 390.000 ;
        RECT 694.770 -38.270 697.870 390.000 ;
        RECT 874.770 -38.270 877.870 390.000 ;
        RECT 1054.770 -38.270 1057.870 390.000 ;
        RECT 1234.770 -38.270 1237.870 3557.950 ;
        RECT 1414.770 -38.270 1417.870 3557.950 ;
        RECT 1594.770 -38.270 1597.870 3557.950 ;
        RECT 1774.770 -38.270 1777.870 3557.950 ;
        RECT 1954.770 -38.270 1957.870 3557.950 ;
        RECT 2134.770 -38.270 2137.870 3557.950 ;
        RECT 2314.770 -38.270 2317.870 3557.950 ;
        RECT 2494.770 -38.270 2497.870 3557.950 ;
        RECT 2674.770 -38.270 2677.870 3557.950 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER via4 ;
        RECT -43.470 3556.610 -42.290 3557.790 ;
        RECT -41.870 3556.610 -40.690 3557.790 ;
        RECT -43.470 3555.010 -42.290 3556.190 ;
        RECT -41.870 3555.010 -40.690 3556.190 ;
        RECT -43.470 3401.890 -42.290 3403.070 ;
        RECT -41.870 3401.890 -40.690 3403.070 ;
        RECT -43.470 3400.290 -42.290 3401.470 ;
        RECT -41.870 3400.290 -40.690 3401.470 ;
        RECT -43.470 3221.890 -42.290 3223.070 ;
        RECT -41.870 3221.890 -40.690 3223.070 ;
        RECT -43.470 3220.290 -42.290 3221.470 ;
        RECT -41.870 3220.290 -40.690 3221.470 ;
        RECT -43.470 3041.890 -42.290 3043.070 ;
        RECT -41.870 3041.890 -40.690 3043.070 ;
        RECT -43.470 3040.290 -42.290 3041.470 ;
        RECT -41.870 3040.290 -40.690 3041.470 ;
        RECT -43.470 2861.890 -42.290 2863.070 ;
        RECT -41.870 2861.890 -40.690 2863.070 ;
        RECT -43.470 2860.290 -42.290 2861.470 ;
        RECT -41.870 2860.290 -40.690 2861.470 ;
        RECT -43.470 2681.890 -42.290 2683.070 ;
        RECT -41.870 2681.890 -40.690 2683.070 ;
        RECT -43.470 2680.290 -42.290 2681.470 ;
        RECT -41.870 2680.290 -40.690 2681.470 ;
        RECT -43.470 2501.890 -42.290 2503.070 ;
        RECT -41.870 2501.890 -40.690 2503.070 ;
        RECT -43.470 2500.290 -42.290 2501.470 ;
        RECT -41.870 2500.290 -40.690 2501.470 ;
        RECT -43.470 2321.890 -42.290 2323.070 ;
        RECT -41.870 2321.890 -40.690 2323.070 ;
        RECT -43.470 2320.290 -42.290 2321.470 ;
        RECT -41.870 2320.290 -40.690 2321.470 ;
        RECT -43.470 2141.890 -42.290 2143.070 ;
        RECT -41.870 2141.890 -40.690 2143.070 ;
        RECT -43.470 2140.290 -42.290 2141.470 ;
        RECT -41.870 2140.290 -40.690 2141.470 ;
        RECT -43.470 1961.890 -42.290 1963.070 ;
        RECT -41.870 1961.890 -40.690 1963.070 ;
        RECT -43.470 1960.290 -42.290 1961.470 ;
        RECT -41.870 1960.290 -40.690 1961.470 ;
        RECT -43.470 1781.890 -42.290 1783.070 ;
        RECT -41.870 1781.890 -40.690 1783.070 ;
        RECT -43.470 1780.290 -42.290 1781.470 ;
        RECT -41.870 1780.290 -40.690 1781.470 ;
        RECT -43.470 1601.890 -42.290 1603.070 ;
        RECT -41.870 1601.890 -40.690 1603.070 ;
        RECT -43.470 1600.290 -42.290 1601.470 ;
        RECT -41.870 1600.290 -40.690 1601.470 ;
        RECT -43.470 1421.890 -42.290 1423.070 ;
        RECT -41.870 1421.890 -40.690 1423.070 ;
        RECT -43.470 1420.290 -42.290 1421.470 ;
        RECT -41.870 1420.290 -40.690 1421.470 ;
        RECT -43.470 1241.890 -42.290 1243.070 ;
        RECT -41.870 1241.890 -40.690 1243.070 ;
        RECT -43.470 1240.290 -42.290 1241.470 ;
        RECT -41.870 1240.290 -40.690 1241.470 ;
        RECT -43.470 1061.890 -42.290 1063.070 ;
        RECT -41.870 1061.890 -40.690 1063.070 ;
        RECT -43.470 1060.290 -42.290 1061.470 ;
        RECT -41.870 1060.290 -40.690 1061.470 ;
        RECT -43.470 881.890 -42.290 883.070 ;
        RECT -41.870 881.890 -40.690 883.070 ;
        RECT -43.470 880.290 -42.290 881.470 ;
        RECT -41.870 880.290 -40.690 881.470 ;
        RECT -43.470 701.890 -42.290 703.070 ;
        RECT -41.870 701.890 -40.690 703.070 ;
        RECT -43.470 700.290 -42.290 701.470 ;
        RECT -41.870 700.290 -40.690 701.470 ;
        RECT -43.470 521.890 -42.290 523.070 ;
        RECT -41.870 521.890 -40.690 523.070 ;
        RECT -43.470 520.290 -42.290 521.470 ;
        RECT -41.870 520.290 -40.690 521.470 ;
        RECT -43.470 341.890 -42.290 343.070 ;
        RECT -41.870 341.890 -40.690 343.070 ;
        RECT -43.470 340.290 -42.290 341.470 ;
        RECT -41.870 340.290 -40.690 341.470 ;
        RECT -43.470 161.890 -42.290 163.070 ;
        RECT -41.870 161.890 -40.690 163.070 ;
        RECT -43.470 160.290 -42.290 161.470 ;
        RECT -41.870 160.290 -40.690 161.470 ;
        RECT -43.470 -36.510 -42.290 -35.330 ;
        RECT -41.870 -36.510 -40.690 -35.330 ;
        RECT -43.470 -38.110 -42.290 -36.930 ;
        RECT -41.870 -38.110 -40.690 -36.930 ;
        RECT 154.930 3556.610 156.110 3557.790 ;
        RECT 156.530 3556.610 157.710 3557.790 ;
        RECT 154.930 3555.010 156.110 3556.190 ;
        RECT 156.530 3555.010 157.710 3556.190 ;
        RECT 154.930 3401.890 156.110 3403.070 ;
        RECT 156.530 3401.890 157.710 3403.070 ;
        RECT 154.930 3400.290 156.110 3401.470 ;
        RECT 156.530 3400.290 157.710 3401.470 ;
        RECT 154.930 3221.890 156.110 3223.070 ;
        RECT 156.530 3221.890 157.710 3223.070 ;
        RECT 154.930 3220.290 156.110 3221.470 ;
        RECT 156.530 3220.290 157.710 3221.470 ;
        RECT 154.930 3041.890 156.110 3043.070 ;
        RECT 156.530 3041.890 157.710 3043.070 ;
        RECT 154.930 3040.290 156.110 3041.470 ;
        RECT 156.530 3040.290 157.710 3041.470 ;
        RECT 154.930 2861.890 156.110 2863.070 ;
        RECT 156.530 2861.890 157.710 2863.070 ;
        RECT 154.930 2860.290 156.110 2861.470 ;
        RECT 156.530 2860.290 157.710 2861.470 ;
        RECT 154.930 2681.890 156.110 2683.070 ;
        RECT 156.530 2681.890 157.710 2683.070 ;
        RECT 154.930 2680.290 156.110 2681.470 ;
        RECT 156.530 2680.290 157.710 2681.470 ;
        RECT 154.930 2501.890 156.110 2503.070 ;
        RECT 156.530 2501.890 157.710 2503.070 ;
        RECT 154.930 2500.290 156.110 2501.470 ;
        RECT 156.530 2500.290 157.710 2501.470 ;
        RECT 154.930 2321.890 156.110 2323.070 ;
        RECT 156.530 2321.890 157.710 2323.070 ;
        RECT 154.930 2320.290 156.110 2321.470 ;
        RECT 156.530 2320.290 157.710 2321.470 ;
        RECT 154.930 2141.890 156.110 2143.070 ;
        RECT 156.530 2141.890 157.710 2143.070 ;
        RECT 154.930 2140.290 156.110 2141.470 ;
        RECT 156.530 2140.290 157.710 2141.470 ;
        RECT 154.930 1961.890 156.110 1963.070 ;
        RECT 156.530 1961.890 157.710 1963.070 ;
        RECT 154.930 1960.290 156.110 1961.470 ;
        RECT 156.530 1960.290 157.710 1961.470 ;
        RECT 154.930 1781.890 156.110 1783.070 ;
        RECT 156.530 1781.890 157.710 1783.070 ;
        RECT 154.930 1780.290 156.110 1781.470 ;
        RECT 156.530 1780.290 157.710 1781.470 ;
        RECT 154.930 1601.890 156.110 1603.070 ;
        RECT 156.530 1601.890 157.710 1603.070 ;
        RECT 154.930 1600.290 156.110 1601.470 ;
        RECT 156.530 1600.290 157.710 1601.470 ;
        RECT 154.930 1421.890 156.110 1423.070 ;
        RECT 156.530 1421.890 157.710 1423.070 ;
        RECT 154.930 1420.290 156.110 1421.470 ;
        RECT 156.530 1420.290 157.710 1421.470 ;
        RECT 154.930 1241.890 156.110 1243.070 ;
        RECT 156.530 1241.890 157.710 1243.070 ;
        RECT 154.930 1240.290 156.110 1241.470 ;
        RECT 156.530 1240.290 157.710 1241.470 ;
        RECT 154.930 1061.890 156.110 1063.070 ;
        RECT 156.530 1061.890 157.710 1063.070 ;
        RECT 154.930 1060.290 156.110 1061.470 ;
        RECT 156.530 1060.290 157.710 1061.470 ;
        RECT 334.930 3556.610 336.110 3557.790 ;
        RECT 336.530 3556.610 337.710 3557.790 ;
        RECT 334.930 3555.010 336.110 3556.190 ;
        RECT 336.530 3555.010 337.710 3556.190 ;
        RECT 334.930 3401.890 336.110 3403.070 ;
        RECT 336.530 3401.890 337.710 3403.070 ;
        RECT 334.930 3400.290 336.110 3401.470 ;
        RECT 336.530 3400.290 337.710 3401.470 ;
        RECT 334.930 3221.890 336.110 3223.070 ;
        RECT 336.530 3221.890 337.710 3223.070 ;
        RECT 334.930 3220.290 336.110 3221.470 ;
        RECT 336.530 3220.290 337.710 3221.470 ;
        RECT 334.930 3041.890 336.110 3043.070 ;
        RECT 336.530 3041.890 337.710 3043.070 ;
        RECT 334.930 3040.290 336.110 3041.470 ;
        RECT 336.530 3040.290 337.710 3041.470 ;
        RECT 334.930 2861.890 336.110 2863.070 ;
        RECT 336.530 2861.890 337.710 2863.070 ;
        RECT 334.930 2860.290 336.110 2861.470 ;
        RECT 336.530 2860.290 337.710 2861.470 ;
        RECT 334.930 2681.890 336.110 2683.070 ;
        RECT 336.530 2681.890 337.710 2683.070 ;
        RECT 334.930 2680.290 336.110 2681.470 ;
        RECT 336.530 2680.290 337.710 2681.470 ;
        RECT 334.930 2501.890 336.110 2503.070 ;
        RECT 336.530 2501.890 337.710 2503.070 ;
        RECT 334.930 2500.290 336.110 2501.470 ;
        RECT 336.530 2500.290 337.710 2501.470 ;
        RECT 334.930 2321.890 336.110 2323.070 ;
        RECT 336.530 2321.890 337.710 2323.070 ;
        RECT 334.930 2320.290 336.110 2321.470 ;
        RECT 336.530 2320.290 337.710 2321.470 ;
        RECT 334.930 2141.890 336.110 2143.070 ;
        RECT 336.530 2141.890 337.710 2143.070 ;
        RECT 334.930 2140.290 336.110 2141.470 ;
        RECT 336.530 2140.290 337.710 2141.470 ;
        RECT 334.930 1961.890 336.110 1963.070 ;
        RECT 336.530 1961.890 337.710 1963.070 ;
        RECT 334.930 1960.290 336.110 1961.470 ;
        RECT 336.530 1960.290 337.710 1961.470 ;
        RECT 334.930 1781.890 336.110 1783.070 ;
        RECT 336.530 1781.890 337.710 1783.070 ;
        RECT 334.930 1780.290 336.110 1781.470 ;
        RECT 336.530 1780.290 337.710 1781.470 ;
        RECT 334.930 1601.890 336.110 1603.070 ;
        RECT 336.530 1601.890 337.710 1603.070 ;
        RECT 334.930 1600.290 336.110 1601.470 ;
        RECT 336.530 1600.290 337.710 1601.470 ;
        RECT 334.930 1421.890 336.110 1423.070 ;
        RECT 336.530 1421.890 337.710 1423.070 ;
        RECT 334.930 1420.290 336.110 1421.470 ;
        RECT 336.530 1420.290 337.710 1421.470 ;
        RECT 334.930 1241.890 336.110 1243.070 ;
        RECT 336.530 1241.890 337.710 1243.070 ;
        RECT 334.930 1240.290 336.110 1241.470 ;
        RECT 336.530 1240.290 337.710 1241.470 ;
        RECT 334.930 1061.890 336.110 1063.070 ;
        RECT 336.530 1061.890 337.710 1063.070 ;
        RECT 334.930 1060.290 336.110 1061.470 ;
        RECT 336.530 1060.290 337.710 1061.470 ;
        RECT 514.930 3556.610 516.110 3557.790 ;
        RECT 516.530 3556.610 517.710 3557.790 ;
        RECT 514.930 3555.010 516.110 3556.190 ;
        RECT 516.530 3555.010 517.710 3556.190 ;
        RECT 514.930 3401.890 516.110 3403.070 ;
        RECT 516.530 3401.890 517.710 3403.070 ;
        RECT 514.930 3400.290 516.110 3401.470 ;
        RECT 516.530 3400.290 517.710 3401.470 ;
        RECT 514.930 3221.890 516.110 3223.070 ;
        RECT 516.530 3221.890 517.710 3223.070 ;
        RECT 514.930 3220.290 516.110 3221.470 ;
        RECT 516.530 3220.290 517.710 3221.470 ;
        RECT 514.930 3041.890 516.110 3043.070 ;
        RECT 516.530 3041.890 517.710 3043.070 ;
        RECT 514.930 3040.290 516.110 3041.470 ;
        RECT 516.530 3040.290 517.710 3041.470 ;
        RECT 514.930 2861.890 516.110 2863.070 ;
        RECT 516.530 2861.890 517.710 2863.070 ;
        RECT 514.930 2860.290 516.110 2861.470 ;
        RECT 516.530 2860.290 517.710 2861.470 ;
        RECT 514.930 2681.890 516.110 2683.070 ;
        RECT 516.530 2681.890 517.710 2683.070 ;
        RECT 514.930 2680.290 516.110 2681.470 ;
        RECT 516.530 2680.290 517.710 2681.470 ;
        RECT 514.930 2501.890 516.110 2503.070 ;
        RECT 516.530 2501.890 517.710 2503.070 ;
        RECT 514.930 2500.290 516.110 2501.470 ;
        RECT 516.530 2500.290 517.710 2501.470 ;
        RECT 514.930 2321.890 516.110 2323.070 ;
        RECT 516.530 2321.890 517.710 2323.070 ;
        RECT 514.930 2320.290 516.110 2321.470 ;
        RECT 516.530 2320.290 517.710 2321.470 ;
        RECT 514.930 2141.890 516.110 2143.070 ;
        RECT 516.530 2141.890 517.710 2143.070 ;
        RECT 514.930 2140.290 516.110 2141.470 ;
        RECT 516.530 2140.290 517.710 2141.470 ;
        RECT 514.930 1961.890 516.110 1963.070 ;
        RECT 516.530 1961.890 517.710 1963.070 ;
        RECT 514.930 1960.290 516.110 1961.470 ;
        RECT 516.530 1960.290 517.710 1961.470 ;
        RECT 514.930 1781.890 516.110 1783.070 ;
        RECT 516.530 1781.890 517.710 1783.070 ;
        RECT 514.930 1780.290 516.110 1781.470 ;
        RECT 516.530 1780.290 517.710 1781.470 ;
        RECT 514.930 1601.890 516.110 1603.070 ;
        RECT 516.530 1601.890 517.710 1603.070 ;
        RECT 514.930 1600.290 516.110 1601.470 ;
        RECT 516.530 1600.290 517.710 1601.470 ;
        RECT 514.930 1421.890 516.110 1423.070 ;
        RECT 516.530 1421.890 517.710 1423.070 ;
        RECT 514.930 1420.290 516.110 1421.470 ;
        RECT 516.530 1420.290 517.710 1421.470 ;
        RECT 514.930 1241.890 516.110 1243.070 ;
        RECT 516.530 1241.890 517.710 1243.070 ;
        RECT 514.930 1240.290 516.110 1241.470 ;
        RECT 516.530 1240.290 517.710 1241.470 ;
        RECT 514.930 1061.890 516.110 1063.070 ;
        RECT 516.530 1061.890 517.710 1063.070 ;
        RECT 514.930 1060.290 516.110 1061.470 ;
        RECT 516.530 1060.290 517.710 1061.470 ;
        RECT 694.930 3556.610 696.110 3557.790 ;
        RECT 696.530 3556.610 697.710 3557.790 ;
        RECT 694.930 3555.010 696.110 3556.190 ;
        RECT 696.530 3555.010 697.710 3556.190 ;
        RECT 694.930 3401.890 696.110 3403.070 ;
        RECT 696.530 3401.890 697.710 3403.070 ;
        RECT 694.930 3400.290 696.110 3401.470 ;
        RECT 696.530 3400.290 697.710 3401.470 ;
        RECT 694.930 3221.890 696.110 3223.070 ;
        RECT 696.530 3221.890 697.710 3223.070 ;
        RECT 694.930 3220.290 696.110 3221.470 ;
        RECT 696.530 3220.290 697.710 3221.470 ;
        RECT 694.930 3041.890 696.110 3043.070 ;
        RECT 696.530 3041.890 697.710 3043.070 ;
        RECT 694.930 3040.290 696.110 3041.470 ;
        RECT 696.530 3040.290 697.710 3041.470 ;
        RECT 694.930 2861.890 696.110 2863.070 ;
        RECT 696.530 2861.890 697.710 2863.070 ;
        RECT 694.930 2860.290 696.110 2861.470 ;
        RECT 696.530 2860.290 697.710 2861.470 ;
        RECT 694.930 2681.890 696.110 2683.070 ;
        RECT 696.530 2681.890 697.710 2683.070 ;
        RECT 694.930 2680.290 696.110 2681.470 ;
        RECT 696.530 2680.290 697.710 2681.470 ;
        RECT 694.930 2501.890 696.110 2503.070 ;
        RECT 696.530 2501.890 697.710 2503.070 ;
        RECT 694.930 2500.290 696.110 2501.470 ;
        RECT 696.530 2500.290 697.710 2501.470 ;
        RECT 694.930 2321.890 696.110 2323.070 ;
        RECT 696.530 2321.890 697.710 2323.070 ;
        RECT 694.930 2320.290 696.110 2321.470 ;
        RECT 696.530 2320.290 697.710 2321.470 ;
        RECT 694.930 2141.890 696.110 2143.070 ;
        RECT 696.530 2141.890 697.710 2143.070 ;
        RECT 694.930 2140.290 696.110 2141.470 ;
        RECT 696.530 2140.290 697.710 2141.470 ;
        RECT 694.930 1961.890 696.110 1963.070 ;
        RECT 696.530 1961.890 697.710 1963.070 ;
        RECT 694.930 1960.290 696.110 1961.470 ;
        RECT 696.530 1960.290 697.710 1961.470 ;
        RECT 694.930 1781.890 696.110 1783.070 ;
        RECT 696.530 1781.890 697.710 1783.070 ;
        RECT 694.930 1780.290 696.110 1781.470 ;
        RECT 696.530 1780.290 697.710 1781.470 ;
        RECT 694.930 1601.890 696.110 1603.070 ;
        RECT 696.530 1601.890 697.710 1603.070 ;
        RECT 694.930 1600.290 696.110 1601.470 ;
        RECT 696.530 1600.290 697.710 1601.470 ;
        RECT 694.930 1421.890 696.110 1423.070 ;
        RECT 696.530 1421.890 697.710 1423.070 ;
        RECT 694.930 1420.290 696.110 1421.470 ;
        RECT 696.530 1420.290 697.710 1421.470 ;
        RECT 694.930 1241.890 696.110 1243.070 ;
        RECT 696.530 1241.890 697.710 1243.070 ;
        RECT 694.930 1240.290 696.110 1241.470 ;
        RECT 696.530 1240.290 697.710 1241.470 ;
        RECT 694.930 1061.890 696.110 1063.070 ;
        RECT 696.530 1061.890 697.710 1063.070 ;
        RECT 694.930 1060.290 696.110 1061.470 ;
        RECT 696.530 1060.290 697.710 1061.470 ;
        RECT 874.930 3556.610 876.110 3557.790 ;
        RECT 876.530 3556.610 877.710 3557.790 ;
        RECT 874.930 3555.010 876.110 3556.190 ;
        RECT 876.530 3555.010 877.710 3556.190 ;
        RECT 874.930 3401.890 876.110 3403.070 ;
        RECT 876.530 3401.890 877.710 3403.070 ;
        RECT 874.930 3400.290 876.110 3401.470 ;
        RECT 876.530 3400.290 877.710 3401.470 ;
        RECT 874.930 3221.890 876.110 3223.070 ;
        RECT 876.530 3221.890 877.710 3223.070 ;
        RECT 874.930 3220.290 876.110 3221.470 ;
        RECT 876.530 3220.290 877.710 3221.470 ;
        RECT 874.930 3041.890 876.110 3043.070 ;
        RECT 876.530 3041.890 877.710 3043.070 ;
        RECT 874.930 3040.290 876.110 3041.470 ;
        RECT 876.530 3040.290 877.710 3041.470 ;
        RECT 874.930 2861.890 876.110 2863.070 ;
        RECT 876.530 2861.890 877.710 2863.070 ;
        RECT 874.930 2860.290 876.110 2861.470 ;
        RECT 876.530 2860.290 877.710 2861.470 ;
        RECT 874.930 2681.890 876.110 2683.070 ;
        RECT 876.530 2681.890 877.710 2683.070 ;
        RECT 874.930 2680.290 876.110 2681.470 ;
        RECT 876.530 2680.290 877.710 2681.470 ;
        RECT 874.930 2501.890 876.110 2503.070 ;
        RECT 876.530 2501.890 877.710 2503.070 ;
        RECT 874.930 2500.290 876.110 2501.470 ;
        RECT 876.530 2500.290 877.710 2501.470 ;
        RECT 874.930 2321.890 876.110 2323.070 ;
        RECT 876.530 2321.890 877.710 2323.070 ;
        RECT 874.930 2320.290 876.110 2321.470 ;
        RECT 876.530 2320.290 877.710 2321.470 ;
        RECT 874.930 2141.890 876.110 2143.070 ;
        RECT 876.530 2141.890 877.710 2143.070 ;
        RECT 874.930 2140.290 876.110 2141.470 ;
        RECT 876.530 2140.290 877.710 2141.470 ;
        RECT 874.930 1961.890 876.110 1963.070 ;
        RECT 876.530 1961.890 877.710 1963.070 ;
        RECT 874.930 1960.290 876.110 1961.470 ;
        RECT 876.530 1960.290 877.710 1961.470 ;
        RECT 874.930 1781.890 876.110 1783.070 ;
        RECT 876.530 1781.890 877.710 1783.070 ;
        RECT 874.930 1780.290 876.110 1781.470 ;
        RECT 876.530 1780.290 877.710 1781.470 ;
        RECT 874.930 1601.890 876.110 1603.070 ;
        RECT 876.530 1601.890 877.710 1603.070 ;
        RECT 874.930 1600.290 876.110 1601.470 ;
        RECT 876.530 1600.290 877.710 1601.470 ;
        RECT 874.930 1421.890 876.110 1423.070 ;
        RECT 876.530 1421.890 877.710 1423.070 ;
        RECT 874.930 1420.290 876.110 1421.470 ;
        RECT 876.530 1420.290 877.710 1421.470 ;
        RECT 874.930 1241.890 876.110 1243.070 ;
        RECT 876.530 1241.890 877.710 1243.070 ;
        RECT 874.930 1240.290 876.110 1241.470 ;
        RECT 876.530 1240.290 877.710 1241.470 ;
        RECT 874.930 1061.890 876.110 1063.070 ;
        RECT 876.530 1061.890 877.710 1063.070 ;
        RECT 874.930 1060.290 876.110 1061.470 ;
        RECT 876.530 1060.290 877.710 1061.470 ;
        RECT 1054.930 3556.610 1056.110 3557.790 ;
        RECT 1056.530 3556.610 1057.710 3557.790 ;
        RECT 1054.930 3555.010 1056.110 3556.190 ;
        RECT 1056.530 3555.010 1057.710 3556.190 ;
        RECT 1054.930 3401.890 1056.110 3403.070 ;
        RECT 1056.530 3401.890 1057.710 3403.070 ;
        RECT 1054.930 3400.290 1056.110 3401.470 ;
        RECT 1056.530 3400.290 1057.710 3401.470 ;
        RECT 1054.930 3221.890 1056.110 3223.070 ;
        RECT 1056.530 3221.890 1057.710 3223.070 ;
        RECT 1054.930 3220.290 1056.110 3221.470 ;
        RECT 1056.530 3220.290 1057.710 3221.470 ;
        RECT 1054.930 3041.890 1056.110 3043.070 ;
        RECT 1056.530 3041.890 1057.710 3043.070 ;
        RECT 1054.930 3040.290 1056.110 3041.470 ;
        RECT 1056.530 3040.290 1057.710 3041.470 ;
        RECT 1054.930 2861.890 1056.110 2863.070 ;
        RECT 1056.530 2861.890 1057.710 2863.070 ;
        RECT 1054.930 2860.290 1056.110 2861.470 ;
        RECT 1056.530 2860.290 1057.710 2861.470 ;
        RECT 1054.930 2681.890 1056.110 2683.070 ;
        RECT 1056.530 2681.890 1057.710 2683.070 ;
        RECT 1054.930 2680.290 1056.110 2681.470 ;
        RECT 1056.530 2680.290 1057.710 2681.470 ;
        RECT 1054.930 2501.890 1056.110 2503.070 ;
        RECT 1056.530 2501.890 1057.710 2503.070 ;
        RECT 1054.930 2500.290 1056.110 2501.470 ;
        RECT 1056.530 2500.290 1057.710 2501.470 ;
        RECT 1054.930 2321.890 1056.110 2323.070 ;
        RECT 1056.530 2321.890 1057.710 2323.070 ;
        RECT 1054.930 2320.290 1056.110 2321.470 ;
        RECT 1056.530 2320.290 1057.710 2321.470 ;
        RECT 1054.930 2141.890 1056.110 2143.070 ;
        RECT 1056.530 2141.890 1057.710 2143.070 ;
        RECT 1054.930 2140.290 1056.110 2141.470 ;
        RECT 1056.530 2140.290 1057.710 2141.470 ;
        RECT 1054.930 1961.890 1056.110 1963.070 ;
        RECT 1056.530 1961.890 1057.710 1963.070 ;
        RECT 1054.930 1960.290 1056.110 1961.470 ;
        RECT 1056.530 1960.290 1057.710 1961.470 ;
        RECT 1054.930 1781.890 1056.110 1783.070 ;
        RECT 1056.530 1781.890 1057.710 1783.070 ;
        RECT 1054.930 1780.290 1056.110 1781.470 ;
        RECT 1056.530 1780.290 1057.710 1781.470 ;
        RECT 1054.930 1601.890 1056.110 1603.070 ;
        RECT 1056.530 1601.890 1057.710 1603.070 ;
        RECT 1054.930 1600.290 1056.110 1601.470 ;
        RECT 1056.530 1600.290 1057.710 1601.470 ;
        RECT 1054.930 1421.890 1056.110 1423.070 ;
        RECT 1056.530 1421.890 1057.710 1423.070 ;
        RECT 1054.930 1420.290 1056.110 1421.470 ;
        RECT 1056.530 1420.290 1057.710 1421.470 ;
        RECT 1054.930 1241.890 1056.110 1243.070 ;
        RECT 1056.530 1241.890 1057.710 1243.070 ;
        RECT 1054.930 1240.290 1056.110 1241.470 ;
        RECT 1056.530 1240.290 1057.710 1241.470 ;
        RECT 1054.930 1061.890 1056.110 1063.070 ;
        RECT 1056.530 1061.890 1057.710 1063.070 ;
        RECT 1054.930 1060.290 1056.110 1061.470 ;
        RECT 1056.530 1060.290 1057.710 1061.470 ;
        RECT 1234.930 3556.610 1236.110 3557.790 ;
        RECT 1236.530 3556.610 1237.710 3557.790 ;
        RECT 1234.930 3555.010 1236.110 3556.190 ;
        RECT 1236.530 3555.010 1237.710 3556.190 ;
        RECT 1234.930 3401.890 1236.110 3403.070 ;
        RECT 1236.530 3401.890 1237.710 3403.070 ;
        RECT 1234.930 3400.290 1236.110 3401.470 ;
        RECT 1236.530 3400.290 1237.710 3401.470 ;
        RECT 1234.930 3221.890 1236.110 3223.070 ;
        RECT 1236.530 3221.890 1237.710 3223.070 ;
        RECT 1234.930 3220.290 1236.110 3221.470 ;
        RECT 1236.530 3220.290 1237.710 3221.470 ;
        RECT 1234.930 3041.890 1236.110 3043.070 ;
        RECT 1236.530 3041.890 1237.710 3043.070 ;
        RECT 1234.930 3040.290 1236.110 3041.470 ;
        RECT 1236.530 3040.290 1237.710 3041.470 ;
        RECT 1234.930 2861.890 1236.110 2863.070 ;
        RECT 1236.530 2861.890 1237.710 2863.070 ;
        RECT 1234.930 2860.290 1236.110 2861.470 ;
        RECT 1236.530 2860.290 1237.710 2861.470 ;
        RECT 1234.930 2681.890 1236.110 2683.070 ;
        RECT 1236.530 2681.890 1237.710 2683.070 ;
        RECT 1234.930 2680.290 1236.110 2681.470 ;
        RECT 1236.530 2680.290 1237.710 2681.470 ;
        RECT 1234.930 2501.890 1236.110 2503.070 ;
        RECT 1236.530 2501.890 1237.710 2503.070 ;
        RECT 1234.930 2500.290 1236.110 2501.470 ;
        RECT 1236.530 2500.290 1237.710 2501.470 ;
        RECT 1234.930 2321.890 1236.110 2323.070 ;
        RECT 1236.530 2321.890 1237.710 2323.070 ;
        RECT 1234.930 2320.290 1236.110 2321.470 ;
        RECT 1236.530 2320.290 1237.710 2321.470 ;
        RECT 1234.930 2141.890 1236.110 2143.070 ;
        RECT 1236.530 2141.890 1237.710 2143.070 ;
        RECT 1234.930 2140.290 1236.110 2141.470 ;
        RECT 1236.530 2140.290 1237.710 2141.470 ;
        RECT 1234.930 1961.890 1236.110 1963.070 ;
        RECT 1236.530 1961.890 1237.710 1963.070 ;
        RECT 1234.930 1960.290 1236.110 1961.470 ;
        RECT 1236.530 1960.290 1237.710 1961.470 ;
        RECT 1234.930 1781.890 1236.110 1783.070 ;
        RECT 1236.530 1781.890 1237.710 1783.070 ;
        RECT 1234.930 1780.290 1236.110 1781.470 ;
        RECT 1236.530 1780.290 1237.710 1781.470 ;
        RECT 1234.930 1601.890 1236.110 1603.070 ;
        RECT 1236.530 1601.890 1237.710 1603.070 ;
        RECT 1234.930 1600.290 1236.110 1601.470 ;
        RECT 1236.530 1600.290 1237.710 1601.470 ;
        RECT 1234.930 1421.890 1236.110 1423.070 ;
        RECT 1236.530 1421.890 1237.710 1423.070 ;
        RECT 1234.930 1420.290 1236.110 1421.470 ;
        RECT 1236.530 1420.290 1237.710 1421.470 ;
        RECT 1234.930 1241.890 1236.110 1243.070 ;
        RECT 1236.530 1241.890 1237.710 1243.070 ;
        RECT 1234.930 1240.290 1236.110 1241.470 ;
        RECT 1236.530 1240.290 1237.710 1241.470 ;
        RECT 1234.930 1061.890 1236.110 1063.070 ;
        RECT 1236.530 1061.890 1237.710 1063.070 ;
        RECT 1234.930 1060.290 1236.110 1061.470 ;
        RECT 1236.530 1060.290 1237.710 1061.470 ;
        RECT 154.930 881.890 156.110 883.070 ;
        RECT 156.530 881.890 157.710 883.070 ;
        RECT 154.930 880.290 156.110 881.470 ;
        RECT 156.530 880.290 157.710 881.470 ;
        RECT 154.930 701.890 156.110 703.070 ;
        RECT 156.530 701.890 157.710 703.070 ;
        RECT 154.930 700.290 156.110 701.470 ;
        RECT 156.530 700.290 157.710 701.470 ;
        RECT 154.930 521.890 156.110 523.070 ;
        RECT 156.530 521.890 157.710 523.070 ;
        RECT 154.930 520.290 156.110 521.470 ;
        RECT 156.530 520.290 157.710 521.470 ;
        RECT 1234.930 881.890 1236.110 883.070 ;
        RECT 1236.530 881.890 1237.710 883.070 ;
        RECT 1234.930 880.290 1236.110 881.470 ;
        RECT 1236.530 880.290 1237.710 881.470 ;
        RECT 1234.930 701.890 1236.110 703.070 ;
        RECT 1236.530 701.890 1237.710 703.070 ;
        RECT 1234.930 700.290 1236.110 701.470 ;
        RECT 1236.530 700.290 1237.710 701.470 ;
        RECT 1234.930 521.890 1236.110 523.070 ;
        RECT 1236.530 521.890 1237.710 523.070 ;
        RECT 1234.930 520.290 1236.110 521.470 ;
        RECT 1236.530 520.290 1237.710 521.470 ;
        RECT 154.930 341.890 156.110 343.070 ;
        RECT 156.530 341.890 157.710 343.070 ;
        RECT 154.930 340.290 156.110 341.470 ;
        RECT 156.530 340.290 157.710 341.470 ;
        RECT 154.930 161.890 156.110 163.070 ;
        RECT 156.530 161.890 157.710 163.070 ;
        RECT 154.930 160.290 156.110 161.470 ;
        RECT 156.530 160.290 157.710 161.470 ;
        RECT 154.930 -36.510 156.110 -35.330 ;
        RECT 156.530 -36.510 157.710 -35.330 ;
        RECT 154.930 -38.110 156.110 -36.930 ;
        RECT 156.530 -38.110 157.710 -36.930 ;
        RECT 334.930 341.890 336.110 343.070 ;
        RECT 336.530 341.890 337.710 343.070 ;
        RECT 334.930 340.290 336.110 341.470 ;
        RECT 336.530 340.290 337.710 341.470 ;
        RECT 334.930 161.890 336.110 163.070 ;
        RECT 336.530 161.890 337.710 163.070 ;
        RECT 334.930 160.290 336.110 161.470 ;
        RECT 336.530 160.290 337.710 161.470 ;
        RECT 334.930 -36.510 336.110 -35.330 ;
        RECT 336.530 -36.510 337.710 -35.330 ;
        RECT 334.930 -38.110 336.110 -36.930 ;
        RECT 336.530 -38.110 337.710 -36.930 ;
        RECT 514.930 341.890 516.110 343.070 ;
        RECT 516.530 341.890 517.710 343.070 ;
        RECT 514.930 340.290 516.110 341.470 ;
        RECT 516.530 340.290 517.710 341.470 ;
        RECT 514.930 161.890 516.110 163.070 ;
        RECT 516.530 161.890 517.710 163.070 ;
        RECT 514.930 160.290 516.110 161.470 ;
        RECT 516.530 160.290 517.710 161.470 ;
        RECT 514.930 -36.510 516.110 -35.330 ;
        RECT 516.530 -36.510 517.710 -35.330 ;
        RECT 514.930 -38.110 516.110 -36.930 ;
        RECT 516.530 -38.110 517.710 -36.930 ;
        RECT 694.930 341.890 696.110 343.070 ;
        RECT 696.530 341.890 697.710 343.070 ;
        RECT 694.930 340.290 696.110 341.470 ;
        RECT 696.530 340.290 697.710 341.470 ;
        RECT 694.930 161.890 696.110 163.070 ;
        RECT 696.530 161.890 697.710 163.070 ;
        RECT 694.930 160.290 696.110 161.470 ;
        RECT 696.530 160.290 697.710 161.470 ;
        RECT 694.930 -36.510 696.110 -35.330 ;
        RECT 696.530 -36.510 697.710 -35.330 ;
        RECT 694.930 -38.110 696.110 -36.930 ;
        RECT 696.530 -38.110 697.710 -36.930 ;
        RECT 874.930 341.890 876.110 343.070 ;
        RECT 876.530 341.890 877.710 343.070 ;
        RECT 874.930 340.290 876.110 341.470 ;
        RECT 876.530 340.290 877.710 341.470 ;
        RECT 874.930 161.890 876.110 163.070 ;
        RECT 876.530 161.890 877.710 163.070 ;
        RECT 874.930 160.290 876.110 161.470 ;
        RECT 876.530 160.290 877.710 161.470 ;
        RECT 874.930 -36.510 876.110 -35.330 ;
        RECT 876.530 -36.510 877.710 -35.330 ;
        RECT 874.930 -38.110 876.110 -36.930 ;
        RECT 876.530 -38.110 877.710 -36.930 ;
        RECT 1054.930 341.890 1056.110 343.070 ;
        RECT 1056.530 341.890 1057.710 343.070 ;
        RECT 1054.930 340.290 1056.110 341.470 ;
        RECT 1056.530 340.290 1057.710 341.470 ;
        RECT 1054.930 161.890 1056.110 163.070 ;
        RECT 1056.530 161.890 1057.710 163.070 ;
        RECT 1054.930 160.290 1056.110 161.470 ;
        RECT 1056.530 160.290 1057.710 161.470 ;
        RECT 1054.930 -36.510 1056.110 -35.330 ;
        RECT 1056.530 -36.510 1057.710 -35.330 ;
        RECT 1054.930 -38.110 1056.110 -36.930 ;
        RECT 1056.530 -38.110 1057.710 -36.930 ;
        RECT 1234.930 341.890 1236.110 343.070 ;
        RECT 1236.530 341.890 1237.710 343.070 ;
        RECT 1234.930 340.290 1236.110 341.470 ;
        RECT 1236.530 340.290 1237.710 341.470 ;
        RECT 1234.930 161.890 1236.110 163.070 ;
        RECT 1236.530 161.890 1237.710 163.070 ;
        RECT 1234.930 160.290 1236.110 161.470 ;
        RECT 1236.530 160.290 1237.710 161.470 ;
        RECT 1234.930 -36.510 1236.110 -35.330 ;
        RECT 1236.530 -36.510 1237.710 -35.330 ;
        RECT 1234.930 -38.110 1236.110 -36.930 ;
        RECT 1236.530 -38.110 1237.710 -36.930 ;
        RECT 1414.930 3556.610 1416.110 3557.790 ;
        RECT 1416.530 3556.610 1417.710 3557.790 ;
        RECT 1414.930 3555.010 1416.110 3556.190 ;
        RECT 1416.530 3555.010 1417.710 3556.190 ;
        RECT 1414.930 3401.890 1416.110 3403.070 ;
        RECT 1416.530 3401.890 1417.710 3403.070 ;
        RECT 1414.930 3400.290 1416.110 3401.470 ;
        RECT 1416.530 3400.290 1417.710 3401.470 ;
        RECT 1414.930 3221.890 1416.110 3223.070 ;
        RECT 1416.530 3221.890 1417.710 3223.070 ;
        RECT 1414.930 3220.290 1416.110 3221.470 ;
        RECT 1416.530 3220.290 1417.710 3221.470 ;
        RECT 1414.930 3041.890 1416.110 3043.070 ;
        RECT 1416.530 3041.890 1417.710 3043.070 ;
        RECT 1414.930 3040.290 1416.110 3041.470 ;
        RECT 1416.530 3040.290 1417.710 3041.470 ;
        RECT 1414.930 2861.890 1416.110 2863.070 ;
        RECT 1416.530 2861.890 1417.710 2863.070 ;
        RECT 1414.930 2860.290 1416.110 2861.470 ;
        RECT 1416.530 2860.290 1417.710 2861.470 ;
        RECT 1414.930 2681.890 1416.110 2683.070 ;
        RECT 1416.530 2681.890 1417.710 2683.070 ;
        RECT 1414.930 2680.290 1416.110 2681.470 ;
        RECT 1416.530 2680.290 1417.710 2681.470 ;
        RECT 1414.930 2501.890 1416.110 2503.070 ;
        RECT 1416.530 2501.890 1417.710 2503.070 ;
        RECT 1414.930 2500.290 1416.110 2501.470 ;
        RECT 1416.530 2500.290 1417.710 2501.470 ;
        RECT 1414.930 2321.890 1416.110 2323.070 ;
        RECT 1416.530 2321.890 1417.710 2323.070 ;
        RECT 1414.930 2320.290 1416.110 2321.470 ;
        RECT 1416.530 2320.290 1417.710 2321.470 ;
        RECT 1414.930 2141.890 1416.110 2143.070 ;
        RECT 1416.530 2141.890 1417.710 2143.070 ;
        RECT 1414.930 2140.290 1416.110 2141.470 ;
        RECT 1416.530 2140.290 1417.710 2141.470 ;
        RECT 1414.930 1961.890 1416.110 1963.070 ;
        RECT 1416.530 1961.890 1417.710 1963.070 ;
        RECT 1414.930 1960.290 1416.110 1961.470 ;
        RECT 1416.530 1960.290 1417.710 1961.470 ;
        RECT 1414.930 1781.890 1416.110 1783.070 ;
        RECT 1416.530 1781.890 1417.710 1783.070 ;
        RECT 1414.930 1780.290 1416.110 1781.470 ;
        RECT 1416.530 1780.290 1417.710 1781.470 ;
        RECT 1414.930 1601.890 1416.110 1603.070 ;
        RECT 1416.530 1601.890 1417.710 1603.070 ;
        RECT 1414.930 1600.290 1416.110 1601.470 ;
        RECT 1416.530 1600.290 1417.710 1601.470 ;
        RECT 1414.930 1421.890 1416.110 1423.070 ;
        RECT 1416.530 1421.890 1417.710 1423.070 ;
        RECT 1414.930 1420.290 1416.110 1421.470 ;
        RECT 1416.530 1420.290 1417.710 1421.470 ;
        RECT 1414.930 1241.890 1416.110 1243.070 ;
        RECT 1416.530 1241.890 1417.710 1243.070 ;
        RECT 1414.930 1240.290 1416.110 1241.470 ;
        RECT 1416.530 1240.290 1417.710 1241.470 ;
        RECT 1414.930 1061.890 1416.110 1063.070 ;
        RECT 1416.530 1061.890 1417.710 1063.070 ;
        RECT 1414.930 1060.290 1416.110 1061.470 ;
        RECT 1416.530 1060.290 1417.710 1061.470 ;
        RECT 1414.930 881.890 1416.110 883.070 ;
        RECT 1416.530 881.890 1417.710 883.070 ;
        RECT 1414.930 880.290 1416.110 881.470 ;
        RECT 1416.530 880.290 1417.710 881.470 ;
        RECT 1414.930 701.890 1416.110 703.070 ;
        RECT 1416.530 701.890 1417.710 703.070 ;
        RECT 1414.930 700.290 1416.110 701.470 ;
        RECT 1416.530 700.290 1417.710 701.470 ;
        RECT 1414.930 521.890 1416.110 523.070 ;
        RECT 1416.530 521.890 1417.710 523.070 ;
        RECT 1414.930 520.290 1416.110 521.470 ;
        RECT 1416.530 520.290 1417.710 521.470 ;
        RECT 1414.930 341.890 1416.110 343.070 ;
        RECT 1416.530 341.890 1417.710 343.070 ;
        RECT 1414.930 340.290 1416.110 341.470 ;
        RECT 1416.530 340.290 1417.710 341.470 ;
        RECT 1414.930 161.890 1416.110 163.070 ;
        RECT 1416.530 161.890 1417.710 163.070 ;
        RECT 1414.930 160.290 1416.110 161.470 ;
        RECT 1416.530 160.290 1417.710 161.470 ;
        RECT 1414.930 -36.510 1416.110 -35.330 ;
        RECT 1416.530 -36.510 1417.710 -35.330 ;
        RECT 1414.930 -38.110 1416.110 -36.930 ;
        RECT 1416.530 -38.110 1417.710 -36.930 ;
        RECT 1594.930 3556.610 1596.110 3557.790 ;
        RECT 1596.530 3556.610 1597.710 3557.790 ;
        RECT 1594.930 3555.010 1596.110 3556.190 ;
        RECT 1596.530 3555.010 1597.710 3556.190 ;
        RECT 1594.930 3401.890 1596.110 3403.070 ;
        RECT 1596.530 3401.890 1597.710 3403.070 ;
        RECT 1594.930 3400.290 1596.110 3401.470 ;
        RECT 1596.530 3400.290 1597.710 3401.470 ;
        RECT 1594.930 3221.890 1596.110 3223.070 ;
        RECT 1596.530 3221.890 1597.710 3223.070 ;
        RECT 1594.930 3220.290 1596.110 3221.470 ;
        RECT 1596.530 3220.290 1597.710 3221.470 ;
        RECT 1594.930 3041.890 1596.110 3043.070 ;
        RECT 1596.530 3041.890 1597.710 3043.070 ;
        RECT 1594.930 3040.290 1596.110 3041.470 ;
        RECT 1596.530 3040.290 1597.710 3041.470 ;
        RECT 1594.930 2861.890 1596.110 2863.070 ;
        RECT 1596.530 2861.890 1597.710 2863.070 ;
        RECT 1594.930 2860.290 1596.110 2861.470 ;
        RECT 1596.530 2860.290 1597.710 2861.470 ;
        RECT 1594.930 2681.890 1596.110 2683.070 ;
        RECT 1596.530 2681.890 1597.710 2683.070 ;
        RECT 1594.930 2680.290 1596.110 2681.470 ;
        RECT 1596.530 2680.290 1597.710 2681.470 ;
        RECT 1594.930 2501.890 1596.110 2503.070 ;
        RECT 1596.530 2501.890 1597.710 2503.070 ;
        RECT 1594.930 2500.290 1596.110 2501.470 ;
        RECT 1596.530 2500.290 1597.710 2501.470 ;
        RECT 1594.930 2321.890 1596.110 2323.070 ;
        RECT 1596.530 2321.890 1597.710 2323.070 ;
        RECT 1594.930 2320.290 1596.110 2321.470 ;
        RECT 1596.530 2320.290 1597.710 2321.470 ;
        RECT 1594.930 2141.890 1596.110 2143.070 ;
        RECT 1596.530 2141.890 1597.710 2143.070 ;
        RECT 1594.930 2140.290 1596.110 2141.470 ;
        RECT 1596.530 2140.290 1597.710 2141.470 ;
        RECT 1594.930 1961.890 1596.110 1963.070 ;
        RECT 1596.530 1961.890 1597.710 1963.070 ;
        RECT 1594.930 1960.290 1596.110 1961.470 ;
        RECT 1596.530 1960.290 1597.710 1961.470 ;
        RECT 1594.930 1781.890 1596.110 1783.070 ;
        RECT 1596.530 1781.890 1597.710 1783.070 ;
        RECT 1594.930 1780.290 1596.110 1781.470 ;
        RECT 1596.530 1780.290 1597.710 1781.470 ;
        RECT 1594.930 1601.890 1596.110 1603.070 ;
        RECT 1596.530 1601.890 1597.710 1603.070 ;
        RECT 1594.930 1600.290 1596.110 1601.470 ;
        RECT 1596.530 1600.290 1597.710 1601.470 ;
        RECT 1594.930 1421.890 1596.110 1423.070 ;
        RECT 1596.530 1421.890 1597.710 1423.070 ;
        RECT 1594.930 1420.290 1596.110 1421.470 ;
        RECT 1596.530 1420.290 1597.710 1421.470 ;
        RECT 1594.930 1241.890 1596.110 1243.070 ;
        RECT 1596.530 1241.890 1597.710 1243.070 ;
        RECT 1594.930 1240.290 1596.110 1241.470 ;
        RECT 1596.530 1240.290 1597.710 1241.470 ;
        RECT 1594.930 1061.890 1596.110 1063.070 ;
        RECT 1596.530 1061.890 1597.710 1063.070 ;
        RECT 1594.930 1060.290 1596.110 1061.470 ;
        RECT 1596.530 1060.290 1597.710 1061.470 ;
        RECT 1594.930 881.890 1596.110 883.070 ;
        RECT 1596.530 881.890 1597.710 883.070 ;
        RECT 1594.930 880.290 1596.110 881.470 ;
        RECT 1596.530 880.290 1597.710 881.470 ;
        RECT 1594.930 701.890 1596.110 703.070 ;
        RECT 1596.530 701.890 1597.710 703.070 ;
        RECT 1594.930 700.290 1596.110 701.470 ;
        RECT 1596.530 700.290 1597.710 701.470 ;
        RECT 1594.930 521.890 1596.110 523.070 ;
        RECT 1596.530 521.890 1597.710 523.070 ;
        RECT 1594.930 520.290 1596.110 521.470 ;
        RECT 1596.530 520.290 1597.710 521.470 ;
        RECT 1594.930 341.890 1596.110 343.070 ;
        RECT 1596.530 341.890 1597.710 343.070 ;
        RECT 1594.930 340.290 1596.110 341.470 ;
        RECT 1596.530 340.290 1597.710 341.470 ;
        RECT 1594.930 161.890 1596.110 163.070 ;
        RECT 1596.530 161.890 1597.710 163.070 ;
        RECT 1594.930 160.290 1596.110 161.470 ;
        RECT 1596.530 160.290 1597.710 161.470 ;
        RECT 1594.930 -36.510 1596.110 -35.330 ;
        RECT 1596.530 -36.510 1597.710 -35.330 ;
        RECT 1594.930 -38.110 1596.110 -36.930 ;
        RECT 1596.530 -38.110 1597.710 -36.930 ;
        RECT 1774.930 3556.610 1776.110 3557.790 ;
        RECT 1776.530 3556.610 1777.710 3557.790 ;
        RECT 1774.930 3555.010 1776.110 3556.190 ;
        RECT 1776.530 3555.010 1777.710 3556.190 ;
        RECT 1774.930 3401.890 1776.110 3403.070 ;
        RECT 1776.530 3401.890 1777.710 3403.070 ;
        RECT 1774.930 3400.290 1776.110 3401.470 ;
        RECT 1776.530 3400.290 1777.710 3401.470 ;
        RECT 1774.930 3221.890 1776.110 3223.070 ;
        RECT 1776.530 3221.890 1777.710 3223.070 ;
        RECT 1774.930 3220.290 1776.110 3221.470 ;
        RECT 1776.530 3220.290 1777.710 3221.470 ;
        RECT 1774.930 3041.890 1776.110 3043.070 ;
        RECT 1776.530 3041.890 1777.710 3043.070 ;
        RECT 1774.930 3040.290 1776.110 3041.470 ;
        RECT 1776.530 3040.290 1777.710 3041.470 ;
        RECT 1774.930 2861.890 1776.110 2863.070 ;
        RECT 1776.530 2861.890 1777.710 2863.070 ;
        RECT 1774.930 2860.290 1776.110 2861.470 ;
        RECT 1776.530 2860.290 1777.710 2861.470 ;
        RECT 1774.930 2681.890 1776.110 2683.070 ;
        RECT 1776.530 2681.890 1777.710 2683.070 ;
        RECT 1774.930 2680.290 1776.110 2681.470 ;
        RECT 1776.530 2680.290 1777.710 2681.470 ;
        RECT 1774.930 2501.890 1776.110 2503.070 ;
        RECT 1776.530 2501.890 1777.710 2503.070 ;
        RECT 1774.930 2500.290 1776.110 2501.470 ;
        RECT 1776.530 2500.290 1777.710 2501.470 ;
        RECT 1774.930 2321.890 1776.110 2323.070 ;
        RECT 1776.530 2321.890 1777.710 2323.070 ;
        RECT 1774.930 2320.290 1776.110 2321.470 ;
        RECT 1776.530 2320.290 1777.710 2321.470 ;
        RECT 1774.930 2141.890 1776.110 2143.070 ;
        RECT 1776.530 2141.890 1777.710 2143.070 ;
        RECT 1774.930 2140.290 1776.110 2141.470 ;
        RECT 1776.530 2140.290 1777.710 2141.470 ;
        RECT 1774.930 1961.890 1776.110 1963.070 ;
        RECT 1776.530 1961.890 1777.710 1963.070 ;
        RECT 1774.930 1960.290 1776.110 1961.470 ;
        RECT 1776.530 1960.290 1777.710 1961.470 ;
        RECT 1774.930 1781.890 1776.110 1783.070 ;
        RECT 1776.530 1781.890 1777.710 1783.070 ;
        RECT 1774.930 1780.290 1776.110 1781.470 ;
        RECT 1776.530 1780.290 1777.710 1781.470 ;
        RECT 1774.930 1601.890 1776.110 1603.070 ;
        RECT 1776.530 1601.890 1777.710 1603.070 ;
        RECT 1774.930 1600.290 1776.110 1601.470 ;
        RECT 1776.530 1600.290 1777.710 1601.470 ;
        RECT 1774.930 1421.890 1776.110 1423.070 ;
        RECT 1776.530 1421.890 1777.710 1423.070 ;
        RECT 1774.930 1420.290 1776.110 1421.470 ;
        RECT 1776.530 1420.290 1777.710 1421.470 ;
        RECT 1774.930 1241.890 1776.110 1243.070 ;
        RECT 1776.530 1241.890 1777.710 1243.070 ;
        RECT 1774.930 1240.290 1776.110 1241.470 ;
        RECT 1776.530 1240.290 1777.710 1241.470 ;
        RECT 1774.930 1061.890 1776.110 1063.070 ;
        RECT 1776.530 1061.890 1777.710 1063.070 ;
        RECT 1774.930 1060.290 1776.110 1061.470 ;
        RECT 1776.530 1060.290 1777.710 1061.470 ;
        RECT 1774.930 881.890 1776.110 883.070 ;
        RECT 1776.530 881.890 1777.710 883.070 ;
        RECT 1774.930 880.290 1776.110 881.470 ;
        RECT 1776.530 880.290 1777.710 881.470 ;
        RECT 1774.930 701.890 1776.110 703.070 ;
        RECT 1776.530 701.890 1777.710 703.070 ;
        RECT 1774.930 700.290 1776.110 701.470 ;
        RECT 1776.530 700.290 1777.710 701.470 ;
        RECT 1774.930 521.890 1776.110 523.070 ;
        RECT 1776.530 521.890 1777.710 523.070 ;
        RECT 1774.930 520.290 1776.110 521.470 ;
        RECT 1776.530 520.290 1777.710 521.470 ;
        RECT 1774.930 341.890 1776.110 343.070 ;
        RECT 1776.530 341.890 1777.710 343.070 ;
        RECT 1774.930 340.290 1776.110 341.470 ;
        RECT 1776.530 340.290 1777.710 341.470 ;
        RECT 1774.930 161.890 1776.110 163.070 ;
        RECT 1776.530 161.890 1777.710 163.070 ;
        RECT 1774.930 160.290 1776.110 161.470 ;
        RECT 1776.530 160.290 1777.710 161.470 ;
        RECT 1774.930 -36.510 1776.110 -35.330 ;
        RECT 1776.530 -36.510 1777.710 -35.330 ;
        RECT 1774.930 -38.110 1776.110 -36.930 ;
        RECT 1776.530 -38.110 1777.710 -36.930 ;
        RECT 1954.930 3556.610 1956.110 3557.790 ;
        RECT 1956.530 3556.610 1957.710 3557.790 ;
        RECT 1954.930 3555.010 1956.110 3556.190 ;
        RECT 1956.530 3555.010 1957.710 3556.190 ;
        RECT 1954.930 3401.890 1956.110 3403.070 ;
        RECT 1956.530 3401.890 1957.710 3403.070 ;
        RECT 1954.930 3400.290 1956.110 3401.470 ;
        RECT 1956.530 3400.290 1957.710 3401.470 ;
        RECT 1954.930 3221.890 1956.110 3223.070 ;
        RECT 1956.530 3221.890 1957.710 3223.070 ;
        RECT 1954.930 3220.290 1956.110 3221.470 ;
        RECT 1956.530 3220.290 1957.710 3221.470 ;
        RECT 1954.930 3041.890 1956.110 3043.070 ;
        RECT 1956.530 3041.890 1957.710 3043.070 ;
        RECT 1954.930 3040.290 1956.110 3041.470 ;
        RECT 1956.530 3040.290 1957.710 3041.470 ;
        RECT 1954.930 2861.890 1956.110 2863.070 ;
        RECT 1956.530 2861.890 1957.710 2863.070 ;
        RECT 1954.930 2860.290 1956.110 2861.470 ;
        RECT 1956.530 2860.290 1957.710 2861.470 ;
        RECT 1954.930 2681.890 1956.110 2683.070 ;
        RECT 1956.530 2681.890 1957.710 2683.070 ;
        RECT 1954.930 2680.290 1956.110 2681.470 ;
        RECT 1956.530 2680.290 1957.710 2681.470 ;
        RECT 1954.930 2501.890 1956.110 2503.070 ;
        RECT 1956.530 2501.890 1957.710 2503.070 ;
        RECT 1954.930 2500.290 1956.110 2501.470 ;
        RECT 1956.530 2500.290 1957.710 2501.470 ;
        RECT 1954.930 2321.890 1956.110 2323.070 ;
        RECT 1956.530 2321.890 1957.710 2323.070 ;
        RECT 1954.930 2320.290 1956.110 2321.470 ;
        RECT 1956.530 2320.290 1957.710 2321.470 ;
        RECT 1954.930 2141.890 1956.110 2143.070 ;
        RECT 1956.530 2141.890 1957.710 2143.070 ;
        RECT 1954.930 2140.290 1956.110 2141.470 ;
        RECT 1956.530 2140.290 1957.710 2141.470 ;
        RECT 1954.930 1961.890 1956.110 1963.070 ;
        RECT 1956.530 1961.890 1957.710 1963.070 ;
        RECT 1954.930 1960.290 1956.110 1961.470 ;
        RECT 1956.530 1960.290 1957.710 1961.470 ;
        RECT 1954.930 1781.890 1956.110 1783.070 ;
        RECT 1956.530 1781.890 1957.710 1783.070 ;
        RECT 1954.930 1780.290 1956.110 1781.470 ;
        RECT 1956.530 1780.290 1957.710 1781.470 ;
        RECT 1954.930 1601.890 1956.110 1603.070 ;
        RECT 1956.530 1601.890 1957.710 1603.070 ;
        RECT 1954.930 1600.290 1956.110 1601.470 ;
        RECT 1956.530 1600.290 1957.710 1601.470 ;
        RECT 1954.930 1421.890 1956.110 1423.070 ;
        RECT 1956.530 1421.890 1957.710 1423.070 ;
        RECT 1954.930 1420.290 1956.110 1421.470 ;
        RECT 1956.530 1420.290 1957.710 1421.470 ;
        RECT 1954.930 1241.890 1956.110 1243.070 ;
        RECT 1956.530 1241.890 1957.710 1243.070 ;
        RECT 1954.930 1240.290 1956.110 1241.470 ;
        RECT 1956.530 1240.290 1957.710 1241.470 ;
        RECT 1954.930 1061.890 1956.110 1063.070 ;
        RECT 1956.530 1061.890 1957.710 1063.070 ;
        RECT 1954.930 1060.290 1956.110 1061.470 ;
        RECT 1956.530 1060.290 1957.710 1061.470 ;
        RECT 1954.930 881.890 1956.110 883.070 ;
        RECT 1956.530 881.890 1957.710 883.070 ;
        RECT 1954.930 880.290 1956.110 881.470 ;
        RECT 1956.530 880.290 1957.710 881.470 ;
        RECT 1954.930 701.890 1956.110 703.070 ;
        RECT 1956.530 701.890 1957.710 703.070 ;
        RECT 1954.930 700.290 1956.110 701.470 ;
        RECT 1956.530 700.290 1957.710 701.470 ;
        RECT 1954.930 521.890 1956.110 523.070 ;
        RECT 1956.530 521.890 1957.710 523.070 ;
        RECT 1954.930 520.290 1956.110 521.470 ;
        RECT 1956.530 520.290 1957.710 521.470 ;
        RECT 1954.930 341.890 1956.110 343.070 ;
        RECT 1956.530 341.890 1957.710 343.070 ;
        RECT 1954.930 340.290 1956.110 341.470 ;
        RECT 1956.530 340.290 1957.710 341.470 ;
        RECT 1954.930 161.890 1956.110 163.070 ;
        RECT 1956.530 161.890 1957.710 163.070 ;
        RECT 1954.930 160.290 1956.110 161.470 ;
        RECT 1956.530 160.290 1957.710 161.470 ;
        RECT 1954.930 -36.510 1956.110 -35.330 ;
        RECT 1956.530 -36.510 1957.710 -35.330 ;
        RECT 1954.930 -38.110 1956.110 -36.930 ;
        RECT 1956.530 -38.110 1957.710 -36.930 ;
        RECT 2134.930 3556.610 2136.110 3557.790 ;
        RECT 2136.530 3556.610 2137.710 3557.790 ;
        RECT 2134.930 3555.010 2136.110 3556.190 ;
        RECT 2136.530 3555.010 2137.710 3556.190 ;
        RECT 2134.930 3401.890 2136.110 3403.070 ;
        RECT 2136.530 3401.890 2137.710 3403.070 ;
        RECT 2134.930 3400.290 2136.110 3401.470 ;
        RECT 2136.530 3400.290 2137.710 3401.470 ;
        RECT 2134.930 3221.890 2136.110 3223.070 ;
        RECT 2136.530 3221.890 2137.710 3223.070 ;
        RECT 2134.930 3220.290 2136.110 3221.470 ;
        RECT 2136.530 3220.290 2137.710 3221.470 ;
        RECT 2134.930 3041.890 2136.110 3043.070 ;
        RECT 2136.530 3041.890 2137.710 3043.070 ;
        RECT 2134.930 3040.290 2136.110 3041.470 ;
        RECT 2136.530 3040.290 2137.710 3041.470 ;
        RECT 2134.930 2861.890 2136.110 2863.070 ;
        RECT 2136.530 2861.890 2137.710 2863.070 ;
        RECT 2134.930 2860.290 2136.110 2861.470 ;
        RECT 2136.530 2860.290 2137.710 2861.470 ;
        RECT 2134.930 2681.890 2136.110 2683.070 ;
        RECT 2136.530 2681.890 2137.710 2683.070 ;
        RECT 2134.930 2680.290 2136.110 2681.470 ;
        RECT 2136.530 2680.290 2137.710 2681.470 ;
        RECT 2134.930 2501.890 2136.110 2503.070 ;
        RECT 2136.530 2501.890 2137.710 2503.070 ;
        RECT 2134.930 2500.290 2136.110 2501.470 ;
        RECT 2136.530 2500.290 2137.710 2501.470 ;
        RECT 2134.930 2321.890 2136.110 2323.070 ;
        RECT 2136.530 2321.890 2137.710 2323.070 ;
        RECT 2134.930 2320.290 2136.110 2321.470 ;
        RECT 2136.530 2320.290 2137.710 2321.470 ;
        RECT 2134.930 2141.890 2136.110 2143.070 ;
        RECT 2136.530 2141.890 2137.710 2143.070 ;
        RECT 2134.930 2140.290 2136.110 2141.470 ;
        RECT 2136.530 2140.290 2137.710 2141.470 ;
        RECT 2134.930 1961.890 2136.110 1963.070 ;
        RECT 2136.530 1961.890 2137.710 1963.070 ;
        RECT 2134.930 1960.290 2136.110 1961.470 ;
        RECT 2136.530 1960.290 2137.710 1961.470 ;
        RECT 2134.930 1781.890 2136.110 1783.070 ;
        RECT 2136.530 1781.890 2137.710 1783.070 ;
        RECT 2134.930 1780.290 2136.110 1781.470 ;
        RECT 2136.530 1780.290 2137.710 1781.470 ;
        RECT 2134.930 1601.890 2136.110 1603.070 ;
        RECT 2136.530 1601.890 2137.710 1603.070 ;
        RECT 2134.930 1600.290 2136.110 1601.470 ;
        RECT 2136.530 1600.290 2137.710 1601.470 ;
        RECT 2134.930 1421.890 2136.110 1423.070 ;
        RECT 2136.530 1421.890 2137.710 1423.070 ;
        RECT 2134.930 1420.290 2136.110 1421.470 ;
        RECT 2136.530 1420.290 2137.710 1421.470 ;
        RECT 2134.930 1241.890 2136.110 1243.070 ;
        RECT 2136.530 1241.890 2137.710 1243.070 ;
        RECT 2134.930 1240.290 2136.110 1241.470 ;
        RECT 2136.530 1240.290 2137.710 1241.470 ;
        RECT 2134.930 1061.890 2136.110 1063.070 ;
        RECT 2136.530 1061.890 2137.710 1063.070 ;
        RECT 2134.930 1060.290 2136.110 1061.470 ;
        RECT 2136.530 1060.290 2137.710 1061.470 ;
        RECT 2134.930 881.890 2136.110 883.070 ;
        RECT 2136.530 881.890 2137.710 883.070 ;
        RECT 2134.930 880.290 2136.110 881.470 ;
        RECT 2136.530 880.290 2137.710 881.470 ;
        RECT 2134.930 701.890 2136.110 703.070 ;
        RECT 2136.530 701.890 2137.710 703.070 ;
        RECT 2134.930 700.290 2136.110 701.470 ;
        RECT 2136.530 700.290 2137.710 701.470 ;
        RECT 2134.930 521.890 2136.110 523.070 ;
        RECT 2136.530 521.890 2137.710 523.070 ;
        RECT 2134.930 520.290 2136.110 521.470 ;
        RECT 2136.530 520.290 2137.710 521.470 ;
        RECT 2134.930 341.890 2136.110 343.070 ;
        RECT 2136.530 341.890 2137.710 343.070 ;
        RECT 2134.930 340.290 2136.110 341.470 ;
        RECT 2136.530 340.290 2137.710 341.470 ;
        RECT 2134.930 161.890 2136.110 163.070 ;
        RECT 2136.530 161.890 2137.710 163.070 ;
        RECT 2134.930 160.290 2136.110 161.470 ;
        RECT 2136.530 160.290 2137.710 161.470 ;
        RECT 2134.930 -36.510 2136.110 -35.330 ;
        RECT 2136.530 -36.510 2137.710 -35.330 ;
        RECT 2134.930 -38.110 2136.110 -36.930 ;
        RECT 2136.530 -38.110 2137.710 -36.930 ;
        RECT 2314.930 3556.610 2316.110 3557.790 ;
        RECT 2316.530 3556.610 2317.710 3557.790 ;
        RECT 2314.930 3555.010 2316.110 3556.190 ;
        RECT 2316.530 3555.010 2317.710 3556.190 ;
        RECT 2314.930 3401.890 2316.110 3403.070 ;
        RECT 2316.530 3401.890 2317.710 3403.070 ;
        RECT 2314.930 3400.290 2316.110 3401.470 ;
        RECT 2316.530 3400.290 2317.710 3401.470 ;
        RECT 2314.930 3221.890 2316.110 3223.070 ;
        RECT 2316.530 3221.890 2317.710 3223.070 ;
        RECT 2314.930 3220.290 2316.110 3221.470 ;
        RECT 2316.530 3220.290 2317.710 3221.470 ;
        RECT 2314.930 3041.890 2316.110 3043.070 ;
        RECT 2316.530 3041.890 2317.710 3043.070 ;
        RECT 2314.930 3040.290 2316.110 3041.470 ;
        RECT 2316.530 3040.290 2317.710 3041.470 ;
        RECT 2314.930 2861.890 2316.110 2863.070 ;
        RECT 2316.530 2861.890 2317.710 2863.070 ;
        RECT 2314.930 2860.290 2316.110 2861.470 ;
        RECT 2316.530 2860.290 2317.710 2861.470 ;
        RECT 2314.930 2681.890 2316.110 2683.070 ;
        RECT 2316.530 2681.890 2317.710 2683.070 ;
        RECT 2314.930 2680.290 2316.110 2681.470 ;
        RECT 2316.530 2680.290 2317.710 2681.470 ;
        RECT 2314.930 2501.890 2316.110 2503.070 ;
        RECT 2316.530 2501.890 2317.710 2503.070 ;
        RECT 2314.930 2500.290 2316.110 2501.470 ;
        RECT 2316.530 2500.290 2317.710 2501.470 ;
        RECT 2314.930 2321.890 2316.110 2323.070 ;
        RECT 2316.530 2321.890 2317.710 2323.070 ;
        RECT 2314.930 2320.290 2316.110 2321.470 ;
        RECT 2316.530 2320.290 2317.710 2321.470 ;
        RECT 2314.930 2141.890 2316.110 2143.070 ;
        RECT 2316.530 2141.890 2317.710 2143.070 ;
        RECT 2314.930 2140.290 2316.110 2141.470 ;
        RECT 2316.530 2140.290 2317.710 2141.470 ;
        RECT 2314.930 1961.890 2316.110 1963.070 ;
        RECT 2316.530 1961.890 2317.710 1963.070 ;
        RECT 2314.930 1960.290 2316.110 1961.470 ;
        RECT 2316.530 1960.290 2317.710 1961.470 ;
        RECT 2314.930 1781.890 2316.110 1783.070 ;
        RECT 2316.530 1781.890 2317.710 1783.070 ;
        RECT 2314.930 1780.290 2316.110 1781.470 ;
        RECT 2316.530 1780.290 2317.710 1781.470 ;
        RECT 2314.930 1601.890 2316.110 1603.070 ;
        RECT 2316.530 1601.890 2317.710 1603.070 ;
        RECT 2314.930 1600.290 2316.110 1601.470 ;
        RECT 2316.530 1600.290 2317.710 1601.470 ;
        RECT 2314.930 1421.890 2316.110 1423.070 ;
        RECT 2316.530 1421.890 2317.710 1423.070 ;
        RECT 2314.930 1420.290 2316.110 1421.470 ;
        RECT 2316.530 1420.290 2317.710 1421.470 ;
        RECT 2314.930 1241.890 2316.110 1243.070 ;
        RECT 2316.530 1241.890 2317.710 1243.070 ;
        RECT 2314.930 1240.290 2316.110 1241.470 ;
        RECT 2316.530 1240.290 2317.710 1241.470 ;
        RECT 2314.930 1061.890 2316.110 1063.070 ;
        RECT 2316.530 1061.890 2317.710 1063.070 ;
        RECT 2314.930 1060.290 2316.110 1061.470 ;
        RECT 2316.530 1060.290 2317.710 1061.470 ;
        RECT 2314.930 881.890 2316.110 883.070 ;
        RECT 2316.530 881.890 2317.710 883.070 ;
        RECT 2314.930 880.290 2316.110 881.470 ;
        RECT 2316.530 880.290 2317.710 881.470 ;
        RECT 2314.930 701.890 2316.110 703.070 ;
        RECT 2316.530 701.890 2317.710 703.070 ;
        RECT 2314.930 700.290 2316.110 701.470 ;
        RECT 2316.530 700.290 2317.710 701.470 ;
        RECT 2314.930 521.890 2316.110 523.070 ;
        RECT 2316.530 521.890 2317.710 523.070 ;
        RECT 2314.930 520.290 2316.110 521.470 ;
        RECT 2316.530 520.290 2317.710 521.470 ;
        RECT 2314.930 341.890 2316.110 343.070 ;
        RECT 2316.530 341.890 2317.710 343.070 ;
        RECT 2314.930 340.290 2316.110 341.470 ;
        RECT 2316.530 340.290 2317.710 341.470 ;
        RECT 2314.930 161.890 2316.110 163.070 ;
        RECT 2316.530 161.890 2317.710 163.070 ;
        RECT 2314.930 160.290 2316.110 161.470 ;
        RECT 2316.530 160.290 2317.710 161.470 ;
        RECT 2314.930 -36.510 2316.110 -35.330 ;
        RECT 2316.530 -36.510 2317.710 -35.330 ;
        RECT 2314.930 -38.110 2316.110 -36.930 ;
        RECT 2316.530 -38.110 2317.710 -36.930 ;
        RECT 2494.930 3556.610 2496.110 3557.790 ;
        RECT 2496.530 3556.610 2497.710 3557.790 ;
        RECT 2494.930 3555.010 2496.110 3556.190 ;
        RECT 2496.530 3555.010 2497.710 3556.190 ;
        RECT 2494.930 3401.890 2496.110 3403.070 ;
        RECT 2496.530 3401.890 2497.710 3403.070 ;
        RECT 2494.930 3400.290 2496.110 3401.470 ;
        RECT 2496.530 3400.290 2497.710 3401.470 ;
        RECT 2494.930 3221.890 2496.110 3223.070 ;
        RECT 2496.530 3221.890 2497.710 3223.070 ;
        RECT 2494.930 3220.290 2496.110 3221.470 ;
        RECT 2496.530 3220.290 2497.710 3221.470 ;
        RECT 2494.930 3041.890 2496.110 3043.070 ;
        RECT 2496.530 3041.890 2497.710 3043.070 ;
        RECT 2494.930 3040.290 2496.110 3041.470 ;
        RECT 2496.530 3040.290 2497.710 3041.470 ;
        RECT 2494.930 2861.890 2496.110 2863.070 ;
        RECT 2496.530 2861.890 2497.710 2863.070 ;
        RECT 2494.930 2860.290 2496.110 2861.470 ;
        RECT 2496.530 2860.290 2497.710 2861.470 ;
        RECT 2494.930 2681.890 2496.110 2683.070 ;
        RECT 2496.530 2681.890 2497.710 2683.070 ;
        RECT 2494.930 2680.290 2496.110 2681.470 ;
        RECT 2496.530 2680.290 2497.710 2681.470 ;
        RECT 2494.930 2501.890 2496.110 2503.070 ;
        RECT 2496.530 2501.890 2497.710 2503.070 ;
        RECT 2494.930 2500.290 2496.110 2501.470 ;
        RECT 2496.530 2500.290 2497.710 2501.470 ;
        RECT 2494.930 2321.890 2496.110 2323.070 ;
        RECT 2496.530 2321.890 2497.710 2323.070 ;
        RECT 2494.930 2320.290 2496.110 2321.470 ;
        RECT 2496.530 2320.290 2497.710 2321.470 ;
        RECT 2494.930 2141.890 2496.110 2143.070 ;
        RECT 2496.530 2141.890 2497.710 2143.070 ;
        RECT 2494.930 2140.290 2496.110 2141.470 ;
        RECT 2496.530 2140.290 2497.710 2141.470 ;
        RECT 2494.930 1961.890 2496.110 1963.070 ;
        RECT 2496.530 1961.890 2497.710 1963.070 ;
        RECT 2494.930 1960.290 2496.110 1961.470 ;
        RECT 2496.530 1960.290 2497.710 1961.470 ;
        RECT 2494.930 1781.890 2496.110 1783.070 ;
        RECT 2496.530 1781.890 2497.710 1783.070 ;
        RECT 2494.930 1780.290 2496.110 1781.470 ;
        RECT 2496.530 1780.290 2497.710 1781.470 ;
        RECT 2494.930 1601.890 2496.110 1603.070 ;
        RECT 2496.530 1601.890 2497.710 1603.070 ;
        RECT 2494.930 1600.290 2496.110 1601.470 ;
        RECT 2496.530 1600.290 2497.710 1601.470 ;
        RECT 2494.930 1421.890 2496.110 1423.070 ;
        RECT 2496.530 1421.890 2497.710 1423.070 ;
        RECT 2494.930 1420.290 2496.110 1421.470 ;
        RECT 2496.530 1420.290 2497.710 1421.470 ;
        RECT 2494.930 1241.890 2496.110 1243.070 ;
        RECT 2496.530 1241.890 2497.710 1243.070 ;
        RECT 2494.930 1240.290 2496.110 1241.470 ;
        RECT 2496.530 1240.290 2497.710 1241.470 ;
        RECT 2494.930 1061.890 2496.110 1063.070 ;
        RECT 2496.530 1061.890 2497.710 1063.070 ;
        RECT 2494.930 1060.290 2496.110 1061.470 ;
        RECT 2496.530 1060.290 2497.710 1061.470 ;
        RECT 2494.930 881.890 2496.110 883.070 ;
        RECT 2496.530 881.890 2497.710 883.070 ;
        RECT 2494.930 880.290 2496.110 881.470 ;
        RECT 2496.530 880.290 2497.710 881.470 ;
        RECT 2494.930 701.890 2496.110 703.070 ;
        RECT 2496.530 701.890 2497.710 703.070 ;
        RECT 2494.930 700.290 2496.110 701.470 ;
        RECT 2496.530 700.290 2497.710 701.470 ;
        RECT 2494.930 521.890 2496.110 523.070 ;
        RECT 2496.530 521.890 2497.710 523.070 ;
        RECT 2494.930 520.290 2496.110 521.470 ;
        RECT 2496.530 520.290 2497.710 521.470 ;
        RECT 2494.930 341.890 2496.110 343.070 ;
        RECT 2496.530 341.890 2497.710 343.070 ;
        RECT 2494.930 340.290 2496.110 341.470 ;
        RECT 2496.530 340.290 2497.710 341.470 ;
        RECT 2494.930 161.890 2496.110 163.070 ;
        RECT 2496.530 161.890 2497.710 163.070 ;
        RECT 2494.930 160.290 2496.110 161.470 ;
        RECT 2496.530 160.290 2497.710 161.470 ;
        RECT 2494.930 -36.510 2496.110 -35.330 ;
        RECT 2496.530 -36.510 2497.710 -35.330 ;
        RECT 2494.930 -38.110 2496.110 -36.930 ;
        RECT 2496.530 -38.110 2497.710 -36.930 ;
        RECT 2674.930 3556.610 2676.110 3557.790 ;
        RECT 2676.530 3556.610 2677.710 3557.790 ;
        RECT 2674.930 3555.010 2676.110 3556.190 ;
        RECT 2676.530 3555.010 2677.710 3556.190 ;
        RECT 2674.930 3401.890 2676.110 3403.070 ;
        RECT 2676.530 3401.890 2677.710 3403.070 ;
        RECT 2674.930 3400.290 2676.110 3401.470 ;
        RECT 2676.530 3400.290 2677.710 3401.470 ;
        RECT 2674.930 3221.890 2676.110 3223.070 ;
        RECT 2676.530 3221.890 2677.710 3223.070 ;
        RECT 2674.930 3220.290 2676.110 3221.470 ;
        RECT 2676.530 3220.290 2677.710 3221.470 ;
        RECT 2674.930 3041.890 2676.110 3043.070 ;
        RECT 2676.530 3041.890 2677.710 3043.070 ;
        RECT 2674.930 3040.290 2676.110 3041.470 ;
        RECT 2676.530 3040.290 2677.710 3041.470 ;
        RECT 2674.930 2861.890 2676.110 2863.070 ;
        RECT 2676.530 2861.890 2677.710 2863.070 ;
        RECT 2674.930 2860.290 2676.110 2861.470 ;
        RECT 2676.530 2860.290 2677.710 2861.470 ;
        RECT 2674.930 2681.890 2676.110 2683.070 ;
        RECT 2676.530 2681.890 2677.710 2683.070 ;
        RECT 2674.930 2680.290 2676.110 2681.470 ;
        RECT 2676.530 2680.290 2677.710 2681.470 ;
        RECT 2674.930 2501.890 2676.110 2503.070 ;
        RECT 2676.530 2501.890 2677.710 2503.070 ;
        RECT 2674.930 2500.290 2676.110 2501.470 ;
        RECT 2676.530 2500.290 2677.710 2501.470 ;
        RECT 2674.930 2321.890 2676.110 2323.070 ;
        RECT 2676.530 2321.890 2677.710 2323.070 ;
        RECT 2674.930 2320.290 2676.110 2321.470 ;
        RECT 2676.530 2320.290 2677.710 2321.470 ;
        RECT 2674.930 2141.890 2676.110 2143.070 ;
        RECT 2676.530 2141.890 2677.710 2143.070 ;
        RECT 2674.930 2140.290 2676.110 2141.470 ;
        RECT 2676.530 2140.290 2677.710 2141.470 ;
        RECT 2674.930 1961.890 2676.110 1963.070 ;
        RECT 2676.530 1961.890 2677.710 1963.070 ;
        RECT 2674.930 1960.290 2676.110 1961.470 ;
        RECT 2676.530 1960.290 2677.710 1961.470 ;
        RECT 2674.930 1781.890 2676.110 1783.070 ;
        RECT 2676.530 1781.890 2677.710 1783.070 ;
        RECT 2674.930 1780.290 2676.110 1781.470 ;
        RECT 2676.530 1780.290 2677.710 1781.470 ;
        RECT 2674.930 1601.890 2676.110 1603.070 ;
        RECT 2676.530 1601.890 2677.710 1603.070 ;
        RECT 2674.930 1600.290 2676.110 1601.470 ;
        RECT 2676.530 1600.290 2677.710 1601.470 ;
        RECT 2674.930 1421.890 2676.110 1423.070 ;
        RECT 2676.530 1421.890 2677.710 1423.070 ;
        RECT 2674.930 1420.290 2676.110 1421.470 ;
        RECT 2676.530 1420.290 2677.710 1421.470 ;
        RECT 2674.930 1241.890 2676.110 1243.070 ;
        RECT 2676.530 1241.890 2677.710 1243.070 ;
        RECT 2674.930 1240.290 2676.110 1241.470 ;
        RECT 2676.530 1240.290 2677.710 1241.470 ;
        RECT 2674.930 1061.890 2676.110 1063.070 ;
        RECT 2676.530 1061.890 2677.710 1063.070 ;
        RECT 2674.930 1060.290 2676.110 1061.470 ;
        RECT 2676.530 1060.290 2677.710 1061.470 ;
        RECT 2674.930 881.890 2676.110 883.070 ;
        RECT 2676.530 881.890 2677.710 883.070 ;
        RECT 2674.930 880.290 2676.110 881.470 ;
        RECT 2676.530 880.290 2677.710 881.470 ;
        RECT 2674.930 701.890 2676.110 703.070 ;
        RECT 2676.530 701.890 2677.710 703.070 ;
        RECT 2674.930 700.290 2676.110 701.470 ;
        RECT 2676.530 700.290 2677.710 701.470 ;
        RECT 2674.930 521.890 2676.110 523.070 ;
        RECT 2676.530 521.890 2677.710 523.070 ;
        RECT 2674.930 520.290 2676.110 521.470 ;
        RECT 2676.530 520.290 2677.710 521.470 ;
        RECT 2674.930 341.890 2676.110 343.070 ;
        RECT 2676.530 341.890 2677.710 343.070 ;
        RECT 2674.930 340.290 2676.110 341.470 ;
        RECT 2676.530 340.290 2677.710 341.470 ;
        RECT 2674.930 161.890 2676.110 163.070 ;
        RECT 2676.530 161.890 2677.710 163.070 ;
        RECT 2674.930 160.290 2676.110 161.470 ;
        RECT 2676.530 160.290 2677.710 161.470 ;
        RECT 2674.930 -36.510 2676.110 -35.330 ;
        RECT 2676.530 -36.510 2677.710 -35.330 ;
        RECT 2674.930 -38.110 2676.110 -36.930 ;
        RECT 2676.530 -38.110 2677.710 -36.930 ;
        RECT 2854.930 3556.610 2856.110 3557.790 ;
        RECT 2856.530 3556.610 2857.710 3557.790 ;
        RECT 2854.930 3555.010 2856.110 3556.190 ;
        RECT 2856.530 3555.010 2857.710 3556.190 ;
        RECT 2854.930 3401.890 2856.110 3403.070 ;
        RECT 2856.530 3401.890 2857.710 3403.070 ;
        RECT 2854.930 3400.290 2856.110 3401.470 ;
        RECT 2856.530 3400.290 2857.710 3401.470 ;
        RECT 2854.930 3221.890 2856.110 3223.070 ;
        RECT 2856.530 3221.890 2857.710 3223.070 ;
        RECT 2854.930 3220.290 2856.110 3221.470 ;
        RECT 2856.530 3220.290 2857.710 3221.470 ;
        RECT 2854.930 3041.890 2856.110 3043.070 ;
        RECT 2856.530 3041.890 2857.710 3043.070 ;
        RECT 2854.930 3040.290 2856.110 3041.470 ;
        RECT 2856.530 3040.290 2857.710 3041.470 ;
        RECT 2854.930 2861.890 2856.110 2863.070 ;
        RECT 2856.530 2861.890 2857.710 2863.070 ;
        RECT 2854.930 2860.290 2856.110 2861.470 ;
        RECT 2856.530 2860.290 2857.710 2861.470 ;
        RECT 2854.930 2681.890 2856.110 2683.070 ;
        RECT 2856.530 2681.890 2857.710 2683.070 ;
        RECT 2854.930 2680.290 2856.110 2681.470 ;
        RECT 2856.530 2680.290 2857.710 2681.470 ;
        RECT 2854.930 2501.890 2856.110 2503.070 ;
        RECT 2856.530 2501.890 2857.710 2503.070 ;
        RECT 2854.930 2500.290 2856.110 2501.470 ;
        RECT 2856.530 2500.290 2857.710 2501.470 ;
        RECT 2854.930 2321.890 2856.110 2323.070 ;
        RECT 2856.530 2321.890 2857.710 2323.070 ;
        RECT 2854.930 2320.290 2856.110 2321.470 ;
        RECT 2856.530 2320.290 2857.710 2321.470 ;
        RECT 2854.930 2141.890 2856.110 2143.070 ;
        RECT 2856.530 2141.890 2857.710 2143.070 ;
        RECT 2854.930 2140.290 2856.110 2141.470 ;
        RECT 2856.530 2140.290 2857.710 2141.470 ;
        RECT 2854.930 1961.890 2856.110 1963.070 ;
        RECT 2856.530 1961.890 2857.710 1963.070 ;
        RECT 2854.930 1960.290 2856.110 1961.470 ;
        RECT 2856.530 1960.290 2857.710 1961.470 ;
        RECT 2854.930 1781.890 2856.110 1783.070 ;
        RECT 2856.530 1781.890 2857.710 1783.070 ;
        RECT 2854.930 1780.290 2856.110 1781.470 ;
        RECT 2856.530 1780.290 2857.710 1781.470 ;
        RECT 2854.930 1601.890 2856.110 1603.070 ;
        RECT 2856.530 1601.890 2857.710 1603.070 ;
        RECT 2854.930 1600.290 2856.110 1601.470 ;
        RECT 2856.530 1600.290 2857.710 1601.470 ;
        RECT 2854.930 1421.890 2856.110 1423.070 ;
        RECT 2856.530 1421.890 2857.710 1423.070 ;
        RECT 2854.930 1420.290 2856.110 1421.470 ;
        RECT 2856.530 1420.290 2857.710 1421.470 ;
        RECT 2854.930 1241.890 2856.110 1243.070 ;
        RECT 2856.530 1241.890 2857.710 1243.070 ;
        RECT 2854.930 1240.290 2856.110 1241.470 ;
        RECT 2856.530 1240.290 2857.710 1241.470 ;
        RECT 2854.930 1061.890 2856.110 1063.070 ;
        RECT 2856.530 1061.890 2857.710 1063.070 ;
        RECT 2854.930 1060.290 2856.110 1061.470 ;
        RECT 2856.530 1060.290 2857.710 1061.470 ;
        RECT 2854.930 881.890 2856.110 883.070 ;
        RECT 2856.530 881.890 2857.710 883.070 ;
        RECT 2854.930 880.290 2856.110 881.470 ;
        RECT 2856.530 880.290 2857.710 881.470 ;
        RECT 2854.930 701.890 2856.110 703.070 ;
        RECT 2856.530 701.890 2857.710 703.070 ;
        RECT 2854.930 700.290 2856.110 701.470 ;
        RECT 2856.530 700.290 2857.710 701.470 ;
        RECT 2854.930 521.890 2856.110 523.070 ;
        RECT 2856.530 521.890 2857.710 523.070 ;
        RECT 2854.930 520.290 2856.110 521.470 ;
        RECT 2856.530 520.290 2857.710 521.470 ;
        RECT 2854.930 341.890 2856.110 343.070 ;
        RECT 2856.530 341.890 2857.710 343.070 ;
        RECT 2854.930 340.290 2856.110 341.470 ;
        RECT 2856.530 340.290 2857.710 341.470 ;
        RECT 2854.930 161.890 2856.110 163.070 ;
        RECT 2856.530 161.890 2857.710 163.070 ;
        RECT 2854.930 160.290 2856.110 161.470 ;
        RECT 2856.530 160.290 2857.710 161.470 ;
        RECT 2854.930 -36.510 2856.110 -35.330 ;
        RECT 2856.530 -36.510 2857.710 -35.330 ;
        RECT 2854.930 -38.110 2856.110 -36.930 ;
        RECT 2856.530 -38.110 2857.710 -36.930 ;
        RECT 2960.310 3556.610 2961.490 3557.790 ;
        RECT 2961.910 3556.610 2963.090 3557.790 ;
        RECT 2960.310 3555.010 2961.490 3556.190 ;
        RECT 2961.910 3555.010 2963.090 3556.190 ;
        RECT 2960.310 3401.890 2961.490 3403.070 ;
        RECT 2961.910 3401.890 2963.090 3403.070 ;
        RECT 2960.310 3400.290 2961.490 3401.470 ;
        RECT 2961.910 3400.290 2963.090 3401.470 ;
        RECT 2960.310 3221.890 2961.490 3223.070 ;
        RECT 2961.910 3221.890 2963.090 3223.070 ;
        RECT 2960.310 3220.290 2961.490 3221.470 ;
        RECT 2961.910 3220.290 2963.090 3221.470 ;
        RECT 2960.310 3041.890 2961.490 3043.070 ;
        RECT 2961.910 3041.890 2963.090 3043.070 ;
        RECT 2960.310 3040.290 2961.490 3041.470 ;
        RECT 2961.910 3040.290 2963.090 3041.470 ;
        RECT 2960.310 2861.890 2961.490 2863.070 ;
        RECT 2961.910 2861.890 2963.090 2863.070 ;
        RECT 2960.310 2860.290 2961.490 2861.470 ;
        RECT 2961.910 2860.290 2963.090 2861.470 ;
        RECT 2960.310 2681.890 2961.490 2683.070 ;
        RECT 2961.910 2681.890 2963.090 2683.070 ;
        RECT 2960.310 2680.290 2961.490 2681.470 ;
        RECT 2961.910 2680.290 2963.090 2681.470 ;
        RECT 2960.310 2501.890 2961.490 2503.070 ;
        RECT 2961.910 2501.890 2963.090 2503.070 ;
        RECT 2960.310 2500.290 2961.490 2501.470 ;
        RECT 2961.910 2500.290 2963.090 2501.470 ;
        RECT 2960.310 2321.890 2961.490 2323.070 ;
        RECT 2961.910 2321.890 2963.090 2323.070 ;
        RECT 2960.310 2320.290 2961.490 2321.470 ;
        RECT 2961.910 2320.290 2963.090 2321.470 ;
        RECT 2960.310 2141.890 2961.490 2143.070 ;
        RECT 2961.910 2141.890 2963.090 2143.070 ;
        RECT 2960.310 2140.290 2961.490 2141.470 ;
        RECT 2961.910 2140.290 2963.090 2141.470 ;
        RECT 2960.310 1961.890 2961.490 1963.070 ;
        RECT 2961.910 1961.890 2963.090 1963.070 ;
        RECT 2960.310 1960.290 2961.490 1961.470 ;
        RECT 2961.910 1960.290 2963.090 1961.470 ;
        RECT 2960.310 1781.890 2961.490 1783.070 ;
        RECT 2961.910 1781.890 2963.090 1783.070 ;
        RECT 2960.310 1780.290 2961.490 1781.470 ;
        RECT 2961.910 1780.290 2963.090 1781.470 ;
        RECT 2960.310 1601.890 2961.490 1603.070 ;
        RECT 2961.910 1601.890 2963.090 1603.070 ;
        RECT 2960.310 1600.290 2961.490 1601.470 ;
        RECT 2961.910 1600.290 2963.090 1601.470 ;
        RECT 2960.310 1421.890 2961.490 1423.070 ;
        RECT 2961.910 1421.890 2963.090 1423.070 ;
        RECT 2960.310 1420.290 2961.490 1421.470 ;
        RECT 2961.910 1420.290 2963.090 1421.470 ;
        RECT 2960.310 1241.890 2961.490 1243.070 ;
        RECT 2961.910 1241.890 2963.090 1243.070 ;
        RECT 2960.310 1240.290 2961.490 1241.470 ;
        RECT 2961.910 1240.290 2963.090 1241.470 ;
        RECT 2960.310 1061.890 2961.490 1063.070 ;
        RECT 2961.910 1061.890 2963.090 1063.070 ;
        RECT 2960.310 1060.290 2961.490 1061.470 ;
        RECT 2961.910 1060.290 2963.090 1061.470 ;
        RECT 2960.310 881.890 2961.490 883.070 ;
        RECT 2961.910 881.890 2963.090 883.070 ;
        RECT 2960.310 880.290 2961.490 881.470 ;
        RECT 2961.910 880.290 2963.090 881.470 ;
        RECT 2960.310 701.890 2961.490 703.070 ;
        RECT 2961.910 701.890 2963.090 703.070 ;
        RECT 2960.310 700.290 2961.490 701.470 ;
        RECT 2961.910 700.290 2963.090 701.470 ;
        RECT 2960.310 521.890 2961.490 523.070 ;
        RECT 2961.910 521.890 2963.090 523.070 ;
        RECT 2960.310 520.290 2961.490 521.470 ;
        RECT 2961.910 520.290 2963.090 521.470 ;
        RECT 2960.310 341.890 2961.490 343.070 ;
        RECT 2961.910 341.890 2963.090 343.070 ;
        RECT 2960.310 340.290 2961.490 341.470 ;
        RECT 2961.910 340.290 2963.090 341.470 ;
        RECT 2960.310 161.890 2961.490 163.070 ;
        RECT 2961.910 161.890 2963.090 163.070 ;
        RECT 2960.310 160.290 2961.490 161.470 ;
        RECT 2961.910 160.290 2963.090 161.470 ;
        RECT 2960.310 -36.510 2961.490 -35.330 ;
        RECT 2961.910 -36.510 2963.090 -35.330 ;
        RECT 2960.310 -38.110 2961.490 -36.930 ;
        RECT 2961.910 -38.110 2963.090 -36.930 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
        RECT -43.630 880.130 2963.250 883.230 ;
        RECT -43.630 700.130 2963.250 703.230 ;
        RECT -43.630 520.130 2963.250 523.230 ;
        RECT -43.630 340.130 2963.250 343.230 ;
        RECT -43.630 160.130 2963.250 163.230 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
        RECT 278.970 1010.000 282.070 3529.150 ;
        RECT 458.970 1010.000 462.070 3529.150 ;
        RECT 638.970 1010.000 642.070 3529.150 ;
        RECT 818.970 1010.000 822.070 3529.150 ;
        RECT 998.970 1010.000 1002.070 3529.150 ;
        RECT 297.840 410.640 299.440 987.760 ;
        RECT 451.440 410.640 453.040 987.760 ;
        RECT 605.040 410.640 606.640 987.760 ;
        RECT 758.640 410.640 760.240 987.760 ;
        RECT 912.240 410.640 913.840 987.760 ;
        RECT 1065.840 410.640 1067.440 987.760 ;
        RECT 278.970 -9.470 282.070 390.000 ;
        RECT 458.970 -9.470 462.070 390.000 ;
        RECT 638.970 -9.470 642.070 390.000 ;
        RECT 818.970 -9.470 822.070 390.000 ;
        RECT 998.970 -9.470 1002.070 390.000 ;
        RECT 1178.970 -9.470 1182.070 3529.150 ;
        RECT 1358.970 -9.470 1362.070 3529.150 ;
        RECT 1538.970 -9.470 1542.070 3529.150 ;
        RECT 1718.970 -9.470 1722.070 3529.150 ;
        RECT 1898.970 -9.470 1902.070 3529.150 ;
        RECT 2078.970 -9.470 2082.070 3529.150 ;
        RECT 2258.970 -9.470 2262.070 3529.150 ;
        RECT 2438.970 -9.470 2442.070 3529.150 ;
        RECT 2618.970 -9.470 2622.070 3529.150 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER via4 ;
        RECT -14.670 3527.810 -13.490 3528.990 ;
        RECT -13.070 3527.810 -11.890 3528.990 ;
        RECT -14.670 3526.210 -13.490 3527.390 ;
        RECT -13.070 3526.210 -11.890 3527.390 ;
        RECT -14.670 3346.090 -13.490 3347.270 ;
        RECT -13.070 3346.090 -11.890 3347.270 ;
        RECT -14.670 3344.490 -13.490 3345.670 ;
        RECT -13.070 3344.490 -11.890 3345.670 ;
        RECT -14.670 3166.090 -13.490 3167.270 ;
        RECT -13.070 3166.090 -11.890 3167.270 ;
        RECT -14.670 3164.490 -13.490 3165.670 ;
        RECT -13.070 3164.490 -11.890 3165.670 ;
        RECT -14.670 2986.090 -13.490 2987.270 ;
        RECT -13.070 2986.090 -11.890 2987.270 ;
        RECT -14.670 2984.490 -13.490 2985.670 ;
        RECT -13.070 2984.490 -11.890 2985.670 ;
        RECT -14.670 2806.090 -13.490 2807.270 ;
        RECT -13.070 2806.090 -11.890 2807.270 ;
        RECT -14.670 2804.490 -13.490 2805.670 ;
        RECT -13.070 2804.490 -11.890 2805.670 ;
        RECT -14.670 2626.090 -13.490 2627.270 ;
        RECT -13.070 2626.090 -11.890 2627.270 ;
        RECT -14.670 2624.490 -13.490 2625.670 ;
        RECT -13.070 2624.490 -11.890 2625.670 ;
        RECT -14.670 2446.090 -13.490 2447.270 ;
        RECT -13.070 2446.090 -11.890 2447.270 ;
        RECT -14.670 2444.490 -13.490 2445.670 ;
        RECT -13.070 2444.490 -11.890 2445.670 ;
        RECT -14.670 2266.090 -13.490 2267.270 ;
        RECT -13.070 2266.090 -11.890 2267.270 ;
        RECT -14.670 2264.490 -13.490 2265.670 ;
        RECT -13.070 2264.490 -11.890 2265.670 ;
        RECT -14.670 2086.090 -13.490 2087.270 ;
        RECT -13.070 2086.090 -11.890 2087.270 ;
        RECT -14.670 2084.490 -13.490 2085.670 ;
        RECT -13.070 2084.490 -11.890 2085.670 ;
        RECT -14.670 1906.090 -13.490 1907.270 ;
        RECT -13.070 1906.090 -11.890 1907.270 ;
        RECT -14.670 1904.490 -13.490 1905.670 ;
        RECT -13.070 1904.490 -11.890 1905.670 ;
        RECT -14.670 1726.090 -13.490 1727.270 ;
        RECT -13.070 1726.090 -11.890 1727.270 ;
        RECT -14.670 1724.490 -13.490 1725.670 ;
        RECT -13.070 1724.490 -11.890 1725.670 ;
        RECT -14.670 1546.090 -13.490 1547.270 ;
        RECT -13.070 1546.090 -11.890 1547.270 ;
        RECT -14.670 1544.490 -13.490 1545.670 ;
        RECT -13.070 1544.490 -11.890 1545.670 ;
        RECT -14.670 1366.090 -13.490 1367.270 ;
        RECT -13.070 1366.090 -11.890 1367.270 ;
        RECT -14.670 1364.490 -13.490 1365.670 ;
        RECT -13.070 1364.490 -11.890 1365.670 ;
        RECT -14.670 1186.090 -13.490 1187.270 ;
        RECT -13.070 1186.090 -11.890 1187.270 ;
        RECT -14.670 1184.490 -13.490 1185.670 ;
        RECT -13.070 1184.490 -11.890 1185.670 ;
        RECT -14.670 1006.090 -13.490 1007.270 ;
        RECT -13.070 1006.090 -11.890 1007.270 ;
        RECT -14.670 1004.490 -13.490 1005.670 ;
        RECT -13.070 1004.490 -11.890 1005.670 ;
        RECT -14.670 826.090 -13.490 827.270 ;
        RECT -13.070 826.090 -11.890 827.270 ;
        RECT -14.670 824.490 -13.490 825.670 ;
        RECT -13.070 824.490 -11.890 825.670 ;
        RECT -14.670 646.090 -13.490 647.270 ;
        RECT -13.070 646.090 -11.890 647.270 ;
        RECT -14.670 644.490 -13.490 645.670 ;
        RECT -13.070 644.490 -11.890 645.670 ;
        RECT -14.670 466.090 -13.490 467.270 ;
        RECT -13.070 466.090 -11.890 467.270 ;
        RECT -14.670 464.490 -13.490 465.670 ;
        RECT -13.070 464.490 -11.890 465.670 ;
        RECT -14.670 286.090 -13.490 287.270 ;
        RECT -13.070 286.090 -11.890 287.270 ;
        RECT -14.670 284.490 -13.490 285.670 ;
        RECT -13.070 284.490 -11.890 285.670 ;
        RECT -14.670 106.090 -13.490 107.270 ;
        RECT -13.070 106.090 -11.890 107.270 ;
        RECT -14.670 104.490 -13.490 105.670 ;
        RECT -13.070 104.490 -11.890 105.670 ;
        RECT -14.670 -7.710 -13.490 -6.530 ;
        RECT -13.070 -7.710 -11.890 -6.530 ;
        RECT -14.670 -9.310 -13.490 -8.130 ;
        RECT -13.070 -9.310 -11.890 -8.130 ;
        RECT 99.130 3527.810 100.310 3528.990 ;
        RECT 100.730 3527.810 101.910 3528.990 ;
        RECT 99.130 3526.210 100.310 3527.390 ;
        RECT 100.730 3526.210 101.910 3527.390 ;
        RECT 99.130 3346.090 100.310 3347.270 ;
        RECT 100.730 3346.090 101.910 3347.270 ;
        RECT 99.130 3344.490 100.310 3345.670 ;
        RECT 100.730 3344.490 101.910 3345.670 ;
        RECT 99.130 3166.090 100.310 3167.270 ;
        RECT 100.730 3166.090 101.910 3167.270 ;
        RECT 99.130 3164.490 100.310 3165.670 ;
        RECT 100.730 3164.490 101.910 3165.670 ;
        RECT 99.130 2986.090 100.310 2987.270 ;
        RECT 100.730 2986.090 101.910 2987.270 ;
        RECT 99.130 2984.490 100.310 2985.670 ;
        RECT 100.730 2984.490 101.910 2985.670 ;
        RECT 99.130 2806.090 100.310 2807.270 ;
        RECT 100.730 2806.090 101.910 2807.270 ;
        RECT 99.130 2804.490 100.310 2805.670 ;
        RECT 100.730 2804.490 101.910 2805.670 ;
        RECT 99.130 2626.090 100.310 2627.270 ;
        RECT 100.730 2626.090 101.910 2627.270 ;
        RECT 99.130 2624.490 100.310 2625.670 ;
        RECT 100.730 2624.490 101.910 2625.670 ;
        RECT 99.130 2446.090 100.310 2447.270 ;
        RECT 100.730 2446.090 101.910 2447.270 ;
        RECT 99.130 2444.490 100.310 2445.670 ;
        RECT 100.730 2444.490 101.910 2445.670 ;
        RECT 99.130 2266.090 100.310 2267.270 ;
        RECT 100.730 2266.090 101.910 2267.270 ;
        RECT 99.130 2264.490 100.310 2265.670 ;
        RECT 100.730 2264.490 101.910 2265.670 ;
        RECT 99.130 2086.090 100.310 2087.270 ;
        RECT 100.730 2086.090 101.910 2087.270 ;
        RECT 99.130 2084.490 100.310 2085.670 ;
        RECT 100.730 2084.490 101.910 2085.670 ;
        RECT 99.130 1906.090 100.310 1907.270 ;
        RECT 100.730 1906.090 101.910 1907.270 ;
        RECT 99.130 1904.490 100.310 1905.670 ;
        RECT 100.730 1904.490 101.910 1905.670 ;
        RECT 99.130 1726.090 100.310 1727.270 ;
        RECT 100.730 1726.090 101.910 1727.270 ;
        RECT 99.130 1724.490 100.310 1725.670 ;
        RECT 100.730 1724.490 101.910 1725.670 ;
        RECT 99.130 1546.090 100.310 1547.270 ;
        RECT 100.730 1546.090 101.910 1547.270 ;
        RECT 99.130 1544.490 100.310 1545.670 ;
        RECT 100.730 1544.490 101.910 1545.670 ;
        RECT 99.130 1366.090 100.310 1367.270 ;
        RECT 100.730 1366.090 101.910 1367.270 ;
        RECT 99.130 1364.490 100.310 1365.670 ;
        RECT 100.730 1364.490 101.910 1365.670 ;
        RECT 99.130 1186.090 100.310 1187.270 ;
        RECT 100.730 1186.090 101.910 1187.270 ;
        RECT 99.130 1184.490 100.310 1185.670 ;
        RECT 100.730 1184.490 101.910 1185.670 ;
        RECT 279.130 3527.810 280.310 3528.990 ;
        RECT 280.730 3527.810 281.910 3528.990 ;
        RECT 279.130 3526.210 280.310 3527.390 ;
        RECT 280.730 3526.210 281.910 3527.390 ;
        RECT 279.130 3346.090 280.310 3347.270 ;
        RECT 280.730 3346.090 281.910 3347.270 ;
        RECT 279.130 3344.490 280.310 3345.670 ;
        RECT 280.730 3344.490 281.910 3345.670 ;
        RECT 279.130 3166.090 280.310 3167.270 ;
        RECT 280.730 3166.090 281.910 3167.270 ;
        RECT 279.130 3164.490 280.310 3165.670 ;
        RECT 280.730 3164.490 281.910 3165.670 ;
        RECT 279.130 2986.090 280.310 2987.270 ;
        RECT 280.730 2986.090 281.910 2987.270 ;
        RECT 279.130 2984.490 280.310 2985.670 ;
        RECT 280.730 2984.490 281.910 2985.670 ;
        RECT 279.130 2806.090 280.310 2807.270 ;
        RECT 280.730 2806.090 281.910 2807.270 ;
        RECT 279.130 2804.490 280.310 2805.670 ;
        RECT 280.730 2804.490 281.910 2805.670 ;
        RECT 279.130 2626.090 280.310 2627.270 ;
        RECT 280.730 2626.090 281.910 2627.270 ;
        RECT 279.130 2624.490 280.310 2625.670 ;
        RECT 280.730 2624.490 281.910 2625.670 ;
        RECT 279.130 2446.090 280.310 2447.270 ;
        RECT 280.730 2446.090 281.910 2447.270 ;
        RECT 279.130 2444.490 280.310 2445.670 ;
        RECT 280.730 2444.490 281.910 2445.670 ;
        RECT 279.130 2266.090 280.310 2267.270 ;
        RECT 280.730 2266.090 281.910 2267.270 ;
        RECT 279.130 2264.490 280.310 2265.670 ;
        RECT 280.730 2264.490 281.910 2265.670 ;
        RECT 279.130 2086.090 280.310 2087.270 ;
        RECT 280.730 2086.090 281.910 2087.270 ;
        RECT 279.130 2084.490 280.310 2085.670 ;
        RECT 280.730 2084.490 281.910 2085.670 ;
        RECT 279.130 1906.090 280.310 1907.270 ;
        RECT 280.730 1906.090 281.910 1907.270 ;
        RECT 279.130 1904.490 280.310 1905.670 ;
        RECT 280.730 1904.490 281.910 1905.670 ;
        RECT 279.130 1726.090 280.310 1727.270 ;
        RECT 280.730 1726.090 281.910 1727.270 ;
        RECT 279.130 1724.490 280.310 1725.670 ;
        RECT 280.730 1724.490 281.910 1725.670 ;
        RECT 279.130 1546.090 280.310 1547.270 ;
        RECT 280.730 1546.090 281.910 1547.270 ;
        RECT 279.130 1544.490 280.310 1545.670 ;
        RECT 280.730 1544.490 281.910 1545.670 ;
        RECT 279.130 1366.090 280.310 1367.270 ;
        RECT 280.730 1366.090 281.910 1367.270 ;
        RECT 279.130 1364.490 280.310 1365.670 ;
        RECT 280.730 1364.490 281.910 1365.670 ;
        RECT 279.130 1186.090 280.310 1187.270 ;
        RECT 280.730 1186.090 281.910 1187.270 ;
        RECT 279.130 1184.490 280.310 1185.670 ;
        RECT 280.730 1184.490 281.910 1185.670 ;
        RECT 459.130 3527.810 460.310 3528.990 ;
        RECT 460.730 3527.810 461.910 3528.990 ;
        RECT 459.130 3526.210 460.310 3527.390 ;
        RECT 460.730 3526.210 461.910 3527.390 ;
        RECT 459.130 3346.090 460.310 3347.270 ;
        RECT 460.730 3346.090 461.910 3347.270 ;
        RECT 459.130 3344.490 460.310 3345.670 ;
        RECT 460.730 3344.490 461.910 3345.670 ;
        RECT 459.130 3166.090 460.310 3167.270 ;
        RECT 460.730 3166.090 461.910 3167.270 ;
        RECT 459.130 3164.490 460.310 3165.670 ;
        RECT 460.730 3164.490 461.910 3165.670 ;
        RECT 459.130 2986.090 460.310 2987.270 ;
        RECT 460.730 2986.090 461.910 2987.270 ;
        RECT 459.130 2984.490 460.310 2985.670 ;
        RECT 460.730 2984.490 461.910 2985.670 ;
        RECT 459.130 2806.090 460.310 2807.270 ;
        RECT 460.730 2806.090 461.910 2807.270 ;
        RECT 459.130 2804.490 460.310 2805.670 ;
        RECT 460.730 2804.490 461.910 2805.670 ;
        RECT 459.130 2626.090 460.310 2627.270 ;
        RECT 460.730 2626.090 461.910 2627.270 ;
        RECT 459.130 2624.490 460.310 2625.670 ;
        RECT 460.730 2624.490 461.910 2625.670 ;
        RECT 459.130 2446.090 460.310 2447.270 ;
        RECT 460.730 2446.090 461.910 2447.270 ;
        RECT 459.130 2444.490 460.310 2445.670 ;
        RECT 460.730 2444.490 461.910 2445.670 ;
        RECT 459.130 2266.090 460.310 2267.270 ;
        RECT 460.730 2266.090 461.910 2267.270 ;
        RECT 459.130 2264.490 460.310 2265.670 ;
        RECT 460.730 2264.490 461.910 2265.670 ;
        RECT 459.130 2086.090 460.310 2087.270 ;
        RECT 460.730 2086.090 461.910 2087.270 ;
        RECT 459.130 2084.490 460.310 2085.670 ;
        RECT 460.730 2084.490 461.910 2085.670 ;
        RECT 459.130 1906.090 460.310 1907.270 ;
        RECT 460.730 1906.090 461.910 1907.270 ;
        RECT 459.130 1904.490 460.310 1905.670 ;
        RECT 460.730 1904.490 461.910 1905.670 ;
        RECT 459.130 1726.090 460.310 1727.270 ;
        RECT 460.730 1726.090 461.910 1727.270 ;
        RECT 459.130 1724.490 460.310 1725.670 ;
        RECT 460.730 1724.490 461.910 1725.670 ;
        RECT 459.130 1546.090 460.310 1547.270 ;
        RECT 460.730 1546.090 461.910 1547.270 ;
        RECT 459.130 1544.490 460.310 1545.670 ;
        RECT 460.730 1544.490 461.910 1545.670 ;
        RECT 459.130 1366.090 460.310 1367.270 ;
        RECT 460.730 1366.090 461.910 1367.270 ;
        RECT 459.130 1364.490 460.310 1365.670 ;
        RECT 460.730 1364.490 461.910 1365.670 ;
        RECT 459.130 1186.090 460.310 1187.270 ;
        RECT 460.730 1186.090 461.910 1187.270 ;
        RECT 459.130 1184.490 460.310 1185.670 ;
        RECT 460.730 1184.490 461.910 1185.670 ;
        RECT 639.130 3527.810 640.310 3528.990 ;
        RECT 640.730 3527.810 641.910 3528.990 ;
        RECT 639.130 3526.210 640.310 3527.390 ;
        RECT 640.730 3526.210 641.910 3527.390 ;
        RECT 639.130 3346.090 640.310 3347.270 ;
        RECT 640.730 3346.090 641.910 3347.270 ;
        RECT 639.130 3344.490 640.310 3345.670 ;
        RECT 640.730 3344.490 641.910 3345.670 ;
        RECT 639.130 3166.090 640.310 3167.270 ;
        RECT 640.730 3166.090 641.910 3167.270 ;
        RECT 639.130 3164.490 640.310 3165.670 ;
        RECT 640.730 3164.490 641.910 3165.670 ;
        RECT 639.130 2986.090 640.310 2987.270 ;
        RECT 640.730 2986.090 641.910 2987.270 ;
        RECT 639.130 2984.490 640.310 2985.670 ;
        RECT 640.730 2984.490 641.910 2985.670 ;
        RECT 639.130 2806.090 640.310 2807.270 ;
        RECT 640.730 2806.090 641.910 2807.270 ;
        RECT 639.130 2804.490 640.310 2805.670 ;
        RECT 640.730 2804.490 641.910 2805.670 ;
        RECT 639.130 2626.090 640.310 2627.270 ;
        RECT 640.730 2626.090 641.910 2627.270 ;
        RECT 639.130 2624.490 640.310 2625.670 ;
        RECT 640.730 2624.490 641.910 2625.670 ;
        RECT 639.130 2446.090 640.310 2447.270 ;
        RECT 640.730 2446.090 641.910 2447.270 ;
        RECT 639.130 2444.490 640.310 2445.670 ;
        RECT 640.730 2444.490 641.910 2445.670 ;
        RECT 639.130 2266.090 640.310 2267.270 ;
        RECT 640.730 2266.090 641.910 2267.270 ;
        RECT 639.130 2264.490 640.310 2265.670 ;
        RECT 640.730 2264.490 641.910 2265.670 ;
        RECT 639.130 2086.090 640.310 2087.270 ;
        RECT 640.730 2086.090 641.910 2087.270 ;
        RECT 639.130 2084.490 640.310 2085.670 ;
        RECT 640.730 2084.490 641.910 2085.670 ;
        RECT 639.130 1906.090 640.310 1907.270 ;
        RECT 640.730 1906.090 641.910 1907.270 ;
        RECT 639.130 1904.490 640.310 1905.670 ;
        RECT 640.730 1904.490 641.910 1905.670 ;
        RECT 639.130 1726.090 640.310 1727.270 ;
        RECT 640.730 1726.090 641.910 1727.270 ;
        RECT 639.130 1724.490 640.310 1725.670 ;
        RECT 640.730 1724.490 641.910 1725.670 ;
        RECT 639.130 1546.090 640.310 1547.270 ;
        RECT 640.730 1546.090 641.910 1547.270 ;
        RECT 639.130 1544.490 640.310 1545.670 ;
        RECT 640.730 1544.490 641.910 1545.670 ;
        RECT 639.130 1366.090 640.310 1367.270 ;
        RECT 640.730 1366.090 641.910 1367.270 ;
        RECT 639.130 1364.490 640.310 1365.670 ;
        RECT 640.730 1364.490 641.910 1365.670 ;
        RECT 639.130 1186.090 640.310 1187.270 ;
        RECT 640.730 1186.090 641.910 1187.270 ;
        RECT 639.130 1184.490 640.310 1185.670 ;
        RECT 640.730 1184.490 641.910 1185.670 ;
        RECT 819.130 3527.810 820.310 3528.990 ;
        RECT 820.730 3527.810 821.910 3528.990 ;
        RECT 819.130 3526.210 820.310 3527.390 ;
        RECT 820.730 3526.210 821.910 3527.390 ;
        RECT 819.130 3346.090 820.310 3347.270 ;
        RECT 820.730 3346.090 821.910 3347.270 ;
        RECT 819.130 3344.490 820.310 3345.670 ;
        RECT 820.730 3344.490 821.910 3345.670 ;
        RECT 819.130 3166.090 820.310 3167.270 ;
        RECT 820.730 3166.090 821.910 3167.270 ;
        RECT 819.130 3164.490 820.310 3165.670 ;
        RECT 820.730 3164.490 821.910 3165.670 ;
        RECT 819.130 2986.090 820.310 2987.270 ;
        RECT 820.730 2986.090 821.910 2987.270 ;
        RECT 819.130 2984.490 820.310 2985.670 ;
        RECT 820.730 2984.490 821.910 2985.670 ;
        RECT 819.130 2806.090 820.310 2807.270 ;
        RECT 820.730 2806.090 821.910 2807.270 ;
        RECT 819.130 2804.490 820.310 2805.670 ;
        RECT 820.730 2804.490 821.910 2805.670 ;
        RECT 819.130 2626.090 820.310 2627.270 ;
        RECT 820.730 2626.090 821.910 2627.270 ;
        RECT 819.130 2624.490 820.310 2625.670 ;
        RECT 820.730 2624.490 821.910 2625.670 ;
        RECT 819.130 2446.090 820.310 2447.270 ;
        RECT 820.730 2446.090 821.910 2447.270 ;
        RECT 819.130 2444.490 820.310 2445.670 ;
        RECT 820.730 2444.490 821.910 2445.670 ;
        RECT 819.130 2266.090 820.310 2267.270 ;
        RECT 820.730 2266.090 821.910 2267.270 ;
        RECT 819.130 2264.490 820.310 2265.670 ;
        RECT 820.730 2264.490 821.910 2265.670 ;
        RECT 819.130 2086.090 820.310 2087.270 ;
        RECT 820.730 2086.090 821.910 2087.270 ;
        RECT 819.130 2084.490 820.310 2085.670 ;
        RECT 820.730 2084.490 821.910 2085.670 ;
        RECT 819.130 1906.090 820.310 1907.270 ;
        RECT 820.730 1906.090 821.910 1907.270 ;
        RECT 819.130 1904.490 820.310 1905.670 ;
        RECT 820.730 1904.490 821.910 1905.670 ;
        RECT 819.130 1726.090 820.310 1727.270 ;
        RECT 820.730 1726.090 821.910 1727.270 ;
        RECT 819.130 1724.490 820.310 1725.670 ;
        RECT 820.730 1724.490 821.910 1725.670 ;
        RECT 819.130 1546.090 820.310 1547.270 ;
        RECT 820.730 1546.090 821.910 1547.270 ;
        RECT 819.130 1544.490 820.310 1545.670 ;
        RECT 820.730 1544.490 821.910 1545.670 ;
        RECT 819.130 1366.090 820.310 1367.270 ;
        RECT 820.730 1366.090 821.910 1367.270 ;
        RECT 819.130 1364.490 820.310 1365.670 ;
        RECT 820.730 1364.490 821.910 1365.670 ;
        RECT 819.130 1186.090 820.310 1187.270 ;
        RECT 820.730 1186.090 821.910 1187.270 ;
        RECT 819.130 1184.490 820.310 1185.670 ;
        RECT 820.730 1184.490 821.910 1185.670 ;
        RECT 999.130 3527.810 1000.310 3528.990 ;
        RECT 1000.730 3527.810 1001.910 3528.990 ;
        RECT 999.130 3526.210 1000.310 3527.390 ;
        RECT 1000.730 3526.210 1001.910 3527.390 ;
        RECT 999.130 3346.090 1000.310 3347.270 ;
        RECT 1000.730 3346.090 1001.910 3347.270 ;
        RECT 999.130 3344.490 1000.310 3345.670 ;
        RECT 1000.730 3344.490 1001.910 3345.670 ;
        RECT 999.130 3166.090 1000.310 3167.270 ;
        RECT 1000.730 3166.090 1001.910 3167.270 ;
        RECT 999.130 3164.490 1000.310 3165.670 ;
        RECT 1000.730 3164.490 1001.910 3165.670 ;
        RECT 999.130 2986.090 1000.310 2987.270 ;
        RECT 1000.730 2986.090 1001.910 2987.270 ;
        RECT 999.130 2984.490 1000.310 2985.670 ;
        RECT 1000.730 2984.490 1001.910 2985.670 ;
        RECT 999.130 2806.090 1000.310 2807.270 ;
        RECT 1000.730 2806.090 1001.910 2807.270 ;
        RECT 999.130 2804.490 1000.310 2805.670 ;
        RECT 1000.730 2804.490 1001.910 2805.670 ;
        RECT 999.130 2626.090 1000.310 2627.270 ;
        RECT 1000.730 2626.090 1001.910 2627.270 ;
        RECT 999.130 2624.490 1000.310 2625.670 ;
        RECT 1000.730 2624.490 1001.910 2625.670 ;
        RECT 999.130 2446.090 1000.310 2447.270 ;
        RECT 1000.730 2446.090 1001.910 2447.270 ;
        RECT 999.130 2444.490 1000.310 2445.670 ;
        RECT 1000.730 2444.490 1001.910 2445.670 ;
        RECT 999.130 2266.090 1000.310 2267.270 ;
        RECT 1000.730 2266.090 1001.910 2267.270 ;
        RECT 999.130 2264.490 1000.310 2265.670 ;
        RECT 1000.730 2264.490 1001.910 2265.670 ;
        RECT 999.130 2086.090 1000.310 2087.270 ;
        RECT 1000.730 2086.090 1001.910 2087.270 ;
        RECT 999.130 2084.490 1000.310 2085.670 ;
        RECT 1000.730 2084.490 1001.910 2085.670 ;
        RECT 999.130 1906.090 1000.310 1907.270 ;
        RECT 1000.730 1906.090 1001.910 1907.270 ;
        RECT 999.130 1904.490 1000.310 1905.670 ;
        RECT 1000.730 1904.490 1001.910 1905.670 ;
        RECT 999.130 1726.090 1000.310 1727.270 ;
        RECT 1000.730 1726.090 1001.910 1727.270 ;
        RECT 999.130 1724.490 1000.310 1725.670 ;
        RECT 1000.730 1724.490 1001.910 1725.670 ;
        RECT 999.130 1546.090 1000.310 1547.270 ;
        RECT 1000.730 1546.090 1001.910 1547.270 ;
        RECT 999.130 1544.490 1000.310 1545.670 ;
        RECT 1000.730 1544.490 1001.910 1545.670 ;
        RECT 999.130 1366.090 1000.310 1367.270 ;
        RECT 1000.730 1366.090 1001.910 1367.270 ;
        RECT 999.130 1364.490 1000.310 1365.670 ;
        RECT 1000.730 1364.490 1001.910 1365.670 ;
        RECT 999.130 1186.090 1000.310 1187.270 ;
        RECT 1000.730 1186.090 1001.910 1187.270 ;
        RECT 999.130 1184.490 1000.310 1185.670 ;
        RECT 1000.730 1184.490 1001.910 1185.670 ;
        RECT 1179.130 3527.810 1180.310 3528.990 ;
        RECT 1180.730 3527.810 1181.910 3528.990 ;
        RECT 1179.130 3526.210 1180.310 3527.390 ;
        RECT 1180.730 3526.210 1181.910 3527.390 ;
        RECT 1179.130 3346.090 1180.310 3347.270 ;
        RECT 1180.730 3346.090 1181.910 3347.270 ;
        RECT 1179.130 3344.490 1180.310 3345.670 ;
        RECT 1180.730 3344.490 1181.910 3345.670 ;
        RECT 1179.130 3166.090 1180.310 3167.270 ;
        RECT 1180.730 3166.090 1181.910 3167.270 ;
        RECT 1179.130 3164.490 1180.310 3165.670 ;
        RECT 1180.730 3164.490 1181.910 3165.670 ;
        RECT 1179.130 2986.090 1180.310 2987.270 ;
        RECT 1180.730 2986.090 1181.910 2987.270 ;
        RECT 1179.130 2984.490 1180.310 2985.670 ;
        RECT 1180.730 2984.490 1181.910 2985.670 ;
        RECT 1179.130 2806.090 1180.310 2807.270 ;
        RECT 1180.730 2806.090 1181.910 2807.270 ;
        RECT 1179.130 2804.490 1180.310 2805.670 ;
        RECT 1180.730 2804.490 1181.910 2805.670 ;
        RECT 1179.130 2626.090 1180.310 2627.270 ;
        RECT 1180.730 2626.090 1181.910 2627.270 ;
        RECT 1179.130 2624.490 1180.310 2625.670 ;
        RECT 1180.730 2624.490 1181.910 2625.670 ;
        RECT 1179.130 2446.090 1180.310 2447.270 ;
        RECT 1180.730 2446.090 1181.910 2447.270 ;
        RECT 1179.130 2444.490 1180.310 2445.670 ;
        RECT 1180.730 2444.490 1181.910 2445.670 ;
        RECT 1179.130 2266.090 1180.310 2267.270 ;
        RECT 1180.730 2266.090 1181.910 2267.270 ;
        RECT 1179.130 2264.490 1180.310 2265.670 ;
        RECT 1180.730 2264.490 1181.910 2265.670 ;
        RECT 1179.130 2086.090 1180.310 2087.270 ;
        RECT 1180.730 2086.090 1181.910 2087.270 ;
        RECT 1179.130 2084.490 1180.310 2085.670 ;
        RECT 1180.730 2084.490 1181.910 2085.670 ;
        RECT 1179.130 1906.090 1180.310 1907.270 ;
        RECT 1180.730 1906.090 1181.910 1907.270 ;
        RECT 1179.130 1904.490 1180.310 1905.670 ;
        RECT 1180.730 1904.490 1181.910 1905.670 ;
        RECT 1179.130 1726.090 1180.310 1727.270 ;
        RECT 1180.730 1726.090 1181.910 1727.270 ;
        RECT 1179.130 1724.490 1180.310 1725.670 ;
        RECT 1180.730 1724.490 1181.910 1725.670 ;
        RECT 1179.130 1546.090 1180.310 1547.270 ;
        RECT 1180.730 1546.090 1181.910 1547.270 ;
        RECT 1179.130 1544.490 1180.310 1545.670 ;
        RECT 1180.730 1544.490 1181.910 1545.670 ;
        RECT 1179.130 1366.090 1180.310 1367.270 ;
        RECT 1180.730 1366.090 1181.910 1367.270 ;
        RECT 1179.130 1364.490 1180.310 1365.670 ;
        RECT 1180.730 1364.490 1181.910 1365.670 ;
        RECT 1179.130 1186.090 1180.310 1187.270 ;
        RECT 1180.730 1186.090 1181.910 1187.270 ;
        RECT 1179.130 1184.490 1180.310 1185.670 ;
        RECT 1180.730 1184.490 1181.910 1185.670 ;
        RECT 99.130 1006.090 100.310 1007.270 ;
        RECT 100.730 1006.090 101.910 1007.270 ;
        RECT 99.130 1004.490 100.310 1005.670 ;
        RECT 100.730 1004.490 101.910 1005.670 ;
        RECT 1179.130 1006.090 1180.310 1007.270 ;
        RECT 1180.730 1006.090 1181.910 1007.270 ;
        RECT 1179.130 1004.490 1180.310 1005.670 ;
        RECT 1180.730 1004.490 1181.910 1005.670 ;
        RECT 99.130 826.090 100.310 827.270 ;
        RECT 100.730 826.090 101.910 827.270 ;
        RECT 99.130 824.490 100.310 825.670 ;
        RECT 100.730 824.490 101.910 825.670 ;
        RECT 99.130 646.090 100.310 647.270 ;
        RECT 100.730 646.090 101.910 647.270 ;
        RECT 99.130 644.490 100.310 645.670 ;
        RECT 100.730 644.490 101.910 645.670 ;
        RECT 99.130 466.090 100.310 467.270 ;
        RECT 100.730 466.090 101.910 467.270 ;
        RECT 99.130 464.490 100.310 465.670 ;
        RECT 100.730 464.490 101.910 465.670 ;
        RECT 298.050 826.090 299.230 827.270 ;
        RECT 298.050 824.490 299.230 825.670 ;
        RECT 298.050 646.090 299.230 647.270 ;
        RECT 298.050 644.490 299.230 645.670 ;
        RECT 298.050 466.090 299.230 467.270 ;
        RECT 298.050 464.490 299.230 465.670 ;
        RECT 451.650 826.090 452.830 827.270 ;
        RECT 451.650 824.490 452.830 825.670 ;
        RECT 451.650 646.090 452.830 647.270 ;
        RECT 451.650 644.490 452.830 645.670 ;
        RECT 451.650 466.090 452.830 467.270 ;
        RECT 451.650 464.490 452.830 465.670 ;
        RECT 605.250 826.090 606.430 827.270 ;
        RECT 605.250 824.490 606.430 825.670 ;
        RECT 605.250 646.090 606.430 647.270 ;
        RECT 605.250 644.490 606.430 645.670 ;
        RECT 605.250 466.090 606.430 467.270 ;
        RECT 605.250 464.490 606.430 465.670 ;
        RECT 758.850 826.090 760.030 827.270 ;
        RECT 758.850 824.490 760.030 825.670 ;
        RECT 758.850 646.090 760.030 647.270 ;
        RECT 758.850 644.490 760.030 645.670 ;
        RECT 758.850 466.090 760.030 467.270 ;
        RECT 758.850 464.490 760.030 465.670 ;
        RECT 912.450 826.090 913.630 827.270 ;
        RECT 912.450 824.490 913.630 825.670 ;
        RECT 912.450 646.090 913.630 647.270 ;
        RECT 912.450 644.490 913.630 645.670 ;
        RECT 912.450 466.090 913.630 467.270 ;
        RECT 912.450 464.490 913.630 465.670 ;
        RECT 1066.050 826.090 1067.230 827.270 ;
        RECT 1066.050 824.490 1067.230 825.670 ;
        RECT 1066.050 646.090 1067.230 647.270 ;
        RECT 1066.050 644.490 1067.230 645.670 ;
        RECT 1066.050 466.090 1067.230 467.270 ;
        RECT 1066.050 464.490 1067.230 465.670 ;
        RECT 1179.130 826.090 1180.310 827.270 ;
        RECT 1180.730 826.090 1181.910 827.270 ;
        RECT 1179.130 824.490 1180.310 825.670 ;
        RECT 1180.730 824.490 1181.910 825.670 ;
        RECT 1179.130 646.090 1180.310 647.270 ;
        RECT 1180.730 646.090 1181.910 647.270 ;
        RECT 1179.130 644.490 1180.310 645.670 ;
        RECT 1180.730 644.490 1181.910 645.670 ;
        RECT 1179.130 466.090 1180.310 467.270 ;
        RECT 1180.730 466.090 1181.910 467.270 ;
        RECT 1179.130 464.490 1180.310 465.670 ;
        RECT 1180.730 464.490 1181.910 465.670 ;
        RECT 99.130 286.090 100.310 287.270 ;
        RECT 100.730 286.090 101.910 287.270 ;
        RECT 99.130 284.490 100.310 285.670 ;
        RECT 100.730 284.490 101.910 285.670 ;
        RECT 99.130 106.090 100.310 107.270 ;
        RECT 100.730 106.090 101.910 107.270 ;
        RECT 99.130 104.490 100.310 105.670 ;
        RECT 100.730 104.490 101.910 105.670 ;
        RECT 99.130 -7.710 100.310 -6.530 ;
        RECT 100.730 -7.710 101.910 -6.530 ;
        RECT 99.130 -9.310 100.310 -8.130 ;
        RECT 100.730 -9.310 101.910 -8.130 ;
        RECT 279.130 286.090 280.310 287.270 ;
        RECT 280.730 286.090 281.910 287.270 ;
        RECT 279.130 284.490 280.310 285.670 ;
        RECT 280.730 284.490 281.910 285.670 ;
        RECT 279.130 106.090 280.310 107.270 ;
        RECT 280.730 106.090 281.910 107.270 ;
        RECT 279.130 104.490 280.310 105.670 ;
        RECT 280.730 104.490 281.910 105.670 ;
        RECT 279.130 -7.710 280.310 -6.530 ;
        RECT 280.730 -7.710 281.910 -6.530 ;
        RECT 279.130 -9.310 280.310 -8.130 ;
        RECT 280.730 -9.310 281.910 -8.130 ;
        RECT 459.130 286.090 460.310 287.270 ;
        RECT 460.730 286.090 461.910 287.270 ;
        RECT 459.130 284.490 460.310 285.670 ;
        RECT 460.730 284.490 461.910 285.670 ;
        RECT 459.130 106.090 460.310 107.270 ;
        RECT 460.730 106.090 461.910 107.270 ;
        RECT 459.130 104.490 460.310 105.670 ;
        RECT 460.730 104.490 461.910 105.670 ;
        RECT 459.130 -7.710 460.310 -6.530 ;
        RECT 460.730 -7.710 461.910 -6.530 ;
        RECT 459.130 -9.310 460.310 -8.130 ;
        RECT 460.730 -9.310 461.910 -8.130 ;
        RECT 639.130 286.090 640.310 287.270 ;
        RECT 640.730 286.090 641.910 287.270 ;
        RECT 639.130 284.490 640.310 285.670 ;
        RECT 640.730 284.490 641.910 285.670 ;
        RECT 639.130 106.090 640.310 107.270 ;
        RECT 640.730 106.090 641.910 107.270 ;
        RECT 639.130 104.490 640.310 105.670 ;
        RECT 640.730 104.490 641.910 105.670 ;
        RECT 639.130 -7.710 640.310 -6.530 ;
        RECT 640.730 -7.710 641.910 -6.530 ;
        RECT 639.130 -9.310 640.310 -8.130 ;
        RECT 640.730 -9.310 641.910 -8.130 ;
        RECT 819.130 286.090 820.310 287.270 ;
        RECT 820.730 286.090 821.910 287.270 ;
        RECT 819.130 284.490 820.310 285.670 ;
        RECT 820.730 284.490 821.910 285.670 ;
        RECT 819.130 106.090 820.310 107.270 ;
        RECT 820.730 106.090 821.910 107.270 ;
        RECT 819.130 104.490 820.310 105.670 ;
        RECT 820.730 104.490 821.910 105.670 ;
        RECT 819.130 -7.710 820.310 -6.530 ;
        RECT 820.730 -7.710 821.910 -6.530 ;
        RECT 819.130 -9.310 820.310 -8.130 ;
        RECT 820.730 -9.310 821.910 -8.130 ;
        RECT 999.130 286.090 1000.310 287.270 ;
        RECT 1000.730 286.090 1001.910 287.270 ;
        RECT 999.130 284.490 1000.310 285.670 ;
        RECT 1000.730 284.490 1001.910 285.670 ;
        RECT 999.130 106.090 1000.310 107.270 ;
        RECT 1000.730 106.090 1001.910 107.270 ;
        RECT 999.130 104.490 1000.310 105.670 ;
        RECT 1000.730 104.490 1001.910 105.670 ;
        RECT 999.130 -7.710 1000.310 -6.530 ;
        RECT 1000.730 -7.710 1001.910 -6.530 ;
        RECT 999.130 -9.310 1000.310 -8.130 ;
        RECT 1000.730 -9.310 1001.910 -8.130 ;
        RECT 1179.130 286.090 1180.310 287.270 ;
        RECT 1180.730 286.090 1181.910 287.270 ;
        RECT 1179.130 284.490 1180.310 285.670 ;
        RECT 1180.730 284.490 1181.910 285.670 ;
        RECT 1179.130 106.090 1180.310 107.270 ;
        RECT 1180.730 106.090 1181.910 107.270 ;
        RECT 1179.130 104.490 1180.310 105.670 ;
        RECT 1180.730 104.490 1181.910 105.670 ;
        RECT 1179.130 -7.710 1180.310 -6.530 ;
        RECT 1180.730 -7.710 1181.910 -6.530 ;
        RECT 1179.130 -9.310 1180.310 -8.130 ;
        RECT 1180.730 -9.310 1181.910 -8.130 ;
        RECT 1359.130 3527.810 1360.310 3528.990 ;
        RECT 1360.730 3527.810 1361.910 3528.990 ;
        RECT 1359.130 3526.210 1360.310 3527.390 ;
        RECT 1360.730 3526.210 1361.910 3527.390 ;
        RECT 1359.130 3346.090 1360.310 3347.270 ;
        RECT 1360.730 3346.090 1361.910 3347.270 ;
        RECT 1359.130 3344.490 1360.310 3345.670 ;
        RECT 1360.730 3344.490 1361.910 3345.670 ;
        RECT 1359.130 3166.090 1360.310 3167.270 ;
        RECT 1360.730 3166.090 1361.910 3167.270 ;
        RECT 1359.130 3164.490 1360.310 3165.670 ;
        RECT 1360.730 3164.490 1361.910 3165.670 ;
        RECT 1359.130 2986.090 1360.310 2987.270 ;
        RECT 1360.730 2986.090 1361.910 2987.270 ;
        RECT 1359.130 2984.490 1360.310 2985.670 ;
        RECT 1360.730 2984.490 1361.910 2985.670 ;
        RECT 1359.130 2806.090 1360.310 2807.270 ;
        RECT 1360.730 2806.090 1361.910 2807.270 ;
        RECT 1359.130 2804.490 1360.310 2805.670 ;
        RECT 1360.730 2804.490 1361.910 2805.670 ;
        RECT 1359.130 2626.090 1360.310 2627.270 ;
        RECT 1360.730 2626.090 1361.910 2627.270 ;
        RECT 1359.130 2624.490 1360.310 2625.670 ;
        RECT 1360.730 2624.490 1361.910 2625.670 ;
        RECT 1359.130 2446.090 1360.310 2447.270 ;
        RECT 1360.730 2446.090 1361.910 2447.270 ;
        RECT 1359.130 2444.490 1360.310 2445.670 ;
        RECT 1360.730 2444.490 1361.910 2445.670 ;
        RECT 1359.130 2266.090 1360.310 2267.270 ;
        RECT 1360.730 2266.090 1361.910 2267.270 ;
        RECT 1359.130 2264.490 1360.310 2265.670 ;
        RECT 1360.730 2264.490 1361.910 2265.670 ;
        RECT 1359.130 2086.090 1360.310 2087.270 ;
        RECT 1360.730 2086.090 1361.910 2087.270 ;
        RECT 1359.130 2084.490 1360.310 2085.670 ;
        RECT 1360.730 2084.490 1361.910 2085.670 ;
        RECT 1359.130 1906.090 1360.310 1907.270 ;
        RECT 1360.730 1906.090 1361.910 1907.270 ;
        RECT 1359.130 1904.490 1360.310 1905.670 ;
        RECT 1360.730 1904.490 1361.910 1905.670 ;
        RECT 1359.130 1726.090 1360.310 1727.270 ;
        RECT 1360.730 1726.090 1361.910 1727.270 ;
        RECT 1359.130 1724.490 1360.310 1725.670 ;
        RECT 1360.730 1724.490 1361.910 1725.670 ;
        RECT 1359.130 1546.090 1360.310 1547.270 ;
        RECT 1360.730 1546.090 1361.910 1547.270 ;
        RECT 1359.130 1544.490 1360.310 1545.670 ;
        RECT 1360.730 1544.490 1361.910 1545.670 ;
        RECT 1359.130 1366.090 1360.310 1367.270 ;
        RECT 1360.730 1366.090 1361.910 1367.270 ;
        RECT 1359.130 1364.490 1360.310 1365.670 ;
        RECT 1360.730 1364.490 1361.910 1365.670 ;
        RECT 1359.130 1186.090 1360.310 1187.270 ;
        RECT 1360.730 1186.090 1361.910 1187.270 ;
        RECT 1359.130 1184.490 1360.310 1185.670 ;
        RECT 1360.730 1184.490 1361.910 1185.670 ;
        RECT 1359.130 1006.090 1360.310 1007.270 ;
        RECT 1360.730 1006.090 1361.910 1007.270 ;
        RECT 1359.130 1004.490 1360.310 1005.670 ;
        RECT 1360.730 1004.490 1361.910 1005.670 ;
        RECT 1359.130 826.090 1360.310 827.270 ;
        RECT 1360.730 826.090 1361.910 827.270 ;
        RECT 1359.130 824.490 1360.310 825.670 ;
        RECT 1360.730 824.490 1361.910 825.670 ;
        RECT 1359.130 646.090 1360.310 647.270 ;
        RECT 1360.730 646.090 1361.910 647.270 ;
        RECT 1359.130 644.490 1360.310 645.670 ;
        RECT 1360.730 644.490 1361.910 645.670 ;
        RECT 1359.130 466.090 1360.310 467.270 ;
        RECT 1360.730 466.090 1361.910 467.270 ;
        RECT 1359.130 464.490 1360.310 465.670 ;
        RECT 1360.730 464.490 1361.910 465.670 ;
        RECT 1359.130 286.090 1360.310 287.270 ;
        RECT 1360.730 286.090 1361.910 287.270 ;
        RECT 1359.130 284.490 1360.310 285.670 ;
        RECT 1360.730 284.490 1361.910 285.670 ;
        RECT 1359.130 106.090 1360.310 107.270 ;
        RECT 1360.730 106.090 1361.910 107.270 ;
        RECT 1359.130 104.490 1360.310 105.670 ;
        RECT 1360.730 104.490 1361.910 105.670 ;
        RECT 1359.130 -7.710 1360.310 -6.530 ;
        RECT 1360.730 -7.710 1361.910 -6.530 ;
        RECT 1359.130 -9.310 1360.310 -8.130 ;
        RECT 1360.730 -9.310 1361.910 -8.130 ;
        RECT 1539.130 3527.810 1540.310 3528.990 ;
        RECT 1540.730 3527.810 1541.910 3528.990 ;
        RECT 1539.130 3526.210 1540.310 3527.390 ;
        RECT 1540.730 3526.210 1541.910 3527.390 ;
        RECT 1539.130 3346.090 1540.310 3347.270 ;
        RECT 1540.730 3346.090 1541.910 3347.270 ;
        RECT 1539.130 3344.490 1540.310 3345.670 ;
        RECT 1540.730 3344.490 1541.910 3345.670 ;
        RECT 1539.130 3166.090 1540.310 3167.270 ;
        RECT 1540.730 3166.090 1541.910 3167.270 ;
        RECT 1539.130 3164.490 1540.310 3165.670 ;
        RECT 1540.730 3164.490 1541.910 3165.670 ;
        RECT 1539.130 2986.090 1540.310 2987.270 ;
        RECT 1540.730 2986.090 1541.910 2987.270 ;
        RECT 1539.130 2984.490 1540.310 2985.670 ;
        RECT 1540.730 2984.490 1541.910 2985.670 ;
        RECT 1539.130 2806.090 1540.310 2807.270 ;
        RECT 1540.730 2806.090 1541.910 2807.270 ;
        RECT 1539.130 2804.490 1540.310 2805.670 ;
        RECT 1540.730 2804.490 1541.910 2805.670 ;
        RECT 1539.130 2626.090 1540.310 2627.270 ;
        RECT 1540.730 2626.090 1541.910 2627.270 ;
        RECT 1539.130 2624.490 1540.310 2625.670 ;
        RECT 1540.730 2624.490 1541.910 2625.670 ;
        RECT 1539.130 2446.090 1540.310 2447.270 ;
        RECT 1540.730 2446.090 1541.910 2447.270 ;
        RECT 1539.130 2444.490 1540.310 2445.670 ;
        RECT 1540.730 2444.490 1541.910 2445.670 ;
        RECT 1539.130 2266.090 1540.310 2267.270 ;
        RECT 1540.730 2266.090 1541.910 2267.270 ;
        RECT 1539.130 2264.490 1540.310 2265.670 ;
        RECT 1540.730 2264.490 1541.910 2265.670 ;
        RECT 1539.130 2086.090 1540.310 2087.270 ;
        RECT 1540.730 2086.090 1541.910 2087.270 ;
        RECT 1539.130 2084.490 1540.310 2085.670 ;
        RECT 1540.730 2084.490 1541.910 2085.670 ;
        RECT 1539.130 1906.090 1540.310 1907.270 ;
        RECT 1540.730 1906.090 1541.910 1907.270 ;
        RECT 1539.130 1904.490 1540.310 1905.670 ;
        RECT 1540.730 1904.490 1541.910 1905.670 ;
        RECT 1539.130 1726.090 1540.310 1727.270 ;
        RECT 1540.730 1726.090 1541.910 1727.270 ;
        RECT 1539.130 1724.490 1540.310 1725.670 ;
        RECT 1540.730 1724.490 1541.910 1725.670 ;
        RECT 1539.130 1546.090 1540.310 1547.270 ;
        RECT 1540.730 1546.090 1541.910 1547.270 ;
        RECT 1539.130 1544.490 1540.310 1545.670 ;
        RECT 1540.730 1544.490 1541.910 1545.670 ;
        RECT 1539.130 1366.090 1540.310 1367.270 ;
        RECT 1540.730 1366.090 1541.910 1367.270 ;
        RECT 1539.130 1364.490 1540.310 1365.670 ;
        RECT 1540.730 1364.490 1541.910 1365.670 ;
        RECT 1539.130 1186.090 1540.310 1187.270 ;
        RECT 1540.730 1186.090 1541.910 1187.270 ;
        RECT 1539.130 1184.490 1540.310 1185.670 ;
        RECT 1540.730 1184.490 1541.910 1185.670 ;
        RECT 1539.130 1006.090 1540.310 1007.270 ;
        RECT 1540.730 1006.090 1541.910 1007.270 ;
        RECT 1539.130 1004.490 1540.310 1005.670 ;
        RECT 1540.730 1004.490 1541.910 1005.670 ;
        RECT 1539.130 826.090 1540.310 827.270 ;
        RECT 1540.730 826.090 1541.910 827.270 ;
        RECT 1539.130 824.490 1540.310 825.670 ;
        RECT 1540.730 824.490 1541.910 825.670 ;
        RECT 1539.130 646.090 1540.310 647.270 ;
        RECT 1540.730 646.090 1541.910 647.270 ;
        RECT 1539.130 644.490 1540.310 645.670 ;
        RECT 1540.730 644.490 1541.910 645.670 ;
        RECT 1539.130 466.090 1540.310 467.270 ;
        RECT 1540.730 466.090 1541.910 467.270 ;
        RECT 1539.130 464.490 1540.310 465.670 ;
        RECT 1540.730 464.490 1541.910 465.670 ;
        RECT 1539.130 286.090 1540.310 287.270 ;
        RECT 1540.730 286.090 1541.910 287.270 ;
        RECT 1539.130 284.490 1540.310 285.670 ;
        RECT 1540.730 284.490 1541.910 285.670 ;
        RECT 1539.130 106.090 1540.310 107.270 ;
        RECT 1540.730 106.090 1541.910 107.270 ;
        RECT 1539.130 104.490 1540.310 105.670 ;
        RECT 1540.730 104.490 1541.910 105.670 ;
        RECT 1539.130 -7.710 1540.310 -6.530 ;
        RECT 1540.730 -7.710 1541.910 -6.530 ;
        RECT 1539.130 -9.310 1540.310 -8.130 ;
        RECT 1540.730 -9.310 1541.910 -8.130 ;
        RECT 1719.130 3527.810 1720.310 3528.990 ;
        RECT 1720.730 3527.810 1721.910 3528.990 ;
        RECT 1719.130 3526.210 1720.310 3527.390 ;
        RECT 1720.730 3526.210 1721.910 3527.390 ;
        RECT 1719.130 3346.090 1720.310 3347.270 ;
        RECT 1720.730 3346.090 1721.910 3347.270 ;
        RECT 1719.130 3344.490 1720.310 3345.670 ;
        RECT 1720.730 3344.490 1721.910 3345.670 ;
        RECT 1719.130 3166.090 1720.310 3167.270 ;
        RECT 1720.730 3166.090 1721.910 3167.270 ;
        RECT 1719.130 3164.490 1720.310 3165.670 ;
        RECT 1720.730 3164.490 1721.910 3165.670 ;
        RECT 1719.130 2986.090 1720.310 2987.270 ;
        RECT 1720.730 2986.090 1721.910 2987.270 ;
        RECT 1719.130 2984.490 1720.310 2985.670 ;
        RECT 1720.730 2984.490 1721.910 2985.670 ;
        RECT 1719.130 2806.090 1720.310 2807.270 ;
        RECT 1720.730 2806.090 1721.910 2807.270 ;
        RECT 1719.130 2804.490 1720.310 2805.670 ;
        RECT 1720.730 2804.490 1721.910 2805.670 ;
        RECT 1719.130 2626.090 1720.310 2627.270 ;
        RECT 1720.730 2626.090 1721.910 2627.270 ;
        RECT 1719.130 2624.490 1720.310 2625.670 ;
        RECT 1720.730 2624.490 1721.910 2625.670 ;
        RECT 1719.130 2446.090 1720.310 2447.270 ;
        RECT 1720.730 2446.090 1721.910 2447.270 ;
        RECT 1719.130 2444.490 1720.310 2445.670 ;
        RECT 1720.730 2444.490 1721.910 2445.670 ;
        RECT 1719.130 2266.090 1720.310 2267.270 ;
        RECT 1720.730 2266.090 1721.910 2267.270 ;
        RECT 1719.130 2264.490 1720.310 2265.670 ;
        RECT 1720.730 2264.490 1721.910 2265.670 ;
        RECT 1719.130 2086.090 1720.310 2087.270 ;
        RECT 1720.730 2086.090 1721.910 2087.270 ;
        RECT 1719.130 2084.490 1720.310 2085.670 ;
        RECT 1720.730 2084.490 1721.910 2085.670 ;
        RECT 1719.130 1906.090 1720.310 1907.270 ;
        RECT 1720.730 1906.090 1721.910 1907.270 ;
        RECT 1719.130 1904.490 1720.310 1905.670 ;
        RECT 1720.730 1904.490 1721.910 1905.670 ;
        RECT 1719.130 1726.090 1720.310 1727.270 ;
        RECT 1720.730 1726.090 1721.910 1727.270 ;
        RECT 1719.130 1724.490 1720.310 1725.670 ;
        RECT 1720.730 1724.490 1721.910 1725.670 ;
        RECT 1719.130 1546.090 1720.310 1547.270 ;
        RECT 1720.730 1546.090 1721.910 1547.270 ;
        RECT 1719.130 1544.490 1720.310 1545.670 ;
        RECT 1720.730 1544.490 1721.910 1545.670 ;
        RECT 1719.130 1366.090 1720.310 1367.270 ;
        RECT 1720.730 1366.090 1721.910 1367.270 ;
        RECT 1719.130 1364.490 1720.310 1365.670 ;
        RECT 1720.730 1364.490 1721.910 1365.670 ;
        RECT 1719.130 1186.090 1720.310 1187.270 ;
        RECT 1720.730 1186.090 1721.910 1187.270 ;
        RECT 1719.130 1184.490 1720.310 1185.670 ;
        RECT 1720.730 1184.490 1721.910 1185.670 ;
        RECT 1719.130 1006.090 1720.310 1007.270 ;
        RECT 1720.730 1006.090 1721.910 1007.270 ;
        RECT 1719.130 1004.490 1720.310 1005.670 ;
        RECT 1720.730 1004.490 1721.910 1005.670 ;
        RECT 1719.130 826.090 1720.310 827.270 ;
        RECT 1720.730 826.090 1721.910 827.270 ;
        RECT 1719.130 824.490 1720.310 825.670 ;
        RECT 1720.730 824.490 1721.910 825.670 ;
        RECT 1719.130 646.090 1720.310 647.270 ;
        RECT 1720.730 646.090 1721.910 647.270 ;
        RECT 1719.130 644.490 1720.310 645.670 ;
        RECT 1720.730 644.490 1721.910 645.670 ;
        RECT 1719.130 466.090 1720.310 467.270 ;
        RECT 1720.730 466.090 1721.910 467.270 ;
        RECT 1719.130 464.490 1720.310 465.670 ;
        RECT 1720.730 464.490 1721.910 465.670 ;
        RECT 1719.130 286.090 1720.310 287.270 ;
        RECT 1720.730 286.090 1721.910 287.270 ;
        RECT 1719.130 284.490 1720.310 285.670 ;
        RECT 1720.730 284.490 1721.910 285.670 ;
        RECT 1719.130 106.090 1720.310 107.270 ;
        RECT 1720.730 106.090 1721.910 107.270 ;
        RECT 1719.130 104.490 1720.310 105.670 ;
        RECT 1720.730 104.490 1721.910 105.670 ;
        RECT 1719.130 -7.710 1720.310 -6.530 ;
        RECT 1720.730 -7.710 1721.910 -6.530 ;
        RECT 1719.130 -9.310 1720.310 -8.130 ;
        RECT 1720.730 -9.310 1721.910 -8.130 ;
        RECT 1899.130 3527.810 1900.310 3528.990 ;
        RECT 1900.730 3527.810 1901.910 3528.990 ;
        RECT 1899.130 3526.210 1900.310 3527.390 ;
        RECT 1900.730 3526.210 1901.910 3527.390 ;
        RECT 1899.130 3346.090 1900.310 3347.270 ;
        RECT 1900.730 3346.090 1901.910 3347.270 ;
        RECT 1899.130 3344.490 1900.310 3345.670 ;
        RECT 1900.730 3344.490 1901.910 3345.670 ;
        RECT 1899.130 3166.090 1900.310 3167.270 ;
        RECT 1900.730 3166.090 1901.910 3167.270 ;
        RECT 1899.130 3164.490 1900.310 3165.670 ;
        RECT 1900.730 3164.490 1901.910 3165.670 ;
        RECT 1899.130 2986.090 1900.310 2987.270 ;
        RECT 1900.730 2986.090 1901.910 2987.270 ;
        RECT 1899.130 2984.490 1900.310 2985.670 ;
        RECT 1900.730 2984.490 1901.910 2985.670 ;
        RECT 1899.130 2806.090 1900.310 2807.270 ;
        RECT 1900.730 2806.090 1901.910 2807.270 ;
        RECT 1899.130 2804.490 1900.310 2805.670 ;
        RECT 1900.730 2804.490 1901.910 2805.670 ;
        RECT 1899.130 2626.090 1900.310 2627.270 ;
        RECT 1900.730 2626.090 1901.910 2627.270 ;
        RECT 1899.130 2624.490 1900.310 2625.670 ;
        RECT 1900.730 2624.490 1901.910 2625.670 ;
        RECT 1899.130 2446.090 1900.310 2447.270 ;
        RECT 1900.730 2446.090 1901.910 2447.270 ;
        RECT 1899.130 2444.490 1900.310 2445.670 ;
        RECT 1900.730 2444.490 1901.910 2445.670 ;
        RECT 1899.130 2266.090 1900.310 2267.270 ;
        RECT 1900.730 2266.090 1901.910 2267.270 ;
        RECT 1899.130 2264.490 1900.310 2265.670 ;
        RECT 1900.730 2264.490 1901.910 2265.670 ;
        RECT 1899.130 2086.090 1900.310 2087.270 ;
        RECT 1900.730 2086.090 1901.910 2087.270 ;
        RECT 1899.130 2084.490 1900.310 2085.670 ;
        RECT 1900.730 2084.490 1901.910 2085.670 ;
        RECT 1899.130 1906.090 1900.310 1907.270 ;
        RECT 1900.730 1906.090 1901.910 1907.270 ;
        RECT 1899.130 1904.490 1900.310 1905.670 ;
        RECT 1900.730 1904.490 1901.910 1905.670 ;
        RECT 1899.130 1726.090 1900.310 1727.270 ;
        RECT 1900.730 1726.090 1901.910 1727.270 ;
        RECT 1899.130 1724.490 1900.310 1725.670 ;
        RECT 1900.730 1724.490 1901.910 1725.670 ;
        RECT 1899.130 1546.090 1900.310 1547.270 ;
        RECT 1900.730 1546.090 1901.910 1547.270 ;
        RECT 1899.130 1544.490 1900.310 1545.670 ;
        RECT 1900.730 1544.490 1901.910 1545.670 ;
        RECT 1899.130 1366.090 1900.310 1367.270 ;
        RECT 1900.730 1366.090 1901.910 1367.270 ;
        RECT 1899.130 1364.490 1900.310 1365.670 ;
        RECT 1900.730 1364.490 1901.910 1365.670 ;
        RECT 1899.130 1186.090 1900.310 1187.270 ;
        RECT 1900.730 1186.090 1901.910 1187.270 ;
        RECT 1899.130 1184.490 1900.310 1185.670 ;
        RECT 1900.730 1184.490 1901.910 1185.670 ;
        RECT 1899.130 1006.090 1900.310 1007.270 ;
        RECT 1900.730 1006.090 1901.910 1007.270 ;
        RECT 1899.130 1004.490 1900.310 1005.670 ;
        RECT 1900.730 1004.490 1901.910 1005.670 ;
        RECT 1899.130 826.090 1900.310 827.270 ;
        RECT 1900.730 826.090 1901.910 827.270 ;
        RECT 1899.130 824.490 1900.310 825.670 ;
        RECT 1900.730 824.490 1901.910 825.670 ;
        RECT 1899.130 646.090 1900.310 647.270 ;
        RECT 1900.730 646.090 1901.910 647.270 ;
        RECT 1899.130 644.490 1900.310 645.670 ;
        RECT 1900.730 644.490 1901.910 645.670 ;
        RECT 1899.130 466.090 1900.310 467.270 ;
        RECT 1900.730 466.090 1901.910 467.270 ;
        RECT 1899.130 464.490 1900.310 465.670 ;
        RECT 1900.730 464.490 1901.910 465.670 ;
        RECT 1899.130 286.090 1900.310 287.270 ;
        RECT 1900.730 286.090 1901.910 287.270 ;
        RECT 1899.130 284.490 1900.310 285.670 ;
        RECT 1900.730 284.490 1901.910 285.670 ;
        RECT 1899.130 106.090 1900.310 107.270 ;
        RECT 1900.730 106.090 1901.910 107.270 ;
        RECT 1899.130 104.490 1900.310 105.670 ;
        RECT 1900.730 104.490 1901.910 105.670 ;
        RECT 1899.130 -7.710 1900.310 -6.530 ;
        RECT 1900.730 -7.710 1901.910 -6.530 ;
        RECT 1899.130 -9.310 1900.310 -8.130 ;
        RECT 1900.730 -9.310 1901.910 -8.130 ;
        RECT 2079.130 3527.810 2080.310 3528.990 ;
        RECT 2080.730 3527.810 2081.910 3528.990 ;
        RECT 2079.130 3526.210 2080.310 3527.390 ;
        RECT 2080.730 3526.210 2081.910 3527.390 ;
        RECT 2079.130 3346.090 2080.310 3347.270 ;
        RECT 2080.730 3346.090 2081.910 3347.270 ;
        RECT 2079.130 3344.490 2080.310 3345.670 ;
        RECT 2080.730 3344.490 2081.910 3345.670 ;
        RECT 2079.130 3166.090 2080.310 3167.270 ;
        RECT 2080.730 3166.090 2081.910 3167.270 ;
        RECT 2079.130 3164.490 2080.310 3165.670 ;
        RECT 2080.730 3164.490 2081.910 3165.670 ;
        RECT 2079.130 2986.090 2080.310 2987.270 ;
        RECT 2080.730 2986.090 2081.910 2987.270 ;
        RECT 2079.130 2984.490 2080.310 2985.670 ;
        RECT 2080.730 2984.490 2081.910 2985.670 ;
        RECT 2079.130 2806.090 2080.310 2807.270 ;
        RECT 2080.730 2806.090 2081.910 2807.270 ;
        RECT 2079.130 2804.490 2080.310 2805.670 ;
        RECT 2080.730 2804.490 2081.910 2805.670 ;
        RECT 2079.130 2626.090 2080.310 2627.270 ;
        RECT 2080.730 2626.090 2081.910 2627.270 ;
        RECT 2079.130 2624.490 2080.310 2625.670 ;
        RECT 2080.730 2624.490 2081.910 2625.670 ;
        RECT 2079.130 2446.090 2080.310 2447.270 ;
        RECT 2080.730 2446.090 2081.910 2447.270 ;
        RECT 2079.130 2444.490 2080.310 2445.670 ;
        RECT 2080.730 2444.490 2081.910 2445.670 ;
        RECT 2079.130 2266.090 2080.310 2267.270 ;
        RECT 2080.730 2266.090 2081.910 2267.270 ;
        RECT 2079.130 2264.490 2080.310 2265.670 ;
        RECT 2080.730 2264.490 2081.910 2265.670 ;
        RECT 2079.130 2086.090 2080.310 2087.270 ;
        RECT 2080.730 2086.090 2081.910 2087.270 ;
        RECT 2079.130 2084.490 2080.310 2085.670 ;
        RECT 2080.730 2084.490 2081.910 2085.670 ;
        RECT 2079.130 1906.090 2080.310 1907.270 ;
        RECT 2080.730 1906.090 2081.910 1907.270 ;
        RECT 2079.130 1904.490 2080.310 1905.670 ;
        RECT 2080.730 1904.490 2081.910 1905.670 ;
        RECT 2079.130 1726.090 2080.310 1727.270 ;
        RECT 2080.730 1726.090 2081.910 1727.270 ;
        RECT 2079.130 1724.490 2080.310 1725.670 ;
        RECT 2080.730 1724.490 2081.910 1725.670 ;
        RECT 2079.130 1546.090 2080.310 1547.270 ;
        RECT 2080.730 1546.090 2081.910 1547.270 ;
        RECT 2079.130 1544.490 2080.310 1545.670 ;
        RECT 2080.730 1544.490 2081.910 1545.670 ;
        RECT 2079.130 1366.090 2080.310 1367.270 ;
        RECT 2080.730 1366.090 2081.910 1367.270 ;
        RECT 2079.130 1364.490 2080.310 1365.670 ;
        RECT 2080.730 1364.490 2081.910 1365.670 ;
        RECT 2079.130 1186.090 2080.310 1187.270 ;
        RECT 2080.730 1186.090 2081.910 1187.270 ;
        RECT 2079.130 1184.490 2080.310 1185.670 ;
        RECT 2080.730 1184.490 2081.910 1185.670 ;
        RECT 2079.130 1006.090 2080.310 1007.270 ;
        RECT 2080.730 1006.090 2081.910 1007.270 ;
        RECT 2079.130 1004.490 2080.310 1005.670 ;
        RECT 2080.730 1004.490 2081.910 1005.670 ;
        RECT 2079.130 826.090 2080.310 827.270 ;
        RECT 2080.730 826.090 2081.910 827.270 ;
        RECT 2079.130 824.490 2080.310 825.670 ;
        RECT 2080.730 824.490 2081.910 825.670 ;
        RECT 2079.130 646.090 2080.310 647.270 ;
        RECT 2080.730 646.090 2081.910 647.270 ;
        RECT 2079.130 644.490 2080.310 645.670 ;
        RECT 2080.730 644.490 2081.910 645.670 ;
        RECT 2079.130 466.090 2080.310 467.270 ;
        RECT 2080.730 466.090 2081.910 467.270 ;
        RECT 2079.130 464.490 2080.310 465.670 ;
        RECT 2080.730 464.490 2081.910 465.670 ;
        RECT 2079.130 286.090 2080.310 287.270 ;
        RECT 2080.730 286.090 2081.910 287.270 ;
        RECT 2079.130 284.490 2080.310 285.670 ;
        RECT 2080.730 284.490 2081.910 285.670 ;
        RECT 2079.130 106.090 2080.310 107.270 ;
        RECT 2080.730 106.090 2081.910 107.270 ;
        RECT 2079.130 104.490 2080.310 105.670 ;
        RECT 2080.730 104.490 2081.910 105.670 ;
        RECT 2079.130 -7.710 2080.310 -6.530 ;
        RECT 2080.730 -7.710 2081.910 -6.530 ;
        RECT 2079.130 -9.310 2080.310 -8.130 ;
        RECT 2080.730 -9.310 2081.910 -8.130 ;
        RECT 2259.130 3527.810 2260.310 3528.990 ;
        RECT 2260.730 3527.810 2261.910 3528.990 ;
        RECT 2259.130 3526.210 2260.310 3527.390 ;
        RECT 2260.730 3526.210 2261.910 3527.390 ;
        RECT 2259.130 3346.090 2260.310 3347.270 ;
        RECT 2260.730 3346.090 2261.910 3347.270 ;
        RECT 2259.130 3344.490 2260.310 3345.670 ;
        RECT 2260.730 3344.490 2261.910 3345.670 ;
        RECT 2259.130 3166.090 2260.310 3167.270 ;
        RECT 2260.730 3166.090 2261.910 3167.270 ;
        RECT 2259.130 3164.490 2260.310 3165.670 ;
        RECT 2260.730 3164.490 2261.910 3165.670 ;
        RECT 2259.130 2986.090 2260.310 2987.270 ;
        RECT 2260.730 2986.090 2261.910 2987.270 ;
        RECT 2259.130 2984.490 2260.310 2985.670 ;
        RECT 2260.730 2984.490 2261.910 2985.670 ;
        RECT 2259.130 2806.090 2260.310 2807.270 ;
        RECT 2260.730 2806.090 2261.910 2807.270 ;
        RECT 2259.130 2804.490 2260.310 2805.670 ;
        RECT 2260.730 2804.490 2261.910 2805.670 ;
        RECT 2259.130 2626.090 2260.310 2627.270 ;
        RECT 2260.730 2626.090 2261.910 2627.270 ;
        RECT 2259.130 2624.490 2260.310 2625.670 ;
        RECT 2260.730 2624.490 2261.910 2625.670 ;
        RECT 2259.130 2446.090 2260.310 2447.270 ;
        RECT 2260.730 2446.090 2261.910 2447.270 ;
        RECT 2259.130 2444.490 2260.310 2445.670 ;
        RECT 2260.730 2444.490 2261.910 2445.670 ;
        RECT 2259.130 2266.090 2260.310 2267.270 ;
        RECT 2260.730 2266.090 2261.910 2267.270 ;
        RECT 2259.130 2264.490 2260.310 2265.670 ;
        RECT 2260.730 2264.490 2261.910 2265.670 ;
        RECT 2259.130 2086.090 2260.310 2087.270 ;
        RECT 2260.730 2086.090 2261.910 2087.270 ;
        RECT 2259.130 2084.490 2260.310 2085.670 ;
        RECT 2260.730 2084.490 2261.910 2085.670 ;
        RECT 2259.130 1906.090 2260.310 1907.270 ;
        RECT 2260.730 1906.090 2261.910 1907.270 ;
        RECT 2259.130 1904.490 2260.310 1905.670 ;
        RECT 2260.730 1904.490 2261.910 1905.670 ;
        RECT 2259.130 1726.090 2260.310 1727.270 ;
        RECT 2260.730 1726.090 2261.910 1727.270 ;
        RECT 2259.130 1724.490 2260.310 1725.670 ;
        RECT 2260.730 1724.490 2261.910 1725.670 ;
        RECT 2259.130 1546.090 2260.310 1547.270 ;
        RECT 2260.730 1546.090 2261.910 1547.270 ;
        RECT 2259.130 1544.490 2260.310 1545.670 ;
        RECT 2260.730 1544.490 2261.910 1545.670 ;
        RECT 2259.130 1366.090 2260.310 1367.270 ;
        RECT 2260.730 1366.090 2261.910 1367.270 ;
        RECT 2259.130 1364.490 2260.310 1365.670 ;
        RECT 2260.730 1364.490 2261.910 1365.670 ;
        RECT 2259.130 1186.090 2260.310 1187.270 ;
        RECT 2260.730 1186.090 2261.910 1187.270 ;
        RECT 2259.130 1184.490 2260.310 1185.670 ;
        RECT 2260.730 1184.490 2261.910 1185.670 ;
        RECT 2259.130 1006.090 2260.310 1007.270 ;
        RECT 2260.730 1006.090 2261.910 1007.270 ;
        RECT 2259.130 1004.490 2260.310 1005.670 ;
        RECT 2260.730 1004.490 2261.910 1005.670 ;
        RECT 2259.130 826.090 2260.310 827.270 ;
        RECT 2260.730 826.090 2261.910 827.270 ;
        RECT 2259.130 824.490 2260.310 825.670 ;
        RECT 2260.730 824.490 2261.910 825.670 ;
        RECT 2259.130 646.090 2260.310 647.270 ;
        RECT 2260.730 646.090 2261.910 647.270 ;
        RECT 2259.130 644.490 2260.310 645.670 ;
        RECT 2260.730 644.490 2261.910 645.670 ;
        RECT 2259.130 466.090 2260.310 467.270 ;
        RECT 2260.730 466.090 2261.910 467.270 ;
        RECT 2259.130 464.490 2260.310 465.670 ;
        RECT 2260.730 464.490 2261.910 465.670 ;
        RECT 2259.130 286.090 2260.310 287.270 ;
        RECT 2260.730 286.090 2261.910 287.270 ;
        RECT 2259.130 284.490 2260.310 285.670 ;
        RECT 2260.730 284.490 2261.910 285.670 ;
        RECT 2259.130 106.090 2260.310 107.270 ;
        RECT 2260.730 106.090 2261.910 107.270 ;
        RECT 2259.130 104.490 2260.310 105.670 ;
        RECT 2260.730 104.490 2261.910 105.670 ;
        RECT 2259.130 -7.710 2260.310 -6.530 ;
        RECT 2260.730 -7.710 2261.910 -6.530 ;
        RECT 2259.130 -9.310 2260.310 -8.130 ;
        RECT 2260.730 -9.310 2261.910 -8.130 ;
        RECT 2439.130 3527.810 2440.310 3528.990 ;
        RECT 2440.730 3527.810 2441.910 3528.990 ;
        RECT 2439.130 3526.210 2440.310 3527.390 ;
        RECT 2440.730 3526.210 2441.910 3527.390 ;
        RECT 2439.130 3346.090 2440.310 3347.270 ;
        RECT 2440.730 3346.090 2441.910 3347.270 ;
        RECT 2439.130 3344.490 2440.310 3345.670 ;
        RECT 2440.730 3344.490 2441.910 3345.670 ;
        RECT 2439.130 3166.090 2440.310 3167.270 ;
        RECT 2440.730 3166.090 2441.910 3167.270 ;
        RECT 2439.130 3164.490 2440.310 3165.670 ;
        RECT 2440.730 3164.490 2441.910 3165.670 ;
        RECT 2439.130 2986.090 2440.310 2987.270 ;
        RECT 2440.730 2986.090 2441.910 2987.270 ;
        RECT 2439.130 2984.490 2440.310 2985.670 ;
        RECT 2440.730 2984.490 2441.910 2985.670 ;
        RECT 2439.130 2806.090 2440.310 2807.270 ;
        RECT 2440.730 2806.090 2441.910 2807.270 ;
        RECT 2439.130 2804.490 2440.310 2805.670 ;
        RECT 2440.730 2804.490 2441.910 2805.670 ;
        RECT 2439.130 2626.090 2440.310 2627.270 ;
        RECT 2440.730 2626.090 2441.910 2627.270 ;
        RECT 2439.130 2624.490 2440.310 2625.670 ;
        RECT 2440.730 2624.490 2441.910 2625.670 ;
        RECT 2439.130 2446.090 2440.310 2447.270 ;
        RECT 2440.730 2446.090 2441.910 2447.270 ;
        RECT 2439.130 2444.490 2440.310 2445.670 ;
        RECT 2440.730 2444.490 2441.910 2445.670 ;
        RECT 2439.130 2266.090 2440.310 2267.270 ;
        RECT 2440.730 2266.090 2441.910 2267.270 ;
        RECT 2439.130 2264.490 2440.310 2265.670 ;
        RECT 2440.730 2264.490 2441.910 2265.670 ;
        RECT 2439.130 2086.090 2440.310 2087.270 ;
        RECT 2440.730 2086.090 2441.910 2087.270 ;
        RECT 2439.130 2084.490 2440.310 2085.670 ;
        RECT 2440.730 2084.490 2441.910 2085.670 ;
        RECT 2439.130 1906.090 2440.310 1907.270 ;
        RECT 2440.730 1906.090 2441.910 1907.270 ;
        RECT 2439.130 1904.490 2440.310 1905.670 ;
        RECT 2440.730 1904.490 2441.910 1905.670 ;
        RECT 2439.130 1726.090 2440.310 1727.270 ;
        RECT 2440.730 1726.090 2441.910 1727.270 ;
        RECT 2439.130 1724.490 2440.310 1725.670 ;
        RECT 2440.730 1724.490 2441.910 1725.670 ;
        RECT 2439.130 1546.090 2440.310 1547.270 ;
        RECT 2440.730 1546.090 2441.910 1547.270 ;
        RECT 2439.130 1544.490 2440.310 1545.670 ;
        RECT 2440.730 1544.490 2441.910 1545.670 ;
        RECT 2439.130 1366.090 2440.310 1367.270 ;
        RECT 2440.730 1366.090 2441.910 1367.270 ;
        RECT 2439.130 1364.490 2440.310 1365.670 ;
        RECT 2440.730 1364.490 2441.910 1365.670 ;
        RECT 2439.130 1186.090 2440.310 1187.270 ;
        RECT 2440.730 1186.090 2441.910 1187.270 ;
        RECT 2439.130 1184.490 2440.310 1185.670 ;
        RECT 2440.730 1184.490 2441.910 1185.670 ;
        RECT 2439.130 1006.090 2440.310 1007.270 ;
        RECT 2440.730 1006.090 2441.910 1007.270 ;
        RECT 2439.130 1004.490 2440.310 1005.670 ;
        RECT 2440.730 1004.490 2441.910 1005.670 ;
        RECT 2439.130 826.090 2440.310 827.270 ;
        RECT 2440.730 826.090 2441.910 827.270 ;
        RECT 2439.130 824.490 2440.310 825.670 ;
        RECT 2440.730 824.490 2441.910 825.670 ;
        RECT 2439.130 646.090 2440.310 647.270 ;
        RECT 2440.730 646.090 2441.910 647.270 ;
        RECT 2439.130 644.490 2440.310 645.670 ;
        RECT 2440.730 644.490 2441.910 645.670 ;
        RECT 2439.130 466.090 2440.310 467.270 ;
        RECT 2440.730 466.090 2441.910 467.270 ;
        RECT 2439.130 464.490 2440.310 465.670 ;
        RECT 2440.730 464.490 2441.910 465.670 ;
        RECT 2439.130 286.090 2440.310 287.270 ;
        RECT 2440.730 286.090 2441.910 287.270 ;
        RECT 2439.130 284.490 2440.310 285.670 ;
        RECT 2440.730 284.490 2441.910 285.670 ;
        RECT 2439.130 106.090 2440.310 107.270 ;
        RECT 2440.730 106.090 2441.910 107.270 ;
        RECT 2439.130 104.490 2440.310 105.670 ;
        RECT 2440.730 104.490 2441.910 105.670 ;
        RECT 2439.130 -7.710 2440.310 -6.530 ;
        RECT 2440.730 -7.710 2441.910 -6.530 ;
        RECT 2439.130 -9.310 2440.310 -8.130 ;
        RECT 2440.730 -9.310 2441.910 -8.130 ;
        RECT 2619.130 3527.810 2620.310 3528.990 ;
        RECT 2620.730 3527.810 2621.910 3528.990 ;
        RECT 2619.130 3526.210 2620.310 3527.390 ;
        RECT 2620.730 3526.210 2621.910 3527.390 ;
        RECT 2619.130 3346.090 2620.310 3347.270 ;
        RECT 2620.730 3346.090 2621.910 3347.270 ;
        RECT 2619.130 3344.490 2620.310 3345.670 ;
        RECT 2620.730 3344.490 2621.910 3345.670 ;
        RECT 2619.130 3166.090 2620.310 3167.270 ;
        RECT 2620.730 3166.090 2621.910 3167.270 ;
        RECT 2619.130 3164.490 2620.310 3165.670 ;
        RECT 2620.730 3164.490 2621.910 3165.670 ;
        RECT 2619.130 2986.090 2620.310 2987.270 ;
        RECT 2620.730 2986.090 2621.910 2987.270 ;
        RECT 2619.130 2984.490 2620.310 2985.670 ;
        RECT 2620.730 2984.490 2621.910 2985.670 ;
        RECT 2619.130 2806.090 2620.310 2807.270 ;
        RECT 2620.730 2806.090 2621.910 2807.270 ;
        RECT 2619.130 2804.490 2620.310 2805.670 ;
        RECT 2620.730 2804.490 2621.910 2805.670 ;
        RECT 2619.130 2626.090 2620.310 2627.270 ;
        RECT 2620.730 2626.090 2621.910 2627.270 ;
        RECT 2619.130 2624.490 2620.310 2625.670 ;
        RECT 2620.730 2624.490 2621.910 2625.670 ;
        RECT 2619.130 2446.090 2620.310 2447.270 ;
        RECT 2620.730 2446.090 2621.910 2447.270 ;
        RECT 2619.130 2444.490 2620.310 2445.670 ;
        RECT 2620.730 2444.490 2621.910 2445.670 ;
        RECT 2619.130 2266.090 2620.310 2267.270 ;
        RECT 2620.730 2266.090 2621.910 2267.270 ;
        RECT 2619.130 2264.490 2620.310 2265.670 ;
        RECT 2620.730 2264.490 2621.910 2265.670 ;
        RECT 2619.130 2086.090 2620.310 2087.270 ;
        RECT 2620.730 2086.090 2621.910 2087.270 ;
        RECT 2619.130 2084.490 2620.310 2085.670 ;
        RECT 2620.730 2084.490 2621.910 2085.670 ;
        RECT 2619.130 1906.090 2620.310 1907.270 ;
        RECT 2620.730 1906.090 2621.910 1907.270 ;
        RECT 2619.130 1904.490 2620.310 1905.670 ;
        RECT 2620.730 1904.490 2621.910 1905.670 ;
        RECT 2619.130 1726.090 2620.310 1727.270 ;
        RECT 2620.730 1726.090 2621.910 1727.270 ;
        RECT 2619.130 1724.490 2620.310 1725.670 ;
        RECT 2620.730 1724.490 2621.910 1725.670 ;
        RECT 2619.130 1546.090 2620.310 1547.270 ;
        RECT 2620.730 1546.090 2621.910 1547.270 ;
        RECT 2619.130 1544.490 2620.310 1545.670 ;
        RECT 2620.730 1544.490 2621.910 1545.670 ;
        RECT 2619.130 1366.090 2620.310 1367.270 ;
        RECT 2620.730 1366.090 2621.910 1367.270 ;
        RECT 2619.130 1364.490 2620.310 1365.670 ;
        RECT 2620.730 1364.490 2621.910 1365.670 ;
        RECT 2619.130 1186.090 2620.310 1187.270 ;
        RECT 2620.730 1186.090 2621.910 1187.270 ;
        RECT 2619.130 1184.490 2620.310 1185.670 ;
        RECT 2620.730 1184.490 2621.910 1185.670 ;
        RECT 2619.130 1006.090 2620.310 1007.270 ;
        RECT 2620.730 1006.090 2621.910 1007.270 ;
        RECT 2619.130 1004.490 2620.310 1005.670 ;
        RECT 2620.730 1004.490 2621.910 1005.670 ;
        RECT 2619.130 826.090 2620.310 827.270 ;
        RECT 2620.730 826.090 2621.910 827.270 ;
        RECT 2619.130 824.490 2620.310 825.670 ;
        RECT 2620.730 824.490 2621.910 825.670 ;
        RECT 2619.130 646.090 2620.310 647.270 ;
        RECT 2620.730 646.090 2621.910 647.270 ;
        RECT 2619.130 644.490 2620.310 645.670 ;
        RECT 2620.730 644.490 2621.910 645.670 ;
        RECT 2619.130 466.090 2620.310 467.270 ;
        RECT 2620.730 466.090 2621.910 467.270 ;
        RECT 2619.130 464.490 2620.310 465.670 ;
        RECT 2620.730 464.490 2621.910 465.670 ;
        RECT 2619.130 286.090 2620.310 287.270 ;
        RECT 2620.730 286.090 2621.910 287.270 ;
        RECT 2619.130 284.490 2620.310 285.670 ;
        RECT 2620.730 284.490 2621.910 285.670 ;
        RECT 2619.130 106.090 2620.310 107.270 ;
        RECT 2620.730 106.090 2621.910 107.270 ;
        RECT 2619.130 104.490 2620.310 105.670 ;
        RECT 2620.730 104.490 2621.910 105.670 ;
        RECT 2619.130 -7.710 2620.310 -6.530 ;
        RECT 2620.730 -7.710 2621.910 -6.530 ;
        RECT 2619.130 -9.310 2620.310 -8.130 ;
        RECT 2620.730 -9.310 2621.910 -8.130 ;
        RECT 2799.130 3527.810 2800.310 3528.990 ;
        RECT 2800.730 3527.810 2801.910 3528.990 ;
        RECT 2799.130 3526.210 2800.310 3527.390 ;
        RECT 2800.730 3526.210 2801.910 3527.390 ;
        RECT 2799.130 3346.090 2800.310 3347.270 ;
        RECT 2800.730 3346.090 2801.910 3347.270 ;
        RECT 2799.130 3344.490 2800.310 3345.670 ;
        RECT 2800.730 3344.490 2801.910 3345.670 ;
        RECT 2799.130 3166.090 2800.310 3167.270 ;
        RECT 2800.730 3166.090 2801.910 3167.270 ;
        RECT 2799.130 3164.490 2800.310 3165.670 ;
        RECT 2800.730 3164.490 2801.910 3165.670 ;
        RECT 2799.130 2986.090 2800.310 2987.270 ;
        RECT 2800.730 2986.090 2801.910 2987.270 ;
        RECT 2799.130 2984.490 2800.310 2985.670 ;
        RECT 2800.730 2984.490 2801.910 2985.670 ;
        RECT 2799.130 2806.090 2800.310 2807.270 ;
        RECT 2800.730 2806.090 2801.910 2807.270 ;
        RECT 2799.130 2804.490 2800.310 2805.670 ;
        RECT 2800.730 2804.490 2801.910 2805.670 ;
        RECT 2799.130 2626.090 2800.310 2627.270 ;
        RECT 2800.730 2626.090 2801.910 2627.270 ;
        RECT 2799.130 2624.490 2800.310 2625.670 ;
        RECT 2800.730 2624.490 2801.910 2625.670 ;
        RECT 2799.130 2446.090 2800.310 2447.270 ;
        RECT 2800.730 2446.090 2801.910 2447.270 ;
        RECT 2799.130 2444.490 2800.310 2445.670 ;
        RECT 2800.730 2444.490 2801.910 2445.670 ;
        RECT 2799.130 2266.090 2800.310 2267.270 ;
        RECT 2800.730 2266.090 2801.910 2267.270 ;
        RECT 2799.130 2264.490 2800.310 2265.670 ;
        RECT 2800.730 2264.490 2801.910 2265.670 ;
        RECT 2799.130 2086.090 2800.310 2087.270 ;
        RECT 2800.730 2086.090 2801.910 2087.270 ;
        RECT 2799.130 2084.490 2800.310 2085.670 ;
        RECT 2800.730 2084.490 2801.910 2085.670 ;
        RECT 2799.130 1906.090 2800.310 1907.270 ;
        RECT 2800.730 1906.090 2801.910 1907.270 ;
        RECT 2799.130 1904.490 2800.310 1905.670 ;
        RECT 2800.730 1904.490 2801.910 1905.670 ;
        RECT 2799.130 1726.090 2800.310 1727.270 ;
        RECT 2800.730 1726.090 2801.910 1727.270 ;
        RECT 2799.130 1724.490 2800.310 1725.670 ;
        RECT 2800.730 1724.490 2801.910 1725.670 ;
        RECT 2799.130 1546.090 2800.310 1547.270 ;
        RECT 2800.730 1546.090 2801.910 1547.270 ;
        RECT 2799.130 1544.490 2800.310 1545.670 ;
        RECT 2800.730 1544.490 2801.910 1545.670 ;
        RECT 2799.130 1366.090 2800.310 1367.270 ;
        RECT 2800.730 1366.090 2801.910 1367.270 ;
        RECT 2799.130 1364.490 2800.310 1365.670 ;
        RECT 2800.730 1364.490 2801.910 1365.670 ;
        RECT 2799.130 1186.090 2800.310 1187.270 ;
        RECT 2800.730 1186.090 2801.910 1187.270 ;
        RECT 2799.130 1184.490 2800.310 1185.670 ;
        RECT 2800.730 1184.490 2801.910 1185.670 ;
        RECT 2799.130 1006.090 2800.310 1007.270 ;
        RECT 2800.730 1006.090 2801.910 1007.270 ;
        RECT 2799.130 1004.490 2800.310 1005.670 ;
        RECT 2800.730 1004.490 2801.910 1005.670 ;
        RECT 2799.130 826.090 2800.310 827.270 ;
        RECT 2800.730 826.090 2801.910 827.270 ;
        RECT 2799.130 824.490 2800.310 825.670 ;
        RECT 2800.730 824.490 2801.910 825.670 ;
        RECT 2799.130 646.090 2800.310 647.270 ;
        RECT 2800.730 646.090 2801.910 647.270 ;
        RECT 2799.130 644.490 2800.310 645.670 ;
        RECT 2800.730 644.490 2801.910 645.670 ;
        RECT 2799.130 466.090 2800.310 467.270 ;
        RECT 2800.730 466.090 2801.910 467.270 ;
        RECT 2799.130 464.490 2800.310 465.670 ;
        RECT 2800.730 464.490 2801.910 465.670 ;
        RECT 2799.130 286.090 2800.310 287.270 ;
        RECT 2800.730 286.090 2801.910 287.270 ;
        RECT 2799.130 284.490 2800.310 285.670 ;
        RECT 2800.730 284.490 2801.910 285.670 ;
        RECT 2799.130 106.090 2800.310 107.270 ;
        RECT 2800.730 106.090 2801.910 107.270 ;
        RECT 2799.130 104.490 2800.310 105.670 ;
        RECT 2800.730 104.490 2801.910 105.670 ;
        RECT 2799.130 -7.710 2800.310 -6.530 ;
        RECT 2800.730 -7.710 2801.910 -6.530 ;
        RECT 2799.130 -9.310 2800.310 -8.130 ;
        RECT 2800.730 -9.310 2801.910 -8.130 ;
        RECT 2931.510 3527.810 2932.690 3528.990 ;
        RECT 2933.110 3527.810 2934.290 3528.990 ;
        RECT 2931.510 3526.210 2932.690 3527.390 ;
        RECT 2933.110 3526.210 2934.290 3527.390 ;
        RECT 2931.510 3346.090 2932.690 3347.270 ;
        RECT 2933.110 3346.090 2934.290 3347.270 ;
        RECT 2931.510 3344.490 2932.690 3345.670 ;
        RECT 2933.110 3344.490 2934.290 3345.670 ;
        RECT 2931.510 3166.090 2932.690 3167.270 ;
        RECT 2933.110 3166.090 2934.290 3167.270 ;
        RECT 2931.510 3164.490 2932.690 3165.670 ;
        RECT 2933.110 3164.490 2934.290 3165.670 ;
        RECT 2931.510 2986.090 2932.690 2987.270 ;
        RECT 2933.110 2986.090 2934.290 2987.270 ;
        RECT 2931.510 2984.490 2932.690 2985.670 ;
        RECT 2933.110 2984.490 2934.290 2985.670 ;
        RECT 2931.510 2806.090 2932.690 2807.270 ;
        RECT 2933.110 2806.090 2934.290 2807.270 ;
        RECT 2931.510 2804.490 2932.690 2805.670 ;
        RECT 2933.110 2804.490 2934.290 2805.670 ;
        RECT 2931.510 2626.090 2932.690 2627.270 ;
        RECT 2933.110 2626.090 2934.290 2627.270 ;
        RECT 2931.510 2624.490 2932.690 2625.670 ;
        RECT 2933.110 2624.490 2934.290 2625.670 ;
        RECT 2931.510 2446.090 2932.690 2447.270 ;
        RECT 2933.110 2446.090 2934.290 2447.270 ;
        RECT 2931.510 2444.490 2932.690 2445.670 ;
        RECT 2933.110 2444.490 2934.290 2445.670 ;
        RECT 2931.510 2266.090 2932.690 2267.270 ;
        RECT 2933.110 2266.090 2934.290 2267.270 ;
        RECT 2931.510 2264.490 2932.690 2265.670 ;
        RECT 2933.110 2264.490 2934.290 2265.670 ;
        RECT 2931.510 2086.090 2932.690 2087.270 ;
        RECT 2933.110 2086.090 2934.290 2087.270 ;
        RECT 2931.510 2084.490 2932.690 2085.670 ;
        RECT 2933.110 2084.490 2934.290 2085.670 ;
        RECT 2931.510 1906.090 2932.690 1907.270 ;
        RECT 2933.110 1906.090 2934.290 1907.270 ;
        RECT 2931.510 1904.490 2932.690 1905.670 ;
        RECT 2933.110 1904.490 2934.290 1905.670 ;
        RECT 2931.510 1726.090 2932.690 1727.270 ;
        RECT 2933.110 1726.090 2934.290 1727.270 ;
        RECT 2931.510 1724.490 2932.690 1725.670 ;
        RECT 2933.110 1724.490 2934.290 1725.670 ;
        RECT 2931.510 1546.090 2932.690 1547.270 ;
        RECT 2933.110 1546.090 2934.290 1547.270 ;
        RECT 2931.510 1544.490 2932.690 1545.670 ;
        RECT 2933.110 1544.490 2934.290 1545.670 ;
        RECT 2931.510 1366.090 2932.690 1367.270 ;
        RECT 2933.110 1366.090 2934.290 1367.270 ;
        RECT 2931.510 1364.490 2932.690 1365.670 ;
        RECT 2933.110 1364.490 2934.290 1365.670 ;
        RECT 2931.510 1186.090 2932.690 1187.270 ;
        RECT 2933.110 1186.090 2934.290 1187.270 ;
        RECT 2931.510 1184.490 2932.690 1185.670 ;
        RECT 2933.110 1184.490 2934.290 1185.670 ;
        RECT 2931.510 1006.090 2932.690 1007.270 ;
        RECT 2933.110 1006.090 2934.290 1007.270 ;
        RECT 2931.510 1004.490 2932.690 1005.670 ;
        RECT 2933.110 1004.490 2934.290 1005.670 ;
        RECT 2931.510 826.090 2932.690 827.270 ;
        RECT 2933.110 826.090 2934.290 827.270 ;
        RECT 2931.510 824.490 2932.690 825.670 ;
        RECT 2933.110 824.490 2934.290 825.670 ;
        RECT 2931.510 646.090 2932.690 647.270 ;
        RECT 2933.110 646.090 2934.290 647.270 ;
        RECT 2931.510 644.490 2932.690 645.670 ;
        RECT 2933.110 644.490 2934.290 645.670 ;
        RECT 2931.510 466.090 2932.690 467.270 ;
        RECT 2933.110 466.090 2934.290 467.270 ;
        RECT 2931.510 464.490 2932.690 465.670 ;
        RECT 2933.110 464.490 2934.290 465.670 ;
        RECT 2931.510 286.090 2932.690 287.270 ;
        RECT 2933.110 286.090 2934.290 287.270 ;
        RECT 2931.510 284.490 2932.690 285.670 ;
        RECT 2933.110 284.490 2934.290 285.670 ;
        RECT 2931.510 106.090 2932.690 107.270 ;
        RECT 2933.110 106.090 2934.290 107.270 ;
        RECT 2931.510 104.490 2932.690 105.670 ;
        RECT 2933.110 104.490 2934.290 105.670 ;
        RECT 2931.510 -7.710 2932.690 -6.530 ;
        RECT 2933.110 -7.710 2934.290 -6.530 ;
        RECT 2931.510 -9.310 2932.690 -8.130 ;
        RECT 2933.110 -9.310 2934.290 -8.130 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
        RECT -14.830 824.330 2934.450 827.430 ;
        RECT -14.830 644.330 2934.450 647.430 ;
        RECT -14.830 464.330 2934.450 467.430 ;
        RECT -14.830 284.330 2934.450 287.430 ;
        RECT -14.830 104.330 2934.450 107.430 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
        RECT 297.570 1010.000 300.670 3538.750 ;
        RECT 477.570 1010.000 480.670 3538.750 ;
        RECT 657.570 1010.000 660.670 3538.750 ;
        RECT 837.570 1010.000 840.670 3538.750 ;
        RECT 1017.570 1010.000 1020.670 3538.750 ;
        RECT 297.570 -19.070 300.670 390.000 ;
        RECT 477.570 -19.070 480.670 390.000 ;
        RECT 657.570 -19.070 660.670 390.000 ;
        RECT 837.570 -19.070 840.670 390.000 ;
        RECT 1017.570 -19.070 1020.670 390.000 ;
        RECT 1197.570 -19.070 1200.670 3538.750 ;
        RECT 1377.570 -19.070 1380.670 3538.750 ;
        RECT 1557.570 -19.070 1560.670 3538.750 ;
        RECT 1737.570 -19.070 1740.670 3538.750 ;
        RECT 1917.570 -19.070 1920.670 3538.750 ;
        RECT 2097.570 -19.070 2100.670 3538.750 ;
        RECT 2277.570 -19.070 2280.670 3538.750 ;
        RECT 2457.570 -19.070 2460.670 3538.750 ;
        RECT 2637.570 -19.070 2640.670 3538.750 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER via4 ;
        RECT -24.270 3537.410 -23.090 3538.590 ;
        RECT -22.670 3537.410 -21.490 3538.590 ;
        RECT -24.270 3535.810 -23.090 3536.990 ;
        RECT -22.670 3535.810 -21.490 3536.990 ;
        RECT -24.270 3364.690 -23.090 3365.870 ;
        RECT -22.670 3364.690 -21.490 3365.870 ;
        RECT -24.270 3363.090 -23.090 3364.270 ;
        RECT -22.670 3363.090 -21.490 3364.270 ;
        RECT -24.270 3184.690 -23.090 3185.870 ;
        RECT -22.670 3184.690 -21.490 3185.870 ;
        RECT -24.270 3183.090 -23.090 3184.270 ;
        RECT -22.670 3183.090 -21.490 3184.270 ;
        RECT -24.270 3004.690 -23.090 3005.870 ;
        RECT -22.670 3004.690 -21.490 3005.870 ;
        RECT -24.270 3003.090 -23.090 3004.270 ;
        RECT -22.670 3003.090 -21.490 3004.270 ;
        RECT -24.270 2824.690 -23.090 2825.870 ;
        RECT -22.670 2824.690 -21.490 2825.870 ;
        RECT -24.270 2823.090 -23.090 2824.270 ;
        RECT -22.670 2823.090 -21.490 2824.270 ;
        RECT -24.270 2644.690 -23.090 2645.870 ;
        RECT -22.670 2644.690 -21.490 2645.870 ;
        RECT -24.270 2643.090 -23.090 2644.270 ;
        RECT -22.670 2643.090 -21.490 2644.270 ;
        RECT -24.270 2464.690 -23.090 2465.870 ;
        RECT -22.670 2464.690 -21.490 2465.870 ;
        RECT -24.270 2463.090 -23.090 2464.270 ;
        RECT -22.670 2463.090 -21.490 2464.270 ;
        RECT -24.270 2284.690 -23.090 2285.870 ;
        RECT -22.670 2284.690 -21.490 2285.870 ;
        RECT -24.270 2283.090 -23.090 2284.270 ;
        RECT -22.670 2283.090 -21.490 2284.270 ;
        RECT -24.270 2104.690 -23.090 2105.870 ;
        RECT -22.670 2104.690 -21.490 2105.870 ;
        RECT -24.270 2103.090 -23.090 2104.270 ;
        RECT -22.670 2103.090 -21.490 2104.270 ;
        RECT -24.270 1924.690 -23.090 1925.870 ;
        RECT -22.670 1924.690 -21.490 1925.870 ;
        RECT -24.270 1923.090 -23.090 1924.270 ;
        RECT -22.670 1923.090 -21.490 1924.270 ;
        RECT -24.270 1744.690 -23.090 1745.870 ;
        RECT -22.670 1744.690 -21.490 1745.870 ;
        RECT -24.270 1743.090 -23.090 1744.270 ;
        RECT -22.670 1743.090 -21.490 1744.270 ;
        RECT -24.270 1564.690 -23.090 1565.870 ;
        RECT -22.670 1564.690 -21.490 1565.870 ;
        RECT -24.270 1563.090 -23.090 1564.270 ;
        RECT -22.670 1563.090 -21.490 1564.270 ;
        RECT -24.270 1384.690 -23.090 1385.870 ;
        RECT -22.670 1384.690 -21.490 1385.870 ;
        RECT -24.270 1383.090 -23.090 1384.270 ;
        RECT -22.670 1383.090 -21.490 1384.270 ;
        RECT -24.270 1204.690 -23.090 1205.870 ;
        RECT -22.670 1204.690 -21.490 1205.870 ;
        RECT -24.270 1203.090 -23.090 1204.270 ;
        RECT -22.670 1203.090 -21.490 1204.270 ;
        RECT -24.270 1024.690 -23.090 1025.870 ;
        RECT -22.670 1024.690 -21.490 1025.870 ;
        RECT -24.270 1023.090 -23.090 1024.270 ;
        RECT -22.670 1023.090 -21.490 1024.270 ;
        RECT -24.270 844.690 -23.090 845.870 ;
        RECT -22.670 844.690 -21.490 845.870 ;
        RECT -24.270 843.090 -23.090 844.270 ;
        RECT -22.670 843.090 -21.490 844.270 ;
        RECT -24.270 664.690 -23.090 665.870 ;
        RECT -22.670 664.690 -21.490 665.870 ;
        RECT -24.270 663.090 -23.090 664.270 ;
        RECT -22.670 663.090 -21.490 664.270 ;
        RECT -24.270 484.690 -23.090 485.870 ;
        RECT -22.670 484.690 -21.490 485.870 ;
        RECT -24.270 483.090 -23.090 484.270 ;
        RECT -22.670 483.090 -21.490 484.270 ;
        RECT -24.270 304.690 -23.090 305.870 ;
        RECT -22.670 304.690 -21.490 305.870 ;
        RECT -24.270 303.090 -23.090 304.270 ;
        RECT -22.670 303.090 -21.490 304.270 ;
        RECT -24.270 124.690 -23.090 125.870 ;
        RECT -22.670 124.690 -21.490 125.870 ;
        RECT -24.270 123.090 -23.090 124.270 ;
        RECT -22.670 123.090 -21.490 124.270 ;
        RECT -24.270 -17.310 -23.090 -16.130 ;
        RECT -22.670 -17.310 -21.490 -16.130 ;
        RECT -24.270 -18.910 -23.090 -17.730 ;
        RECT -22.670 -18.910 -21.490 -17.730 ;
        RECT 117.730 3537.410 118.910 3538.590 ;
        RECT 119.330 3537.410 120.510 3538.590 ;
        RECT 117.730 3535.810 118.910 3536.990 ;
        RECT 119.330 3535.810 120.510 3536.990 ;
        RECT 117.730 3364.690 118.910 3365.870 ;
        RECT 119.330 3364.690 120.510 3365.870 ;
        RECT 117.730 3363.090 118.910 3364.270 ;
        RECT 119.330 3363.090 120.510 3364.270 ;
        RECT 117.730 3184.690 118.910 3185.870 ;
        RECT 119.330 3184.690 120.510 3185.870 ;
        RECT 117.730 3183.090 118.910 3184.270 ;
        RECT 119.330 3183.090 120.510 3184.270 ;
        RECT 117.730 3004.690 118.910 3005.870 ;
        RECT 119.330 3004.690 120.510 3005.870 ;
        RECT 117.730 3003.090 118.910 3004.270 ;
        RECT 119.330 3003.090 120.510 3004.270 ;
        RECT 117.730 2824.690 118.910 2825.870 ;
        RECT 119.330 2824.690 120.510 2825.870 ;
        RECT 117.730 2823.090 118.910 2824.270 ;
        RECT 119.330 2823.090 120.510 2824.270 ;
        RECT 117.730 2644.690 118.910 2645.870 ;
        RECT 119.330 2644.690 120.510 2645.870 ;
        RECT 117.730 2643.090 118.910 2644.270 ;
        RECT 119.330 2643.090 120.510 2644.270 ;
        RECT 117.730 2464.690 118.910 2465.870 ;
        RECT 119.330 2464.690 120.510 2465.870 ;
        RECT 117.730 2463.090 118.910 2464.270 ;
        RECT 119.330 2463.090 120.510 2464.270 ;
        RECT 117.730 2284.690 118.910 2285.870 ;
        RECT 119.330 2284.690 120.510 2285.870 ;
        RECT 117.730 2283.090 118.910 2284.270 ;
        RECT 119.330 2283.090 120.510 2284.270 ;
        RECT 117.730 2104.690 118.910 2105.870 ;
        RECT 119.330 2104.690 120.510 2105.870 ;
        RECT 117.730 2103.090 118.910 2104.270 ;
        RECT 119.330 2103.090 120.510 2104.270 ;
        RECT 117.730 1924.690 118.910 1925.870 ;
        RECT 119.330 1924.690 120.510 1925.870 ;
        RECT 117.730 1923.090 118.910 1924.270 ;
        RECT 119.330 1923.090 120.510 1924.270 ;
        RECT 117.730 1744.690 118.910 1745.870 ;
        RECT 119.330 1744.690 120.510 1745.870 ;
        RECT 117.730 1743.090 118.910 1744.270 ;
        RECT 119.330 1743.090 120.510 1744.270 ;
        RECT 117.730 1564.690 118.910 1565.870 ;
        RECT 119.330 1564.690 120.510 1565.870 ;
        RECT 117.730 1563.090 118.910 1564.270 ;
        RECT 119.330 1563.090 120.510 1564.270 ;
        RECT 117.730 1384.690 118.910 1385.870 ;
        RECT 119.330 1384.690 120.510 1385.870 ;
        RECT 117.730 1383.090 118.910 1384.270 ;
        RECT 119.330 1383.090 120.510 1384.270 ;
        RECT 117.730 1204.690 118.910 1205.870 ;
        RECT 119.330 1204.690 120.510 1205.870 ;
        RECT 117.730 1203.090 118.910 1204.270 ;
        RECT 119.330 1203.090 120.510 1204.270 ;
        RECT 117.730 1024.690 118.910 1025.870 ;
        RECT 119.330 1024.690 120.510 1025.870 ;
        RECT 117.730 1023.090 118.910 1024.270 ;
        RECT 119.330 1023.090 120.510 1024.270 ;
        RECT 297.730 3537.410 298.910 3538.590 ;
        RECT 299.330 3537.410 300.510 3538.590 ;
        RECT 297.730 3535.810 298.910 3536.990 ;
        RECT 299.330 3535.810 300.510 3536.990 ;
        RECT 297.730 3364.690 298.910 3365.870 ;
        RECT 299.330 3364.690 300.510 3365.870 ;
        RECT 297.730 3363.090 298.910 3364.270 ;
        RECT 299.330 3363.090 300.510 3364.270 ;
        RECT 297.730 3184.690 298.910 3185.870 ;
        RECT 299.330 3184.690 300.510 3185.870 ;
        RECT 297.730 3183.090 298.910 3184.270 ;
        RECT 299.330 3183.090 300.510 3184.270 ;
        RECT 297.730 3004.690 298.910 3005.870 ;
        RECT 299.330 3004.690 300.510 3005.870 ;
        RECT 297.730 3003.090 298.910 3004.270 ;
        RECT 299.330 3003.090 300.510 3004.270 ;
        RECT 297.730 2824.690 298.910 2825.870 ;
        RECT 299.330 2824.690 300.510 2825.870 ;
        RECT 297.730 2823.090 298.910 2824.270 ;
        RECT 299.330 2823.090 300.510 2824.270 ;
        RECT 297.730 2644.690 298.910 2645.870 ;
        RECT 299.330 2644.690 300.510 2645.870 ;
        RECT 297.730 2643.090 298.910 2644.270 ;
        RECT 299.330 2643.090 300.510 2644.270 ;
        RECT 297.730 2464.690 298.910 2465.870 ;
        RECT 299.330 2464.690 300.510 2465.870 ;
        RECT 297.730 2463.090 298.910 2464.270 ;
        RECT 299.330 2463.090 300.510 2464.270 ;
        RECT 297.730 2284.690 298.910 2285.870 ;
        RECT 299.330 2284.690 300.510 2285.870 ;
        RECT 297.730 2283.090 298.910 2284.270 ;
        RECT 299.330 2283.090 300.510 2284.270 ;
        RECT 297.730 2104.690 298.910 2105.870 ;
        RECT 299.330 2104.690 300.510 2105.870 ;
        RECT 297.730 2103.090 298.910 2104.270 ;
        RECT 299.330 2103.090 300.510 2104.270 ;
        RECT 297.730 1924.690 298.910 1925.870 ;
        RECT 299.330 1924.690 300.510 1925.870 ;
        RECT 297.730 1923.090 298.910 1924.270 ;
        RECT 299.330 1923.090 300.510 1924.270 ;
        RECT 297.730 1744.690 298.910 1745.870 ;
        RECT 299.330 1744.690 300.510 1745.870 ;
        RECT 297.730 1743.090 298.910 1744.270 ;
        RECT 299.330 1743.090 300.510 1744.270 ;
        RECT 297.730 1564.690 298.910 1565.870 ;
        RECT 299.330 1564.690 300.510 1565.870 ;
        RECT 297.730 1563.090 298.910 1564.270 ;
        RECT 299.330 1563.090 300.510 1564.270 ;
        RECT 297.730 1384.690 298.910 1385.870 ;
        RECT 299.330 1384.690 300.510 1385.870 ;
        RECT 297.730 1383.090 298.910 1384.270 ;
        RECT 299.330 1383.090 300.510 1384.270 ;
        RECT 297.730 1204.690 298.910 1205.870 ;
        RECT 299.330 1204.690 300.510 1205.870 ;
        RECT 297.730 1203.090 298.910 1204.270 ;
        RECT 299.330 1203.090 300.510 1204.270 ;
        RECT 297.730 1024.690 298.910 1025.870 ;
        RECT 299.330 1024.690 300.510 1025.870 ;
        RECT 297.730 1023.090 298.910 1024.270 ;
        RECT 299.330 1023.090 300.510 1024.270 ;
        RECT 477.730 3537.410 478.910 3538.590 ;
        RECT 479.330 3537.410 480.510 3538.590 ;
        RECT 477.730 3535.810 478.910 3536.990 ;
        RECT 479.330 3535.810 480.510 3536.990 ;
        RECT 477.730 3364.690 478.910 3365.870 ;
        RECT 479.330 3364.690 480.510 3365.870 ;
        RECT 477.730 3363.090 478.910 3364.270 ;
        RECT 479.330 3363.090 480.510 3364.270 ;
        RECT 477.730 3184.690 478.910 3185.870 ;
        RECT 479.330 3184.690 480.510 3185.870 ;
        RECT 477.730 3183.090 478.910 3184.270 ;
        RECT 479.330 3183.090 480.510 3184.270 ;
        RECT 477.730 3004.690 478.910 3005.870 ;
        RECT 479.330 3004.690 480.510 3005.870 ;
        RECT 477.730 3003.090 478.910 3004.270 ;
        RECT 479.330 3003.090 480.510 3004.270 ;
        RECT 477.730 2824.690 478.910 2825.870 ;
        RECT 479.330 2824.690 480.510 2825.870 ;
        RECT 477.730 2823.090 478.910 2824.270 ;
        RECT 479.330 2823.090 480.510 2824.270 ;
        RECT 477.730 2644.690 478.910 2645.870 ;
        RECT 479.330 2644.690 480.510 2645.870 ;
        RECT 477.730 2643.090 478.910 2644.270 ;
        RECT 479.330 2643.090 480.510 2644.270 ;
        RECT 477.730 2464.690 478.910 2465.870 ;
        RECT 479.330 2464.690 480.510 2465.870 ;
        RECT 477.730 2463.090 478.910 2464.270 ;
        RECT 479.330 2463.090 480.510 2464.270 ;
        RECT 477.730 2284.690 478.910 2285.870 ;
        RECT 479.330 2284.690 480.510 2285.870 ;
        RECT 477.730 2283.090 478.910 2284.270 ;
        RECT 479.330 2283.090 480.510 2284.270 ;
        RECT 477.730 2104.690 478.910 2105.870 ;
        RECT 479.330 2104.690 480.510 2105.870 ;
        RECT 477.730 2103.090 478.910 2104.270 ;
        RECT 479.330 2103.090 480.510 2104.270 ;
        RECT 477.730 1924.690 478.910 1925.870 ;
        RECT 479.330 1924.690 480.510 1925.870 ;
        RECT 477.730 1923.090 478.910 1924.270 ;
        RECT 479.330 1923.090 480.510 1924.270 ;
        RECT 477.730 1744.690 478.910 1745.870 ;
        RECT 479.330 1744.690 480.510 1745.870 ;
        RECT 477.730 1743.090 478.910 1744.270 ;
        RECT 479.330 1743.090 480.510 1744.270 ;
        RECT 477.730 1564.690 478.910 1565.870 ;
        RECT 479.330 1564.690 480.510 1565.870 ;
        RECT 477.730 1563.090 478.910 1564.270 ;
        RECT 479.330 1563.090 480.510 1564.270 ;
        RECT 477.730 1384.690 478.910 1385.870 ;
        RECT 479.330 1384.690 480.510 1385.870 ;
        RECT 477.730 1383.090 478.910 1384.270 ;
        RECT 479.330 1383.090 480.510 1384.270 ;
        RECT 477.730 1204.690 478.910 1205.870 ;
        RECT 479.330 1204.690 480.510 1205.870 ;
        RECT 477.730 1203.090 478.910 1204.270 ;
        RECT 479.330 1203.090 480.510 1204.270 ;
        RECT 477.730 1024.690 478.910 1025.870 ;
        RECT 479.330 1024.690 480.510 1025.870 ;
        RECT 477.730 1023.090 478.910 1024.270 ;
        RECT 479.330 1023.090 480.510 1024.270 ;
        RECT 657.730 3537.410 658.910 3538.590 ;
        RECT 659.330 3537.410 660.510 3538.590 ;
        RECT 657.730 3535.810 658.910 3536.990 ;
        RECT 659.330 3535.810 660.510 3536.990 ;
        RECT 657.730 3364.690 658.910 3365.870 ;
        RECT 659.330 3364.690 660.510 3365.870 ;
        RECT 657.730 3363.090 658.910 3364.270 ;
        RECT 659.330 3363.090 660.510 3364.270 ;
        RECT 657.730 3184.690 658.910 3185.870 ;
        RECT 659.330 3184.690 660.510 3185.870 ;
        RECT 657.730 3183.090 658.910 3184.270 ;
        RECT 659.330 3183.090 660.510 3184.270 ;
        RECT 657.730 3004.690 658.910 3005.870 ;
        RECT 659.330 3004.690 660.510 3005.870 ;
        RECT 657.730 3003.090 658.910 3004.270 ;
        RECT 659.330 3003.090 660.510 3004.270 ;
        RECT 657.730 2824.690 658.910 2825.870 ;
        RECT 659.330 2824.690 660.510 2825.870 ;
        RECT 657.730 2823.090 658.910 2824.270 ;
        RECT 659.330 2823.090 660.510 2824.270 ;
        RECT 657.730 2644.690 658.910 2645.870 ;
        RECT 659.330 2644.690 660.510 2645.870 ;
        RECT 657.730 2643.090 658.910 2644.270 ;
        RECT 659.330 2643.090 660.510 2644.270 ;
        RECT 657.730 2464.690 658.910 2465.870 ;
        RECT 659.330 2464.690 660.510 2465.870 ;
        RECT 657.730 2463.090 658.910 2464.270 ;
        RECT 659.330 2463.090 660.510 2464.270 ;
        RECT 657.730 2284.690 658.910 2285.870 ;
        RECT 659.330 2284.690 660.510 2285.870 ;
        RECT 657.730 2283.090 658.910 2284.270 ;
        RECT 659.330 2283.090 660.510 2284.270 ;
        RECT 657.730 2104.690 658.910 2105.870 ;
        RECT 659.330 2104.690 660.510 2105.870 ;
        RECT 657.730 2103.090 658.910 2104.270 ;
        RECT 659.330 2103.090 660.510 2104.270 ;
        RECT 657.730 1924.690 658.910 1925.870 ;
        RECT 659.330 1924.690 660.510 1925.870 ;
        RECT 657.730 1923.090 658.910 1924.270 ;
        RECT 659.330 1923.090 660.510 1924.270 ;
        RECT 657.730 1744.690 658.910 1745.870 ;
        RECT 659.330 1744.690 660.510 1745.870 ;
        RECT 657.730 1743.090 658.910 1744.270 ;
        RECT 659.330 1743.090 660.510 1744.270 ;
        RECT 657.730 1564.690 658.910 1565.870 ;
        RECT 659.330 1564.690 660.510 1565.870 ;
        RECT 657.730 1563.090 658.910 1564.270 ;
        RECT 659.330 1563.090 660.510 1564.270 ;
        RECT 657.730 1384.690 658.910 1385.870 ;
        RECT 659.330 1384.690 660.510 1385.870 ;
        RECT 657.730 1383.090 658.910 1384.270 ;
        RECT 659.330 1383.090 660.510 1384.270 ;
        RECT 657.730 1204.690 658.910 1205.870 ;
        RECT 659.330 1204.690 660.510 1205.870 ;
        RECT 657.730 1203.090 658.910 1204.270 ;
        RECT 659.330 1203.090 660.510 1204.270 ;
        RECT 657.730 1024.690 658.910 1025.870 ;
        RECT 659.330 1024.690 660.510 1025.870 ;
        RECT 657.730 1023.090 658.910 1024.270 ;
        RECT 659.330 1023.090 660.510 1024.270 ;
        RECT 837.730 3537.410 838.910 3538.590 ;
        RECT 839.330 3537.410 840.510 3538.590 ;
        RECT 837.730 3535.810 838.910 3536.990 ;
        RECT 839.330 3535.810 840.510 3536.990 ;
        RECT 837.730 3364.690 838.910 3365.870 ;
        RECT 839.330 3364.690 840.510 3365.870 ;
        RECT 837.730 3363.090 838.910 3364.270 ;
        RECT 839.330 3363.090 840.510 3364.270 ;
        RECT 837.730 3184.690 838.910 3185.870 ;
        RECT 839.330 3184.690 840.510 3185.870 ;
        RECT 837.730 3183.090 838.910 3184.270 ;
        RECT 839.330 3183.090 840.510 3184.270 ;
        RECT 837.730 3004.690 838.910 3005.870 ;
        RECT 839.330 3004.690 840.510 3005.870 ;
        RECT 837.730 3003.090 838.910 3004.270 ;
        RECT 839.330 3003.090 840.510 3004.270 ;
        RECT 837.730 2824.690 838.910 2825.870 ;
        RECT 839.330 2824.690 840.510 2825.870 ;
        RECT 837.730 2823.090 838.910 2824.270 ;
        RECT 839.330 2823.090 840.510 2824.270 ;
        RECT 837.730 2644.690 838.910 2645.870 ;
        RECT 839.330 2644.690 840.510 2645.870 ;
        RECT 837.730 2643.090 838.910 2644.270 ;
        RECT 839.330 2643.090 840.510 2644.270 ;
        RECT 837.730 2464.690 838.910 2465.870 ;
        RECT 839.330 2464.690 840.510 2465.870 ;
        RECT 837.730 2463.090 838.910 2464.270 ;
        RECT 839.330 2463.090 840.510 2464.270 ;
        RECT 837.730 2284.690 838.910 2285.870 ;
        RECT 839.330 2284.690 840.510 2285.870 ;
        RECT 837.730 2283.090 838.910 2284.270 ;
        RECT 839.330 2283.090 840.510 2284.270 ;
        RECT 837.730 2104.690 838.910 2105.870 ;
        RECT 839.330 2104.690 840.510 2105.870 ;
        RECT 837.730 2103.090 838.910 2104.270 ;
        RECT 839.330 2103.090 840.510 2104.270 ;
        RECT 837.730 1924.690 838.910 1925.870 ;
        RECT 839.330 1924.690 840.510 1925.870 ;
        RECT 837.730 1923.090 838.910 1924.270 ;
        RECT 839.330 1923.090 840.510 1924.270 ;
        RECT 837.730 1744.690 838.910 1745.870 ;
        RECT 839.330 1744.690 840.510 1745.870 ;
        RECT 837.730 1743.090 838.910 1744.270 ;
        RECT 839.330 1743.090 840.510 1744.270 ;
        RECT 837.730 1564.690 838.910 1565.870 ;
        RECT 839.330 1564.690 840.510 1565.870 ;
        RECT 837.730 1563.090 838.910 1564.270 ;
        RECT 839.330 1563.090 840.510 1564.270 ;
        RECT 837.730 1384.690 838.910 1385.870 ;
        RECT 839.330 1384.690 840.510 1385.870 ;
        RECT 837.730 1383.090 838.910 1384.270 ;
        RECT 839.330 1383.090 840.510 1384.270 ;
        RECT 837.730 1204.690 838.910 1205.870 ;
        RECT 839.330 1204.690 840.510 1205.870 ;
        RECT 837.730 1203.090 838.910 1204.270 ;
        RECT 839.330 1203.090 840.510 1204.270 ;
        RECT 837.730 1024.690 838.910 1025.870 ;
        RECT 839.330 1024.690 840.510 1025.870 ;
        RECT 837.730 1023.090 838.910 1024.270 ;
        RECT 839.330 1023.090 840.510 1024.270 ;
        RECT 1017.730 3537.410 1018.910 3538.590 ;
        RECT 1019.330 3537.410 1020.510 3538.590 ;
        RECT 1017.730 3535.810 1018.910 3536.990 ;
        RECT 1019.330 3535.810 1020.510 3536.990 ;
        RECT 1017.730 3364.690 1018.910 3365.870 ;
        RECT 1019.330 3364.690 1020.510 3365.870 ;
        RECT 1017.730 3363.090 1018.910 3364.270 ;
        RECT 1019.330 3363.090 1020.510 3364.270 ;
        RECT 1017.730 3184.690 1018.910 3185.870 ;
        RECT 1019.330 3184.690 1020.510 3185.870 ;
        RECT 1017.730 3183.090 1018.910 3184.270 ;
        RECT 1019.330 3183.090 1020.510 3184.270 ;
        RECT 1017.730 3004.690 1018.910 3005.870 ;
        RECT 1019.330 3004.690 1020.510 3005.870 ;
        RECT 1017.730 3003.090 1018.910 3004.270 ;
        RECT 1019.330 3003.090 1020.510 3004.270 ;
        RECT 1017.730 2824.690 1018.910 2825.870 ;
        RECT 1019.330 2824.690 1020.510 2825.870 ;
        RECT 1017.730 2823.090 1018.910 2824.270 ;
        RECT 1019.330 2823.090 1020.510 2824.270 ;
        RECT 1017.730 2644.690 1018.910 2645.870 ;
        RECT 1019.330 2644.690 1020.510 2645.870 ;
        RECT 1017.730 2643.090 1018.910 2644.270 ;
        RECT 1019.330 2643.090 1020.510 2644.270 ;
        RECT 1017.730 2464.690 1018.910 2465.870 ;
        RECT 1019.330 2464.690 1020.510 2465.870 ;
        RECT 1017.730 2463.090 1018.910 2464.270 ;
        RECT 1019.330 2463.090 1020.510 2464.270 ;
        RECT 1017.730 2284.690 1018.910 2285.870 ;
        RECT 1019.330 2284.690 1020.510 2285.870 ;
        RECT 1017.730 2283.090 1018.910 2284.270 ;
        RECT 1019.330 2283.090 1020.510 2284.270 ;
        RECT 1017.730 2104.690 1018.910 2105.870 ;
        RECT 1019.330 2104.690 1020.510 2105.870 ;
        RECT 1017.730 2103.090 1018.910 2104.270 ;
        RECT 1019.330 2103.090 1020.510 2104.270 ;
        RECT 1017.730 1924.690 1018.910 1925.870 ;
        RECT 1019.330 1924.690 1020.510 1925.870 ;
        RECT 1017.730 1923.090 1018.910 1924.270 ;
        RECT 1019.330 1923.090 1020.510 1924.270 ;
        RECT 1017.730 1744.690 1018.910 1745.870 ;
        RECT 1019.330 1744.690 1020.510 1745.870 ;
        RECT 1017.730 1743.090 1018.910 1744.270 ;
        RECT 1019.330 1743.090 1020.510 1744.270 ;
        RECT 1017.730 1564.690 1018.910 1565.870 ;
        RECT 1019.330 1564.690 1020.510 1565.870 ;
        RECT 1017.730 1563.090 1018.910 1564.270 ;
        RECT 1019.330 1563.090 1020.510 1564.270 ;
        RECT 1017.730 1384.690 1018.910 1385.870 ;
        RECT 1019.330 1384.690 1020.510 1385.870 ;
        RECT 1017.730 1383.090 1018.910 1384.270 ;
        RECT 1019.330 1383.090 1020.510 1384.270 ;
        RECT 1017.730 1204.690 1018.910 1205.870 ;
        RECT 1019.330 1204.690 1020.510 1205.870 ;
        RECT 1017.730 1203.090 1018.910 1204.270 ;
        RECT 1019.330 1203.090 1020.510 1204.270 ;
        RECT 1017.730 1024.690 1018.910 1025.870 ;
        RECT 1019.330 1024.690 1020.510 1025.870 ;
        RECT 1017.730 1023.090 1018.910 1024.270 ;
        RECT 1019.330 1023.090 1020.510 1024.270 ;
        RECT 1197.730 3537.410 1198.910 3538.590 ;
        RECT 1199.330 3537.410 1200.510 3538.590 ;
        RECT 1197.730 3535.810 1198.910 3536.990 ;
        RECT 1199.330 3535.810 1200.510 3536.990 ;
        RECT 1197.730 3364.690 1198.910 3365.870 ;
        RECT 1199.330 3364.690 1200.510 3365.870 ;
        RECT 1197.730 3363.090 1198.910 3364.270 ;
        RECT 1199.330 3363.090 1200.510 3364.270 ;
        RECT 1197.730 3184.690 1198.910 3185.870 ;
        RECT 1199.330 3184.690 1200.510 3185.870 ;
        RECT 1197.730 3183.090 1198.910 3184.270 ;
        RECT 1199.330 3183.090 1200.510 3184.270 ;
        RECT 1197.730 3004.690 1198.910 3005.870 ;
        RECT 1199.330 3004.690 1200.510 3005.870 ;
        RECT 1197.730 3003.090 1198.910 3004.270 ;
        RECT 1199.330 3003.090 1200.510 3004.270 ;
        RECT 1197.730 2824.690 1198.910 2825.870 ;
        RECT 1199.330 2824.690 1200.510 2825.870 ;
        RECT 1197.730 2823.090 1198.910 2824.270 ;
        RECT 1199.330 2823.090 1200.510 2824.270 ;
        RECT 1197.730 2644.690 1198.910 2645.870 ;
        RECT 1199.330 2644.690 1200.510 2645.870 ;
        RECT 1197.730 2643.090 1198.910 2644.270 ;
        RECT 1199.330 2643.090 1200.510 2644.270 ;
        RECT 1197.730 2464.690 1198.910 2465.870 ;
        RECT 1199.330 2464.690 1200.510 2465.870 ;
        RECT 1197.730 2463.090 1198.910 2464.270 ;
        RECT 1199.330 2463.090 1200.510 2464.270 ;
        RECT 1197.730 2284.690 1198.910 2285.870 ;
        RECT 1199.330 2284.690 1200.510 2285.870 ;
        RECT 1197.730 2283.090 1198.910 2284.270 ;
        RECT 1199.330 2283.090 1200.510 2284.270 ;
        RECT 1197.730 2104.690 1198.910 2105.870 ;
        RECT 1199.330 2104.690 1200.510 2105.870 ;
        RECT 1197.730 2103.090 1198.910 2104.270 ;
        RECT 1199.330 2103.090 1200.510 2104.270 ;
        RECT 1197.730 1924.690 1198.910 1925.870 ;
        RECT 1199.330 1924.690 1200.510 1925.870 ;
        RECT 1197.730 1923.090 1198.910 1924.270 ;
        RECT 1199.330 1923.090 1200.510 1924.270 ;
        RECT 1197.730 1744.690 1198.910 1745.870 ;
        RECT 1199.330 1744.690 1200.510 1745.870 ;
        RECT 1197.730 1743.090 1198.910 1744.270 ;
        RECT 1199.330 1743.090 1200.510 1744.270 ;
        RECT 1197.730 1564.690 1198.910 1565.870 ;
        RECT 1199.330 1564.690 1200.510 1565.870 ;
        RECT 1197.730 1563.090 1198.910 1564.270 ;
        RECT 1199.330 1563.090 1200.510 1564.270 ;
        RECT 1197.730 1384.690 1198.910 1385.870 ;
        RECT 1199.330 1384.690 1200.510 1385.870 ;
        RECT 1197.730 1383.090 1198.910 1384.270 ;
        RECT 1199.330 1383.090 1200.510 1384.270 ;
        RECT 1197.730 1204.690 1198.910 1205.870 ;
        RECT 1199.330 1204.690 1200.510 1205.870 ;
        RECT 1197.730 1203.090 1198.910 1204.270 ;
        RECT 1199.330 1203.090 1200.510 1204.270 ;
        RECT 1197.730 1024.690 1198.910 1025.870 ;
        RECT 1199.330 1024.690 1200.510 1025.870 ;
        RECT 1197.730 1023.090 1198.910 1024.270 ;
        RECT 1199.330 1023.090 1200.510 1024.270 ;
        RECT 117.730 844.690 118.910 845.870 ;
        RECT 119.330 844.690 120.510 845.870 ;
        RECT 117.730 843.090 118.910 844.270 ;
        RECT 119.330 843.090 120.510 844.270 ;
        RECT 117.730 664.690 118.910 665.870 ;
        RECT 119.330 664.690 120.510 665.870 ;
        RECT 117.730 663.090 118.910 664.270 ;
        RECT 119.330 663.090 120.510 664.270 ;
        RECT 117.730 484.690 118.910 485.870 ;
        RECT 119.330 484.690 120.510 485.870 ;
        RECT 117.730 483.090 118.910 484.270 ;
        RECT 119.330 483.090 120.510 484.270 ;
        RECT 1197.730 844.690 1198.910 845.870 ;
        RECT 1199.330 844.690 1200.510 845.870 ;
        RECT 1197.730 843.090 1198.910 844.270 ;
        RECT 1199.330 843.090 1200.510 844.270 ;
        RECT 1197.730 664.690 1198.910 665.870 ;
        RECT 1199.330 664.690 1200.510 665.870 ;
        RECT 1197.730 663.090 1198.910 664.270 ;
        RECT 1199.330 663.090 1200.510 664.270 ;
        RECT 1197.730 484.690 1198.910 485.870 ;
        RECT 1199.330 484.690 1200.510 485.870 ;
        RECT 1197.730 483.090 1198.910 484.270 ;
        RECT 1199.330 483.090 1200.510 484.270 ;
        RECT 117.730 304.690 118.910 305.870 ;
        RECT 119.330 304.690 120.510 305.870 ;
        RECT 117.730 303.090 118.910 304.270 ;
        RECT 119.330 303.090 120.510 304.270 ;
        RECT 117.730 124.690 118.910 125.870 ;
        RECT 119.330 124.690 120.510 125.870 ;
        RECT 117.730 123.090 118.910 124.270 ;
        RECT 119.330 123.090 120.510 124.270 ;
        RECT 117.730 -17.310 118.910 -16.130 ;
        RECT 119.330 -17.310 120.510 -16.130 ;
        RECT 117.730 -18.910 118.910 -17.730 ;
        RECT 119.330 -18.910 120.510 -17.730 ;
        RECT 297.730 304.690 298.910 305.870 ;
        RECT 299.330 304.690 300.510 305.870 ;
        RECT 297.730 303.090 298.910 304.270 ;
        RECT 299.330 303.090 300.510 304.270 ;
        RECT 297.730 124.690 298.910 125.870 ;
        RECT 299.330 124.690 300.510 125.870 ;
        RECT 297.730 123.090 298.910 124.270 ;
        RECT 299.330 123.090 300.510 124.270 ;
        RECT 297.730 -17.310 298.910 -16.130 ;
        RECT 299.330 -17.310 300.510 -16.130 ;
        RECT 297.730 -18.910 298.910 -17.730 ;
        RECT 299.330 -18.910 300.510 -17.730 ;
        RECT 477.730 304.690 478.910 305.870 ;
        RECT 479.330 304.690 480.510 305.870 ;
        RECT 477.730 303.090 478.910 304.270 ;
        RECT 479.330 303.090 480.510 304.270 ;
        RECT 477.730 124.690 478.910 125.870 ;
        RECT 479.330 124.690 480.510 125.870 ;
        RECT 477.730 123.090 478.910 124.270 ;
        RECT 479.330 123.090 480.510 124.270 ;
        RECT 477.730 -17.310 478.910 -16.130 ;
        RECT 479.330 -17.310 480.510 -16.130 ;
        RECT 477.730 -18.910 478.910 -17.730 ;
        RECT 479.330 -18.910 480.510 -17.730 ;
        RECT 657.730 304.690 658.910 305.870 ;
        RECT 659.330 304.690 660.510 305.870 ;
        RECT 657.730 303.090 658.910 304.270 ;
        RECT 659.330 303.090 660.510 304.270 ;
        RECT 657.730 124.690 658.910 125.870 ;
        RECT 659.330 124.690 660.510 125.870 ;
        RECT 657.730 123.090 658.910 124.270 ;
        RECT 659.330 123.090 660.510 124.270 ;
        RECT 657.730 -17.310 658.910 -16.130 ;
        RECT 659.330 -17.310 660.510 -16.130 ;
        RECT 657.730 -18.910 658.910 -17.730 ;
        RECT 659.330 -18.910 660.510 -17.730 ;
        RECT 837.730 304.690 838.910 305.870 ;
        RECT 839.330 304.690 840.510 305.870 ;
        RECT 837.730 303.090 838.910 304.270 ;
        RECT 839.330 303.090 840.510 304.270 ;
        RECT 837.730 124.690 838.910 125.870 ;
        RECT 839.330 124.690 840.510 125.870 ;
        RECT 837.730 123.090 838.910 124.270 ;
        RECT 839.330 123.090 840.510 124.270 ;
        RECT 837.730 -17.310 838.910 -16.130 ;
        RECT 839.330 -17.310 840.510 -16.130 ;
        RECT 837.730 -18.910 838.910 -17.730 ;
        RECT 839.330 -18.910 840.510 -17.730 ;
        RECT 1017.730 304.690 1018.910 305.870 ;
        RECT 1019.330 304.690 1020.510 305.870 ;
        RECT 1017.730 303.090 1018.910 304.270 ;
        RECT 1019.330 303.090 1020.510 304.270 ;
        RECT 1017.730 124.690 1018.910 125.870 ;
        RECT 1019.330 124.690 1020.510 125.870 ;
        RECT 1017.730 123.090 1018.910 124.270 ;
        RECT 1019.330 123.090 1020.510 124.270 ;
        RECT 1017.730 -17.310 1018.910 -16.130 ;
        RECT 1019.330 -17.310 1020.510 -16.130 ;
        RECT 1017.730 -18.910 1018.910 -17.730 ;
        RECT 1019.330 -18.910 1020.510 -17.730 ;
        RECT 1197.730 304.690 1198.910 305.870 ;
        RECT 1199.330 304.690 1200.510 305.870 ;
        RECT 1197.730 303.090 1198.910 304.270 ;
        RECT 1199.330 303.090 1200.510 304.270 ;
        RECT 1197.730 124.690 1198.910 125.870 ;
        RECT 1199.330 124.690 1200.510 125.870 ;
        RECT 1197.730 123.090 1198.910 124.270 ;
        RECT 1199.330 123.090 1200.510 124.270 ;
        RECT 1197.730 -17.310 1198.910 -16.130 ;
        RECT 1199.330 -17.310 1200.510 -16.130 ;
        RECT 1197.730 -18.910 1198.910 -17.730 ;
        RECT 1199.330 -18.910 1200.510 -17.730 ;
        RECT 1377.730 3537.410 1378.910 3538.590 ;
        RECT 1379.330 3537.410 1380.510 3538.590 ;
        RECT 1377.730 3535.810 1378.910 3536.990 ;
        RECT 1379.330 3535.810 1380.510 3536.990 ;
        RECT 1377.730 3364.690 1378.910 3365.870 ;
        RECT 1379.330 3364.690 1380.510 3365.870 ;
        RECT 1377.730 3363.090 1378.910 3364.270 ;
        RECT 1379.330 3363.090 1380.510 3364.270 ;
        RECT 1377.730 3184.690 1378.910 3185.870 ;
        RECT 1379.330 3184.690 1380.510 3185.870 ;
        RECT 1377.730 3183.090 1378.910 3184.270 ;
        RECT 1379.330 3183.090 1380.510 3184.270 ;
        RECT 1377.730 3004.690 1378.910 3005.870 ;
        RECT 1379.330 3004.690 1380.510 3005.870 ;
        RECT 1377.730 3003.090 1378.910 3004.270 ;
        RECT 1379.330 3003.090 1380.510 3004.270 ;
        RECT 1377.730 2824.690 1378.910 2825.870 ;
        RECT 1379.330 2824.690 1380.510 2825.870 ;
        RECT 1377.730 2823.090 1378.910 2824.270 ;
        RECT 1379.330 2823.090 1380.510 2824.270 ;
        RECT 1377.730 2644.690 1378.910 2645.870 ;
        RECT 1379.330 2644.690 1380.510 2645.870 ;
        RECT 1377.730 2643.090 1378.910 2644.270 ;
        RECT 1379.330 2643.090 1380.510 2644.270 ;
        RECT 1377.730 2464.690 1378.910 2465.870 ;
        RECT 1379.330 2464.690 1380.510 2465.870 ;
        RECT 1377.730 2463.090 1378.910 2464.270 ;
        RECT 1379.330 2463.090 1380.510 2464.270 ;
        RECT 1377.730 2284.690 1378.910 2285.870 ;
        RECT 1379.330 2284.690 1380.510 2285.870 ;
        RECT 1377.730 2283.090 1378.910 2284.270 ;
        RECT 1379.330 2283.090 1380.510 2284.270 ;
        RECT 1377.730 2104.690 1378.910 2105.870 ;
        RECT 1379.330 2104.690 1380.510 2105.870 ;
        RECT 1377.730 2103.090 1378.910 2104.270 ;
        RECT 1379.330 2103.090 1380.510 2104.270 ;
        RECT 1377.730 1924.690 1378.910 1925.870 ;
        RECT 1379.330 1924.690 1380.510 1925.870 ;
        RECT 1377.730 1923.090 1378.910 1924.270 ;
        RECT 1379.330 1923.090 1380.510 1924.270 ;
        RECT 1377.730 1744.690 1378.910 1745.870 ;
        RECT 1379.330 1744.690 1380.510 1745.870 ;
        RECT 1377.730 1743.090 1378.910 1744.270 ;
        RECT 1379.330 1743.090 1380.510 1744.270 ;
        RECT 1377.730 1564.690 1378.910 1565.870 ;
        RECT 1379.330 1564.690 1380.510 1565.870 ;
        RECT 1377.730 1563.090 1378.910 1564.270 ;
        RECT 1379.330 1563.090 1380.510 1564.270 ;
        RECT 1377.730 1384.690 1378.910 1385.870 ;
        RECT 1379.330 1384.690 1380.510 1385.870 ;
        RECT 1377.730 1383.090 1378.910 1384.270 ;
        RECT 1379.330 1383.090 1380.510 1384.270 ;
        RECT 1377.730 1204.690 1378.910 1205.870 ;
        RECT 1379.330 1204.690 1380.510 1205.870 ;
        RECT 1377.730 1203.090 1378.910 1204.270 ;
        RECT 1379.330 1203.090 1380.510 1204.270 ;
        RECT 1377.730 1024.690 1378.910 1025.870 ;
        RECT 1379.330 1024.690 1380.510 1025.870 ;
        RECT 1377.730 1023.090 1378.910 1024.270 ;
        RECT 1379.330 1023.090 1380.510 1024.270 ;
        RECT 1377.730 844.690 1378.910 845.870 ;
        RECT 1379.330 844.690 1380.510 845.870 ;
        RECT 1377.730 843.090 1378.910 844.270 ;
        RECT 1379.330 843.090 1380.510 844.270 ;
        RECT 1377.730 664.690 1378.910 665.870 ;
        RECT 1379.330 664.690 1380.510 665.870 ;
        RECT 1377.730 663.090 1378.910 664.270 ;
        RECT 1379.330 663.090 1380.510 664.270 ;
        RECT 1377.730 484.690 1378.910 485.870 ;
        RECT 1379.330 484.690 1380.510 485.870 ;
        RECT 1377.730 483.090 1378.910 484.270 ;
        RECT 1379.330 483.090 1380.510 484.270 ;
        RECT 1377.730 304.690 1378.910 305.870 ;
        RECT 1379.330 304.690 1380.510 305.870 ;
        RECT 1377.730 303.090 1378.910 304.270 ;
        RECT 1379.330 303.090 1380.510 304.270 ;
        RECT 1377.730 124.690 1378.910 125.870 ;
        RECT 1379.330 124.690 1380.510 125.870 ;
        RECT 1377.730 123.090 1378.910 124.270 ;
        RECT 1379.330 123.090 1380.510 124.270 ;
        RECT 1377.730 -17.310 1378.910 -16.130 ;
        RECT 1379.330 -17.310 1380.510 -16.130 ;
        RECT 1377.730 -18.910 1378.910 -17.730 ;
        RECT 1379.330 -18.910 1380.510 -17.730 ;
        RECT 1557.730 3537.410 1558.910 3538.590 ;
        RECT 1559.330 3537.410 1560.510 3538.590 ;
        RECT 1557.730 3535.810 1558.910 3536.990 ;
        RECT 1559.330 3535.810 1560.510 3536.990 ;
        RECT 1557.730 3364.690 1558.910 3365.870 ;
        RECT 1559.330 3364.690 1560.510 3365.870 ;
        RECT 1557.730 3363.090 1558.910 3364.270 ;
        RECT 1559.330 3363.090 1560.510 3364.270 ;
        RECT 1557.730 3184.690 1558.910 3185.870 ;
        RECT 1559.330 3184.690 1560.510 3185.870 ;
        RECT 1557.730 3183.090 1558.910 3184.270 ;
        RECT 1559.330 3183.090 1560.510 3184.270 ;
        RECT 1557.730 3004.690 1558.910 3005.870 ;
        RECT 1559.330 3004.690 1560.510 3005.870 ;
        RECT 1557.730 3003.090 1558.910 3004.270 ;
        RECT 1559.330 3003.090 1560.510 3004.270 ;
        RECT 1557.730 2824.690 1558.910 2825.870 ;
        RECT 1559.330 2824.690 1560.510 2825.870 ;
        RECT 1557.730 2823.090 1558.910 2824.270 ;
        RECT 1559.330 2823.090 1560.510 2824.270 ;
        RECT 1557.730 2644.690 1558.910 2645.870 ;
        RECT 1559.330 2644.690 1560.510 2645.870 ;
        RECT 1557.730 2643.090 1558.910 2644.270 ;
        RECT 1559.330 2643.090 1560.510 2644.270 ;
        RECT 1557.730 2464.690 1558.910 2465.870 ;
        RECT 1559.330 2464.690 1560.510 2465.870 ;
        RECT 1557.730 2463.090 1558.910 2464.270 ;
        RECT 1559.330 2463.090 1560.510 2464.270 ;
        RECT 1557.730 2284.690 1558.910 2285.870 ;
        RECT 1559.330 2284.690 1560.510 2285.870 ;
        RECT 1557.730 2283.090 1558.910 2284.270 ;
        RECT 1559.330 2283.090 1560.510 2284.270 ;
        RECT 1557.730 2104.690 1558.910 2105.870 ;
        RECT 1559.330 2104.690 1560.510 2105.870 ;
        RECT 1557.730 2103.090 1558.910 2104.270 ;
        RECT 1559.330 2103.090 1560.510 2104.270 ;
        RECT 1557.730 1924.690 1558.910 1925.870 ;
        RECT 1559.330 1924.690 1560.510 1925.870 ;
        RECT 1557.730 1923.090 1558.910 1924.270 ;
        RECT 1559.330 1923.090 1560.510 1924.270 ;
        RECT 1557.730 1744.690 1558.910 1745.870 ;
        RECT 1559.330 1744.690 1560.510 1745.870 ;
        RECT 1557.730 1743.090 1558.910 1744.270 ;
        RECT 1559.330 1743.090 1560.510 1744.270 ;
        RECT 1557.730 1564.690 1558.910 1565.870 ;
        RECT 1559.330 1564.690 1560.510 1565.870 ;
        RECT 1557.730 1563.090 1558.910 1564.270 ;
        RECT 1559.330 1563.090 1560.510 1564.270 ;
        RECT 1557.730 1384.690 1558.910 1385.870 ;
        RECT 1559.330 1384.690 1560.510 1385.870 ;
        RECT 1557.730 1383.090 1558.910 1384.270 ;
        RECT 1559.330 1383.090 1560.510 1384.270 ;
        RECT 1557.730 1204.690 1558.910 1205.870 ;
        RECT 1559.330 1204.690 1560.510 1205.870 ;
        RECT 1557.730 1203.090 1558.910 1204.270 ;
        RECT 1559.330 1203.090 1560.510 1204.270 ;
        RECT 1557.730 1024.690 1558.910 1025.870 ;
        RECT 1559.330 1024.690 1560.510 1025.870 ;
        RECT 1557.730 1023.090 1558.910 1024.270 ;
        RECT 1559.330 1023.090 1560.510 1024.270 ;
        RECT 1557.730 844.690 1558.910 845.870 ;
        RECT 1559.330 844.690 1560.510 845.870 ;
        RECT 1557.730 843.090 1558.910 844.270 ;
        RECT 1559.330 843.090 1560.510 844.270 ;
        RECT 1557.730 664.690 1558.910 665.870 ;
        RECT 1559.330 664.690 1560.510 665.870 ;
        RECT 1557.730 663.090 1558.910 664.270 ;
        RECT 1559.330 663.090 1560.510 664.270 ;
        RECT 1557.730 484.690 1558.910 485.870 ;
        RECT 1559.330 484.690 1560.510 485.870 ;
        RECT 1557.730 483.090 1558.910 484.270 ;
        RECT 1559.330 483.090 1560.510 484.270 ;
        RECT 1557.730 304.690 1558.910 305.870 ;
        RECT 1559.330 304.690 1560.510 305.870 ;
        RECT 1557.730 303.090 1558.910 304.270 ;
        RECT 1559.330 303.090 1560.510 304.270 ;
        RECT 1557.730 124.690 1558.910 125.870 ;
        RECT 1559.330 124.690 1560.510 125.870 ;
        RECT 1557.730 123.090 1558.910 124.270 ;
        RECT 1559.330 123.090 1560.510 124.270 ;
        RECT 1557.730 -17.310 1558.910 -16.130 ;
        RECT 1559.330 -17.310 1560.510 -16.130 ;
        RECT 1557.730 -18.910 1558.910 -17.730 ;
        RECT 1559.330 -18.910 1560.510 -17.730 ;
        RECT 1737.730 3537.410 1738.910 3538.590 ;
        RECT 1739.330 3537.410 1740.510 3538.590 ;
        RECT 1737.730 3535.810 1738.910 3536.990 ;
        RECT 1739.330 3535.810 1740.510 3536.990 ;
        RECT 1737.730 3364.690 1738.910 3365.870 ;
        RECT 1739.330 3364.690 1740.510 3365.870 ;
        RECT 1737.730 3363.090 1738.910 3364.270 ;
        RECT 1739.330 3363.090 1740.510 3364.270 ;
        RECT 1737.730 3184.690 1738.910 3185.870 ;
        RECT 1739.330 3184.690 1740.510 3185.870 ;
        RECT 1737.730 3183.090 1738.910 3184.270 ;
        RECT 1739.330 3183.090 1740.510 3184.270 ;
        RECT 1737.730 3004.690 1738.910 3005.870 ;
        RECT 1739.330 3004.690 1740.510 3005.870 ;
        RECT 1737.730 3003.090 1738.910 3004.270 ;
        RECT 1739.330 3003.090 1740.510 3004.270 ;
        RECT 1737.730 2824.690 1738.910 2825.870 ;
        RECT 1739.330 2824.690 1740.510 2825.870 ;
        RECT 1737.730 2823.090 1738.910 2824.270 ;
        RECT 1739.330 2823.090 1740.510 2824.270 ;
        RECT 1737.730 2644.690 1738.910 2645.870 ;
        RECT 1739.330 2644.690 1740.510 2645.870 ;
        RECT 1737.730 2643.090 1738.910 2644.270 ;
        RECT 1739.330 2643.090 1740.510 2644.270 ;
        RECT 1737.730 2464.690 1738.910 2465.870 ;
        RECT 1739.330 2464.690 1740.510 2465.870 ;
        RECT 1737.730 2463.090 1738.910 2464.270 ;
        RECT 1739.330 2463.090 1740.510 2464.270 ;
        RECT 1737.730 2284.690 1738.910 2285.870 ;
        RECT 1739.330 2284.690 1740.510 2285.870 ;
        RECT 1737.730 2283.090 1738.910 2284.270 ;
        RECT 1739.330 2283.090 1740.510 2284.270 ;
        RECT 1737.730 2104.690 1738.910 2105.870 ;
        RECT 1739.330 2104.690 1740.510 2105.870 ;
        RECT 1737.730 2103.090 1738.910 2104.270 ;
        RECT 1739.330 2103.090 1740.510 2104.270 ;
        RECT 1737.730 1924.690 1738.910 1925.870 ;
        RECT 1739.330 1924.690 1740.510 1925.870 ;
        RECT 1737.730 1923.090 1738.910 1924.270 ;
        RECT 1739.330 1923.090 1740.510 1924.270 ;
        RECT 1737.730 1744.690 1738.910 1745.870 ;
        RECT 1739.330 1744.690 1740.510 1745.870 ;
        RECT 1737.730 1743.090 1738.910 1744.270 ;
        RECT 1739.330 1743.090 1740.510 1744.270 ;
        RECT 1737.730 1564.690 1738.910 1565.870 ;
        RECT 1739.330 1564.690 1740.510 1565.870 ;
        RECT 1737.730 1563.090 1738.910 1564.270 ;
        RECT 1739.330 1563.090 1740.510 1564.270 ;
        RECT 1737.730 1384.690 1738.910 1385.870 ;
        RECT 1739.330 1384.690 1740.510 1385.870 ;
        RECT 1737.730 1383.090 1738.910 1384.270 ;
        RECT 1739.330 1383.090 1740.510 1384.270 ;
        RECT 1737.730 1204.690 1738.910 1205.870 ;
        RECT 1739.330 1204.690 1740.510 1205.870 ;
        RECT 1737.730 1203.090 1738.910 1204.270 ;
        RECT 1739.330 1203.090 1740.510 1204.270 ;
        RECT 1737.730 1024.690 1738.910 1025.870 ;
        RECT 1739.330 1024.690 1740.510 1025.870 ;
        RECT 1737.730 1023.090 1738.910 1024.270 ;
        RECT 1739.330 1023.090 1740.510 1024.270 ;
        RECT 1737.730 844.690 1738.910 845.870 ;
        RECT 1739.330 844.690 1740.510 845.870 ;
        RECT 1737.730 843.090 1738.910 844.270 ;
        RECT 1739.330 843.090 1740.510 844.270 ;
        RECT 1737.730 664.690 1738.910 665.870 ;
        RECT 1739.330 664.690 1740.510 665.870 ;
        RECT 1737.730 663.090 1738.910 664.270 ;
        RECT 1739.330 663.090 1740.510 664.270 ;
        RECT 1737.730 484.690 1738.910 485.870 ;
        RECT 1739.330 484.690 1740.510 485.870 ;
        RECT 1737.730 483.090 1738.910 484.270 ;
        RECT 1739.330 483.090 1740.510 484.270 ;
        RECT 1737.730 304.690 1738.910 305.870 ;
        RECT 1739.330 304.690 1740.510 305.870 ;
        RECT 1737.730 303.090 1738.910 304.270 ;
        RECT 1739.330 303.090 1740.510 304.270 ;
        RECT 1737.730 124.690 1738.910 125.870 ;
        RECT 1739.330 124.690 1740.510 125.870 ;
        RECT 1737.730 123.090 1738.910 124.270 ;
        RECT 1739.330 123.090 1740.510 124.270 ;
        RECT 1737.730 -17.310 1738.910 -16.130 ;
        RECT 1739.330 -17.310 1740.510 -16.130 ;
        RECT 1737.730 -18.910 1738.910 -17.730 ;
        RECT 1739.330 -18.910 1740.510 -17.730 ;
        RECT 1917.730 3537.410 1918.910 3538.590 ;
        RECT 1919.330 3537.410 1920.510 3538.590 ;
        RECT 1917.730 3535.810 1918.910 3536.990 ;
        RECT 1919.330 3535.810 1920.510 3536.990 ;
        RECT 1917.730 3364.690 1918.910 3365.870 ;
        RECT 1919.330 3364.690 1920.510 3365.870 ;
        RECT 1917.730 3363.090 1918.910 3364.270 ;
        RECT 1919.330 3363.090 1920.510 3364.270 ;
        RECT 1917.730 3184.690 1918.910 3185.870 ;
        RECT 1919.330 3184.690 1920.510 3185.870 ;
        RECT 1917.730 3183.090 1918.910 3184.270 ;
        RECT 1919.330 3183.090 1920.510 3184.270 ;
        RECT 1917.730 3004.690 1918.910 3005.870 ;
        RECT 1919.330 3004.690 1920.510 3005.870 ;
        RECT 1917.730 3003.090 1918.910 3004.270 ;
        RECT 1919.330 3003.090 1920.510 3004.270 ;
        RECT 1917.730 2824.690 1918.910 2825.870 ;
        RECT 1919.330 2824.690 1920.510 2825.870 ;
        RECT 1917.730 2823.090 1918.910 2824.270 ;
        RECT 1919.330 2823.090 1920.510 2824.270 ;
        RECT 1917.730 2644.690 1918.910 2645.870 ;
        RECT 1919.330 2644.690 1920.510 2645.870 ;
        RECT 1917.730 2643.090 1918.910 2644.270 ;
        RECT 1919.330 2643.090 1920.510 2644.270 ;
        RECT 1917.730 2464.690 1918.910 2465.870 ;
        RECT 1919.330 2464.690 1920.510 2465.870 ;
        RECT 1917.730 2463.090 1918.910 2464.270 ;
        RECT 1919.330 2463.090 1920.510 2464.270 ;
        RECT 1917.730 2284.690 1918.910 2285.870 ;
        RECT 1919.330 2284.690 1920.510 2285.870 ;
        RECT 1917.730 2283.090 1918.910 2284.270 ;
        RECT 1919.330 2283.090 1920.510 2284.270 ;
        RECT 1917.730 2104.690 1918.910 2105.870 ;
        RECT 1919.330 2104.690 1920.510 2105.870 ;
        RECT 1917.730 2103.090 1918.910 2104.270 ;
        RECT 1919.330 2103.090 1920.510 2104.270 ;
        RECT 1917.730 1924.690 1918.910 1925.870 ;
        RECT 1919.330 1924.690 1920.510 1925.870 ;
        RECT 1917.730 1923.090 1918.910 1924.270 ;
        RECT 1919.330 1923.090 1920.510 1924.270 ;
        RECT 1917.730 1744.690 1918.910 1745.870 ;
        RECT 1919.330 1744.690 1920.510 1745.870 ;
        RECT 1917.730 1743.090 1918.910 1744.270 ;
        RECT 1919.330 1743.090 1920.510 1744.270 ;
        RECT 1917.730 1564.690 1918.910 1565.870 ;
        RECT 1919.330 1564.690 1920.510 1565.870 ;
        RECT 1917.730 1563.090 1918.910 1564.270 ;
        RECT 1919.330 1563.090 1920.510 1564.270 ;
        RECT 1917.730 1384.690 1918.910 1385.870 ;
        RECT 1919.330 1384.690 1920.510 1385.870 ;
        RECT 1917.730 1383.090 1918.910 1384.270 ;
        RECT 1919.330 1383.090 1920.510 1384.270 ;
        RECT 1917.730 1204.690 1918.910 1205.870 ;
        RECT 1919.330 1204.690 1920.510 1205.870 ;
        RECT 1917.730 1203.090 1918.910 1204.270 ;
        RECT 1919.330 1203.090 1920.510 1204.270 ;
        RECT 1917.730 1024.690 1918.910 1025.870 ;
        RECT 1919.330 1024.690 1920.510 1025.870 ;
        RECT 1917.730 1023.090 1918.910 1024.270 ;
        RECT 1919.330 1023.090 1920.510 1024.270 ;
        RECT 1917.730 844.690 1918.910 845.870 ;
        RECT 1919.330 844.690 1920.510 845.870 ;
        RECT 1917.730 843.090 1918.910 844.270 ;
        RECT 1919.330 843.090 1920.510 844.270 ;
        RECT 1917.730 664.690 1918.910 665.870 ;
        RECT 1919.330 664.690 1920.510 665.870 ;
        RECT 1917.730 663.090 1918.910 664.270 ;
        RECT 1919.330 663.090 1920.510 664.270 ;
        RECT 1917.730 484.690 1918.910 485.870 ;
        RECT 1919.330 484.690 1920.510 485.870 ;
        RECT 1917.730 483.090 1918.910 484.270 ;
        RECT 1919.330 483.090 1920.510 484.270 ;
        RECT 1917.730 304.690 1918.910 305.870 ;
        RECT 1919.330 304.690 1920.510 305.870 ;
        RECT 1917.730 303.090 1918.910 304.270 ;
        RECT 1919.330 303.090 1920.510 304.270 ;
        RECT 1917.730 124.690 1918.910 125.870 ;
        RECT 1919.330 124.690 1920.510 125.870 ;
        RECT 1917.730 123.090 1918.910 124.270 ;
        RECT 1919.330 123.090 1920.510 124.270 ;
        RECT 1917.730 -17.310 1918.910 -16.130 ;
        RECT 1919.330 -17.310 1920.510 -16.130 ;
        RECT 1917.730 -18.910 1918.910 -17.730 ;
        RECT 1919.330 -18.910 1920.510 -17.730 ;
        RECT 2097.730 3537.410 2098.910 3538.590 ;
        RECT 2099.330 3537.410 2100.510 3538.590 ;
        RECT 2097.730 3535.810 2098.910 3536.990 ;
        RECT 2099.330 3535.810 2100.510 3536.990 ;
        RECT 2097.730 3364.690 2098.910 3365.870 ;
        RECT 2099.330 3364.690 2100.510 3365.870 ;
        RECT 2097.730 3363.090 2098.910 3364.270 ;
        RECT 2099.330 3363.090 2100.510 3364.270 ;
        RECT 2097.730 3184.690 2098.910 3185.870 ;
        RECT 2099.330 3184.690 2100.510 3185.870 ;
        RECT 2097.730 3183.090 2098.910 3184.270 ;
        RECT 2099.330 3183.090 2100.510 3184.270 ;
        RECT 2097.730 3004.690 2098.910 3005.870 ;
        RECT 2099.330 3004.690 2100.510 3005.870 ;
        RECT 2097.730 3003.090 2098.910 3004.270 ;
        RECT 2099.330 3003.090 2100.510 3004.270 ;
        RECT 2097.730 2824.690 2098.910 2825.870 ;
        RECT 2099.330 2824.690 2100.510 2825.870 ;
        RECT 2097.730 2823.090 2098.910 2824.270 ;
        RECT 2099.330 2823.090 2100.510 2824.270 ;
        RECT 2097.730 2644.690 2098.910 2645.870 ;
        RECT 2099.330 2644.690 2100.510 2645.870 ;
        RECT 2097.730 2643.090 2098.910 2644.270 ;
        RECT 2099.330 2643.090 2100.510 2644.270 ;
        RECT 2097.730 2464.690 2098.910 2465.870 ;
        RECT 2099.330 2464.690 2100.510 2465.870 ;
        RECT 2097.730 2463.090 2098.910 2464.270 ;
        RECT 2099.330 2463.090 2100.510 2464.270 ;
        RECT 2097.730 2284.690 2098.910 2285.870 ;
        RECT 2099.330 2284.690 2100.510 2285.870 ;
        RECT 2097.730 2283.090 2098.910 2284.270 ;
        RECT 2099.330 2283.090 2100.510 2284.270 ;
        RECT 2097.730 2104.690 2098.910 2105.870 ;
        RECT 2099.330 2104.690 2100.510 2105.870 ;
        RECT 2097.730 2103.090 2098.910 2104.270 ;
        RECT 2099.330 2103.090 2100.510 2104.270 ;
        RECT 2097.730 1924.690 2098.910 1925.870 ;
        RECT 2099.330 1924.690 2100.510 1925.870 ;
        RECT 2097.730 1923.090 2098.910 1924.270 ;
        RECT 2099.330 1923.090 2100.510 1924.270 ;
        RECT 2097.730 1744.690 2098.910 1745.870 ;
        RECT 2099.330 1744.690 2100.510 1745.870 ;
        RECT 2097.730 1743.090 2098.910 1744.270 ;
        RECT 2099.330 1743.090 2100.510 1744.270 ;
        RECT 2097.730 1564.690 2098.910 1565.870 ;
        RECT 2099.330 1564.690 2100.510 1565.870 ;
        RECT 2097.730 1563.090 2098.910 1564.270 ;
        RECT 2099.330 1563.090 2100.510 1564.270 ;
        RECT 2097.730 1384.690 2098.910 1385.870 ;
        RECT 2099.330 1384.690 2100.510 1385.870 ;
        RECT 2097.730 1383.090 2098.910 1384.270 ;
        RECT 2099.330 1383.090 2100.510 1384.270 ;
        RECT 2097.730 1204.690 2098.910 1205.870 ;
        RECT 2099.330 1204.690 2100.510 1205.870 ;
        RECT 2097.730 1203.090 2098.910 1204.270 ;
        RECT 2099.330 1203.090 2100.510 1204.270 ;
        RECT 2097.730 1024.690 2098.910 1025.870 ;
        RECT 2099.330 1024.690 2100.510 1025.870 ;
        RECT 2097.730 1023.090 2098.910 1024.270 ;
        RECT 2099.330 1023.090 2100.510 1024.270 ;
        RECT 2097.730 844.690 2098.910 845.870 ;
        RECT 2099.330 844.690 2100.510 845.870 ;
        RECT 2097.730 843.090 2098.910 844.270 ;
        RECT 2099.330 843.090 2100.510 844.270 ;
        RECT 2097.730 664.690 2098.910 665.870 ;
        RECT 2099.330 664.690 2100.510 665.870 ;
        RECT 2097.730 663.090 2098.910 664.270 ;
        RECT 2099.330 663.090 2100.510 664.270 ;
        RECT 2097.730 484.690 2098.910 485.870 ;
        RECT 2099.330 484.690 2100.510 485.870 ;
        RECT 2097.730 483.090 2098.910 484.270 ;
        RECT 2099.330 483.090 2100.510 484.270 ;
        RECT 2097.730 304.690 2098.910 305.870 ;
        RECT 2099.330 304.690 2100.510 305.870 ;
        RECT 2097.730 303.090 2098.910 304.270 ;
        RECT 2099.330 303.090 2100.510 304.270 ;
        RECT 2097.730 124.690 2098.910 125.870 ;
        RECT 2099.330 124.690 2100.510 125.870 ;
        RECT 2097.730 123.090 2098.910 124.270 ;
        RECT 2099.330 123.090 2100.510 124.270 ;
        RECT 2097.730 -17.310 2098.910 -16.130 ;
        RECT 2099.330 -17.310 2100.510 -16.130 ;
        RECT 2097.730 -18.910 2098.910 -17.730 ;
        RECT 2099.330 -18.910 2100.510 -17.730 ;
        RECT 2277.730 3537.410 2278.910 3538.590 ;
        RECT 2279.330 3537.410 2280.510 3538.590 ;
        RECT 2277.730 3535.810 2278.910 3536.990 ;
        RECT 2279.330 3535.810 2280.510 3536.990 ;
        RECT 2277.730 3364.690 2278.910 3365.870 ;
        RECT 2279.330 3364.690 2280.510 3365.870 ;
        RECT 2277.730 3363.090 2278.910 3364.270 ;
        RECT 2279.330 3363.090 2280.510 3364.270 ;
        RECT 2277.730 3184.690 2278.910 3185.870 ;
        RECT 2279.330 3184.690 2280.510 3185.870 ;
        RECT 2277.730 3183.090 2278.910 3184.270 ;
        RECT 2279.330 3183.090 2280.510 3184.270 ;
        RECT 2277.730 3004.690 2278.910 3005.870 ;
        RECT 2279.330 3004.690 2280.510 3005.870 ;
        RECT 2277.730 3003.090 2278.910 3004.270 ;
        RECT 2279.330 3003.090 2280.510 3004.270 ;
        RECT 2277.730 2824.690 2278.910 2825.870 ;
        RECT 2279.330 2824.690 2280.510 2825.870 ;
        RECT 2277.730 2823.090 2278.910 2824.270 ;
        RECT 2279.330 2823.090 2280.510 2824.270 ;
        RECT 2277.730 2644.690 2278.910 2645.870 ;
        RECT 2279.330 2644.690 2280.510 2645.870 ;
        RECT 2277.730 2643.090 2278.910 2644.270 ;
        RECT 2279.330 2643.090 2280.510 2644.270 ;
        RECT 2277.730 2464.690 2278.910 2465.870 ;
        RECT 2279.330 2464.690 2280.510 2465.870 ;
        RECT 2277.730 2463.090 2278.910 2464.270 ;
        RECT 2279.330 2463.090 2280.510 2464.270 ;
        RECT 2277.730 2284.690 2278.910 2285.870 ;
        RECT 2279.330 2284.690 2280.510 2285.870 ;
        RECT 2277.730 2283.090 2278.910 2284.270 ;
        RECT 2279.330 2283.090 2280.510 2284.270 ;
        RECT 2277.730 2104.690 2278.910 2105.870 ;
        RECT 2279.330 2104.690 2280.510 2105.870 ;
        RECT 2277.730 2103.090 2278.910 2104.270 ;
        RECT 2279.330 2103.090 2280.510 2104.270 ;
        RECT 2277.730 1924.690 2278.910 1925.870 ;
        RECT 2279.330 1924.690 2280.510 1925.870 ;
        RECT 2277.730 1923.090 2278.910 1924.270 ;
        RECT 2279.330 1923.090 2280.510 1924.270 ;
        RECT 2277.730 1744.690 2278.910 1745.870 ;
        RECT 2279.330 1744.690 2280.510 1745.870 ;
        RECT 2277.730 1743.090 2278.910 1744.270 ;
        RECT 2279.330 1743.090 2280.510 1744.270 ;
        RECT 2277.730 1564.690 2278.910 1565.870 ;
        RECT 2279.330 1564.690 2280.510 1565.870 ;
        RECT 2277.730 1563.090 2278.910 1564.270 ;
        RECT 2279.330 1563.090 2280.510 1564.270 ;
        RECT 2277.730 1384.690 2278.910 1385.870 ;
        RECT 2279.330 1384.690 2280.510 1385.870 ;
        RECT 2277.730 1383.090 2278.910 1384.270 ;
        RECT 2279.330 1383.090 2280.510 1384.270 ;
        RECT 2277.730 1204.690 2278.910 1205.870 ;
        RECT 2279.330 1204.690 2280.510 1205.870 ;
        RECT 2277.730 1203.090 2278.910 1204.270 ;
        RECT 2279.330 1203.090 2280.510 1204.270 ;
        RECT 2277.730 1024.690 2278.910 1025.870 ;
        RECT 2279.330 1024.690 2280.510 1025.870 ;
        RECT 2277.730 1023.090 2278.910 1024.270 ;
        RECT 2279.330 1023.090 2280.510 1024.270 ;
        RECT 2277.730 844.690 2278.910 845.870 ;
        RECT 2279.330 844.690 2280.510 845.870 ;
        RECT 2277.730 843.090 2278.910 844.270 ;
        RECT 2279.330 843.090 2280.510 844.270 ;
        RECT 2277.730 664.690 2278.910 665.870 ;
        RECT 2279.330 664.690 2280.510 665.870 ;
        RECT 2277.730 663.090 2278.910 664.270 ;
        RECT 2279.330 663.090 2280.510 664.270 ;
        RECT 2277.730 484.690 2278.910 485.870 ;
        RECT 2279.330 484.690 2280.510 485.870 ;
        RECT 2277.730 483.090 2278.910 484.270 ;
        RECT 2279.330 483.090 2280.510 484.270 ;
        RECT 2277.730 304.690 2278.910 305.870 ;
        RECT 2279.330 304.690 2280.510 305.870 ;
        RECT 2277.730 303.090 2278.910 304.270 ;
        RECT 2279.330 303.090 2280.510 304.270 ;
        RECT 2277.730 124.690 2278.910 125.870 ;
        RECT 2279.330 124.690 2280.510 125.870 ;
        RECT 2277.730 123.090 2278.910 124.270 ;
        RECT 2279.330 123.090 2280.510 124.270 ;
        RECT 2277.730 -17.310 2278.910 -16.130 ;
        RECT 2279.330 -17.310 2280.510 -16.130 ;
        RECT 2277.730 -18.910 2278.910 -17.730 ;
        RECT 2279.330 -18.910 2280.510 -17.730 ;
        RECT 2457.730 3537.410 2458.910 3538.590 ;
        RECT 2459.330 3537.410 2460.510 3538.590 ;
        RECT 2457.730 3535.810 2458.910 3536.990 ;
        RECT 2459.330 3535.810 2460.510 3536.990 ;
        RECT 2457.730 3364.690 2458.910 3365.870 ;
        RECT 2459.330 3364.690 2460.510 3365.870 ;
        RECT 2457.730 3363.090 2458.910 3364.270 ;
        RECT 2459.330 3363.090 2460.510 3364.270 ;
        RECT 2457.730 3184.690 2458.910 3185.870 ;
        RECT 2459.330 3184.690 2460.510 3185.870 ;
        RECT 2457.730 3183.090 2458.910 3184.270 ;
        RECT 2459.330 3183.090 2460.510 3184.270 ;
        RECT 2457.730 3004.690 2458.910 3005.870 ;
        RECT 2459.330 3004.690 2460.510 3005.870 ;
        RECT 2457.730 3003.090 2458.910 3004.270 ;
        RECT 2459.330 3003.090 2460.510 3004.270 ;
        RECT 2457.730 2824.690 2458.910 2825.870 ;
        RECT 2459.330 2824.690 2460.510 2825.870 ;
        RECT 2457.730 2823.090 2458.910 2824.270 ;
        RECT 2459.330 2823.090 2460.510 2824.270 ;
        RECT 2457.730 2644.690 2458.910 2645.870 ;
        RECT 2459.330 2644.690 2460.510 2645.870 ;
        RECT 2457.730 2643.090 2458.910 2644.270 ;
        RECT 2459.330 2643.090 2460.510 2644.270 ;
        RECT 2457.730 2464.690 2458.910 2465.870 ;
        RECT 2459.330 2464.690 2460.510 2465.870 ;
        RECT 2457.730 2463.090 2458.910 2464.270 ;
        RECT 2459.330 2463.090 2460.510 2464.270 ;
        RECT 2457.730 2284.690 2458.910 2285.870 ;
        RECT 2459.330 2284.690 2460.510 2285.870 ;
        RECT 2457.730 2283.090 2458.910 2284.270 ;
        RECT 2459.330 2283.090 2460.510 2284.270 ;
        RECT 2457.730 2104.690 2458.910 2105.870 ;
        RECT 2459.330 2104.690 2460.510 2105.870 ;
        RECT 2457.730 2103.090 2458.910 2104.270 ;
        RECT 2459.330 2103.090 2460.510 2104.270 ;
        RECT 2457.730 1924.690 2458.910 1925.870 ;
        RECT 2459.330 1924.690 2460.510 1925.870 ;
        RECT 2457.730 1923.090 2458.910 1924.270 ;
        RECT 2459.330 1923.090 2460.510 1924.270 ;
        RECT 2457.730 1744.690 2458.910 1745.870 ;
        RECT 2459.330 1744.690 2460.510 1745.870 ;
        RECT 2457.730 1743.090 2458.910 1744.270 ;
        RECT 2459.330 1743.090 2460.510 1744.270 ;
        RECT 2457.730 1564.690 2458.910 1565.870 ;
        RECT 2459.330 1564.690 2460.510 1565.870 ;
        RECT 2457.730 1563.090 2458.910 1564.270 ;
        RECT 2459.330 1563.090 2460.510 1564.270 ;
        RECT 2457.730 1384.690 2458.910 1385.870 ;
        RECT 2459.330 1384.690 2460.510 1385.870 ;
        RECT 2457.730 1383.090 2458.910 1384.270 ;
        RECT 2459.330 1383.090 2460.510 1384.270 ;
        RECT 2457.730 1204.690 2458.910 1205.870 ;
        RECT 2459.330 1204.690 2460.510 1205.870 ;
        RECT 2457.730 1203.090 2458.910 1204.270 ;
        RECT 2459.330 1203.090 2460.510 1204.270 ;
        RECT 2457.730 1024.690 2458.910 1025.870 ;
        RECT 2459.330 1024.690 2460.510 1025.870 ;
        RECT 2457.730 1023.090 2458.910 1024.270 ;
        RECT 2459.330 1023.090 2460.510 1024.270 ;
        RECT 2457.730 844.690 2458.910 845.870 ;
        RECT 2459.330 844.690 2460.510 845.870 ;
        RECT 2457.730 843.090 2458.910 844.270 ;
        RECT 2459.330 843.090 2460.510 844.270 ;
        RECT 2457.730 664.690 2458.910 665.870 ;
        RECT 2459.330 664.690 2460.510 665.870 ;
        RECT 2457.730 663.090 2458.910 664.270 ;
        RECT 2459.330 663.090 2460.510 664.270 ;
        RECT 2457.730 484.690 2458.910 485.870 ;
        RECT 2459.330 484.690 2460.510 485.870 ;
        RECT 2457.730 483.090 2458.910 484.270 ;
        RECT 2459.330 483.090 2460.510 484.270 ;
        RECT 2457.730 304.690 2458.910 305.870 ;
        RECT 2459.330 304.690 2460.510 305.870 ;
        RECT 2457.730 303.090 2458.910 304.270 ;
        RECT 2459.330 303.090 2460.510 304.270 ;
        RECT 2457.730 124.690 2458.910 125.870 ;
        RECT 2459.330 124.690 2460.510 125.870 ;
        RECT 2457.730 123.090 2458.910 124.270 ;
        RECT 2459.330 123.090 2460.510 124.270 ;
        RECT 2457.730 -17.310 2458.910 -16.130 ;
        RECT 2459.330 -17.310 2460.510 -16.130 ;
        RECT 2457.730 -18.910 2458.910 -17.730 ;
        RECT 2459.330 -18.910 2460.510 -17.730 ;
        RECT 2637.730 3537.410 2638.910 3538.590 ;
        RECT 2639.330 3537.410 2640.510 3538.590 ;
        RECT 2637.730 3535.810 2638.910 3536.990 ;
        RECT 2639.330 3535.810 2640.510 3536.990 ;
        RECT 2637.730 3364.690 2638.910 3365.870 ;
        RECT 2639.330 3364.690 2640.510 3365.870 ;
        RECT 2637.730 3363.090 2638.910 3364.270 ;
        RECT 2639.330 3363.090 2640.510 3364.270 ;
        RECT 2637.730 3184.690 2638.910 3185.870 ;
        RECT 2639.330 3184.690 2640.510 3185.870 ;
        RECT 2637.730 3183.090 2638.910 3184.270 ;
        RECT 2639.330 3183.090 2640.510 3184.270 ;
        RECT 2637.730 3004.690 2638.910 3005.870 ;
        RECT 2639.330 3004.690 2640.510 3005.870 ;
        RECT 2637.730 3003.090 2638.910 3004.270 ;
        RECT 2639.330 3003.090 2640.510 3004.270 ;
        RECT 2637.730 2824.690 2638.910 2825.870 ;
        RECT 2639.330 2824.690 2640.510 2825.870 ;
        RECT 2637.730 2823.090 2638.910 2824.270 ;
        RECT 2639.330 2823.090 2640.510 2824.270 ;
        RECT 2637.730 2644.690 2638.910 2645.870 ;
        RECT 2639.330 2644.690 2640.510 2645.870 ;
        RECT 2637.730 2643.090 2638.910 2644.270 ;
        RECT 2639.330 2643.090 2640.510 2644.270 ;
        RECT 2637.730 2464.690 2638.910 2465.870 ;
        RECT 2639.330 2464.690 2640.510 2465.870 ;
        RECT 2637.730 2463.090 2638.910 2464.270 ;
        RECT 2639.330 2463.090 2640.510 2464.270 ;
        RECT 2637.730 2284.690 2638.910 2285.870 ;
        RECT 2639.330 2284.690 2640.510 2285.870 ;
        RECT 2637.730 2283.090 2638.910 2284.270 ;
        RECT 2639.330 2283.090 2640.510 2284.270 ;
        RECT 2637.730 2104.690 2638.910 2105.870 ;
        RECT 2639.330 2104.690 2640.510 2105.870 ;
        RECT 2637.730 2103.090 2638.910 2104.270 ;
        RECT 2639.330 2103.090 2640.510 2104.270 ;
        RECT 2637.730 1924.690 2638.910 1925.870 ;
        RECT 2639.330 1924.690 2640.510 1925.870 ;
        RECT 2637.730 1923.090 2638.910 1924.270 ;
        RECT 2639.330 1923.090 2640.510 1924.270 ;
        RECT 2637.730 1744.690 2638.910 1745.870 ;
        RECT 2639.330 1744.690 2640.510 1745.870 ;
        RECT 2637.730 1743.090 2638.910 1744.270 ;
        RECT 2639.330 1743.090 2640.510 1744.270 ;
        RECT 2637.730 1564.690 2638.910 1565.870 ;
        RECT 2639.330 1564.690 2640.510 1565.870 ;
        RECT 2637.730 1563.090 2638.910 1564.270 ;
        RECT 2639.330 1563.090 2640.510 1564.270 ;
        RECT 2637.730 1384.690 2638.910 1385.870 ;
        RECT 2639.330 1384.690 2640.510 1385.870 ;
        RECT 2637.730 1383.090 2638.910 1384.270 ;
        RECT 2639.330 1383.090 2640.510 1384.270 ;
        RECT 2637.730 1204.690 2638.910 1205.870 ;
        RECT 2639.330 1204.690 2640.510 1205.870 ;
        RECT 2637.730 1203.090 2638.910 1204.270 ;
        RECT 2639.330 1203.090 2640.510 1204.270 ;
        RECT 2637.730 1024.690 2638.910 1025.870 ;
        RECT 2639.330 1024.690 2640.510 1025.870 ;
        RECT 2637.730 1023.090 2638.910 1024.270 ;
        RECT 2639.330 1023.090 2640.510 1024.270 ;
        RECT 2637.730 844.690 2638.910 845.870 ;
        RECT 2639.330 844.690 2640.510 845.870 ;
        RECT 2637.730 843.090 2638.910 844.270 ;
        RECT 2639.330 843.090 2640.510 844.270 ;
        RECT 2637.730 664.690 2638.910 665.870 ;
        RECT 2639.330 664.690 2640.510 665.870 ;
        RECT 2637.730 663.090 2638.910 664.270 ;
        RECT 2639.330 663.090 2640.510 664.270 ;
        RECT 2637.730 484.690 2638.910 485.870 ;
        RECT 2639.330 484.690 2640.510 485.870 ;
        RECT 2637.730 483.090 2638.910 484.270 ;
        RECT 2639.330 483.090 2640.510 484.270 ;
        RECT 2637.730 304.690 2638.910 305.870 ;
        RECT 2639.330 304.690 2640.510 305.870 ;
        RECT 2637.730 303.090 2638.910 304.270 ;
        RECT 2639.330 303.090 2640.510 304.270 ;
        RECT 2637.730 124.690 2638.910 125.870 ;
        RECT 2639.330 124.690 2640.510 125.870 ;
        RECT 2637.730 123.090 2638.910 124.270 ;
        RECT 2639.330 123.090 2640.510 124.270 ;
        RECT 2637.730 -17.310 2638.910 -16.130 ;
        RECT 2639.330 -17.310 2640.510 -16.130 ;
        RECT 2637.730 -18.910 2638.910 -17.730 ;
        RECT 2639.330 -18.910 2640.510 -17.730 ;
        RECT 2817.730 3537.410 2818.910 3538.590 ;
        RECT 2819.330 3537.410 2820.510 3538.590 ;
        RECT 2817.730 3535.810 2818.910 3536.990 ;
        RECT 2819.330 3535.810 2820.510 3536.990 ;
        RECT 2817.730 3364.690 2818.910 3365.870 ;
        RECT 2819.330 3364.690 2820.510 3365.870 ;
        RECT 2817.730 3363.090 2818.910 3364.270 ;
        RECT 2819.330 3363.090 2820.510 3364.270 ;
        RECT 2817.730 3184.690 2818.910 3185.870 ;
        RECT 2819.330 3184.690 2820.510 3185.870 ;
        RECT 2817.730 3183.090 2818.910 3184.270 ;
        RECT 2819.330 3183.090 2820.510 3184.270 ;
        RECT 2817.730 3004.690 2818.910 3005.870 ;
        RECT 2819.330 3004.690 2820.510 3005.870 ;
        RECT 2817.730 3003.090 2818.910 3004.270 ;
        RECT 2819.330 3003.090 2820.510 3004.270 ;
        RECT 2817.730 2824.690 2818.910 2825.870 ;
        RECT 2819.330 2824.690 2820.510 2825.870 ;
        RECT 2817.730 2823.090 2818.910 2824.270 ;
        RECT 2819.330 2823.090 2820.510 2824.270 ;
        RECT 2817.730 2644.690 2818.910 2645.870 ;
        RECT 2819.330 2644.690 2820.510 2645.870 ;
        RECT 2817.730 2643.090 2818.910 2644.270 ;
        RECT 2819.330 2643.090 2820.510 2644.270 ;
        RECT 2817.730 2464.690 2818.910 2465.870 ;
        RECT 2819.330 2464.690 2820.510 2465.870 ;
        RECT 2817.730 2463.090 2818.910 2464.270 ;
        RECT 2819.330 2463.090 2820.510 2464.270 ;
        RECT 2817.730 2284.690 2818.910 2285.870 ;
        RECT 2819.330 2284.690 2820.510 2285.870 ;
        RECT 2817.730 2283.090 2818.910 2284.270 ;
        RECT 2819.330 2283.090 2820.510 2284.270 ;
        RECT 2817.730 2104.690 2818.910 2105.870 ;
        RECT 2819.330 2104.690 2820.510 2105.870 ;
        RECT 2817.730 2103.090 2818.910 2104.270 ;
        RECT 2819.330 2103.090 2820.510 2104.270 ;
        RECT 2817.730 1924.690 2818.910 1925.870 ;
        RECT 2819.330 1924.690 2820.510 1925.870 ;
        RECT 2817.730 1923.090 2818.910 1924.270 ;
        RECT 2819.330 1923.090 2820.510 1924.270 ;
        RECT 2817.730 1744.690 2818.910 1745.870 ;
        RECT 2819.330 1744.690 2820.510 1745.870 ;
        RECT 2817.730 1743.090 2818.910 1744.270 ;
        RECT 2819.330 1743.090 2820.510 1744.270 ;
        RECT 2817.730 1564.690 2818.910 1565.870 ;
        RECT 2819.330 1564.690 2820.510 1565.870 ;
        RECT 2817.730 1563.090 2818.910 1564.270 ;
        RECT 2819.330 1563.090 2820.510 1564.270 ;
        RECT 2817.730 1384.690 2818.910 1385.870 ;
        RECT 2819.330 1384.690 2820.510 1385.870 ;
        RECT 2817.730 1383.090 2818.910 1384.270 ;
        RECT 2819.330 1383.090 2820.510 1384.270 ;
        RECT 2817.730 1204.690 2818.910 1205.870 ;
        RECT 2819.330 1204.690 2820.510 1205.870 ;
        RECT 2817.730 1203.090 2818.910 1204.270 ;
        RECT 2819.330 1203.090 2820.510 1204.270 ;
        RECT 2817.730 1024.690 2818.910 1025.870 ;
        RECT 2819.330 1024.690 2820.510 1025.870 ;
        RECT 2817.730 1023.090 2818.910 1024.270 ;
        RECT 2819.330 1023.090 2820.510 1024.270 ;
        RECT 2817.730 844.690 2818.910 845.870 ;
        RECT 2819.330 844.690 2820.510 845.870 ;
        RECT 2817.730 843.090 2818.910 844.270 ;
        RECT 2819.330 843.090 2820.510 844.270 ;
        RECT 2817.730 664.690 2818.910 665.870 ;
        RECT 2819.330 664.690 2820.510 665.870 ;
        RECT 2817.730 663.090 2818.910 664.270 ;
        RECT 2819.330 663.090 2820.510 664.270 ;
        RECT 2817.730 484.690 2818.910 485.870 ;
        RECT 2819.330 484.690 2820.510 485.870 ;
        RECT 2817.730 483.090 2818.910 484.270 ;
        RECT 2819.330 483.090 2820.510 484.270 ;
        RECT 2817.730 304.690 2818.910 305.870 ;
        RECT 2819.330 304.690 2820.510 305.870 ;
        RECT 2817.730 303.090 2818.910 304.270 ;
        RECT 2819.330 303.090 2820.510 304.270 ;
        RECT 2817.730 124.690 2818.910 125.870 ;
        RECT 2819.330 124.690 2820.510 125.870 ;
        RECT 2817.730 123.090 2818.910 124.270 ;
        RECT 2819.330 123.090 2820.510 124.270 ;
        RECT 2817.730 -17.310 2818.910 -16.130 ;
        RECT 2819.330 -17.310 2820.510 -16.130 ;
        RECT 2817.730 -18.910 2818.910 -17.730 ;
        RECT 2819.330 -18.910 2820.510 -17.730 ;
        RECT 2941.110 3537.410 2942.290 3538.590 ;
        RECT 2942.710 3537.410 2943.890 3538.590 ;
        RECT 2941.110 3535.810 2942.290 3536.990 ;
        RECT 2942.710 3535.810 2943.890 3536.990 ;
        RECT 2941.110 3364.690 2942.290 3365.870 ;
        RECT 2942.710 3364.690 2943.890 3365.870 ;
        RECT 2941.110 3363.090 2942.290 3364.270 ;
        RECT 2942.710 3363.090 2943.890 3364.270 ;
        RECT 2941.110 3184.690 2942.290 3185.870 ;
        RECT 2942.710 3184.690 2943.890 3185.870 ;
        RECT 2941.110 3183.090 2942.290 3184.270 ;
        RECT 2942.710 3183.090 2943.890 3184.270 ;
        RECT 2941.110 3004.690 2942.290 3005.870 ;
        RECT 2942.710 3004.690 2943.890 3005.870 ;
        RECT 2941.110 3003.090 2942.290 3004.270 ;
        RECT 2942.710 3003.090 2943.890 3004.270 ;
        RECT 2941.110 2824.690 2942.290 2825.870 ;
        RECT 2942.710 2824.690 2943.890 2825.870 ;
        RECT 2941.110 2823.090 2942.290 2824.270 ;
        RECT 2942.710 2823.090 2943.890 2824.270 ;
        RECT 2941.110 2644.690 2942.290 2645.870 ;
        RECT 2942.710 2644.690 2943.890 2645.870 ;
        RECT 2941.110 2643.090 2942.290 2644.270 ;
        RECT 2942.710 2643.090 2943.890 2644.270 ;
        RECT 2941.110 2464.690 2942.290 2465.870 ;
        RECT 2942.710 2464.690 2943.890 2465.870 ;
        RECT 2941.110 2463.090 2942.290 2464.270 ;
        RECT 2942.710 2463.090 2943.890 2464.270 ;
        RECT 2941.110 2284.690 2942.290 2285.870 ;
        RECT 2942.710 2284.690 2943.890 2285.870 ;
        RECT 2941.110 2283.090 2942.290 2284.270 ;
        RECT 2942.710 2283.090 2943.890 2284.270 ;
        RECT 2941.110 2104.690 2942.290 2105.870 ;
        RECT 2942.710 2104.690 2943.890 2105.870 ;
        RECT 2941.110 2103.090 2942.290 2104.270 ;
        RECT 2942.710 2103.090 2943.890 2104.270 ;
        RECT 2941.110 1924.690 2942.290 1925.870 ;
        RECT 2942.710 1924.690 2943.890 1925.870 ;
        RECT 2941.110 1923.090 2942.290 1924.270 ;
        RECT 2942.710 1923.090 2943.890 1924.270 ;
        RECT 2941.110 1744.690 2942.290 1745.870 ;
        RECT 2942.710 1744.690 2943.890 1745.870 ;
        RECT 2941.110 1743.090 2942.290 1744.270 ;
        RECT 2942.710 1743.090 2943.890 1744.270 ;
        RECT 2941.110 1564.690 2942.290 1565.870 ;
        RECT 2942.710 1564.690 2943.890 1565.870 ;
        RECT 2941.110 1563.090 2942.290 1564.270 ;
        RECT 2942.710 1563.090 2943.890 1564.270 ;
        RECT 2941.110 1384.690 2942.290 1385.870 ;
        RECT 2942.710 1384.690 2943.890 1385.870 ;
        RECT 2941.110 1383.090 2942.290 1384.270 ;
        RECT 2942.710 1383.090 2943.890 1384.270 ;
        RECT 2941.110 1204.690 2942.290 1205.870 ;
        RECT 2942.710 1204.690 2943.890 1205.870 ;
        RECT 2941.110 1203.090 2942.290 1204.270 ;
        RECT 2942.710 1203.090 2943.890 1204.270 ;
        RECT 2941.110 1024.690 2942.290 1025.870 ;
        RECT 2942.710 1024.690 2943.890 1025.870 ;
        RECT 2941.110 1023.090 2942.290 1024.270 ;
        RECT 2942.710 1023.090 2943.890 1024.270 ;
        RECT 2941.110 844.690 2942.290 845.870 ;
        RECT 2942.710 844.690 2943.890 845.870 ;
        RECT 2941.110 843.090 2942.290 844.270 ;
        RECT 2942.710 843.090 2943.890 844.270 ;
        RECT 2941.110 664.690 2942.290 665.870 ;
        RECT 2942.710 664.690 2943.890 665.870 ;
        RECT 2941.110 663.090 2942.290 664.270 ;
        RECT 2942.710 663.090 2943.890 664.270 ;
        RECT 2941.110 484.690 2942.290 485.870 ;
        RECT 2942.710 484.690 2943.890 485.870 ;
        RECT 2941.110 483.090 2942.290 484.270 ;
        RECT 2942.710 483.090 2943.890 484.270 ;
        RECT 2941.110 304.690 2942.290 305.870 ;
        RECT 2942.710 304.690 2943.890 305.870 ;
        RECT 2941.110 303.090 2942.290 304.270 ;
        RECT 2942.710 303.090 2943.890 304.270 ;
        RECT 2941.110 124.690 2942.290 125.870 ;
        RECT 2942.710 124.690 2943.890 125.870 ;
        RECT 2941.110 123.090 2942.290 124.270 ;
        RECT 2942.710 123.090 2943.890 124.270 ;
        RECT 2941.110 -17.310 2942.290 -16.130 ;
        RECT 2942.710 -17.310 2943.890 -16.130 ;
        RECT 2941.110 -18.910 2942.290 -17.730 ;
        RECT 2942.710 -18.910 2943.890 -17.730 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
        RECT -24.430 842.930 2944.050 846.030 ;
        RECT -24.430 662.930 2944.050 666.030 ;
        RECT -24.430 482.930 2944.050 486.030 ;
        RECT -24.430 302.930 2944.050 306.030 ;
        RECT -24.430 122.930 2944.050 126.030 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.930 400.250 202.210 404.000 ;
        RECT 201.640 400.110 202.210 400.250 ;
        RECT 201.640 16.845 201.780 400.110 ;
        RECT 201.930 400.000 202.210 400.110 ;
        RECT 8.370 16.475 8.650 16.845 ;
        RECT 201.570 16.475 201.850 16.845 ;
        RECT 8.440 2.400 8.580 16.475 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 8.370 16.520 8.650 16.800 ;
        RECT 201.570 16.520 201.850 16.800 ;
      LAYER met3 ;
        RECT 8.345 16.810 8.675 16.825 ;
        RECT 201.545 16.810 201.875 16.825 ;
        RECT 8.345 16.510 201.875 16.810 ;
        RECT 8.345 16.495 8.675 16.510 ;
        RECT 201.545 16.495 201.875 16.510 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 201.090 376.280 201.410 376.340 ;
        RECT 202.470 376.280 202.790 376.340 ;
        RECT 201.090 376.140 202.790 376.280 ;
        RECT 201.090 376.080 201.410 376.140 ;
        RECT 202.470 376.080 202.790 376.140 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 201.090 17.580 201.410 17.640 ;
        RECT 14.330 17.440 201.410 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 201.090 17.380 201.410 17.440 ;
      LAYER via ;
        RECT 201.120 376.080 201.380 376.340 ;
        RECT 202.500 376.080 202.760 376.340 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 201.120 17.380 201.380 17.640 ;
      LAYER met2 ;
        RECT 203.770 400.250 204.050 404.000 ;
        RECT 202.560 400.110 204.050 400.250 ;
        RECT 202.560 376.370 202.700 400.110 ;
        RECT 203.770 400.000 204.050 400.110 ;
        RECT 201.120 376.050 201.380 376.370 ;
        RECT 202.500 376.050 202.760 376.370 ;
        RECT 201.180 17.670 201.320 376.050 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 201.120 17.350 201.380 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 207.530 386.480 207.850 386.540 ;
        RECT 209.830 386.480 210.150 386.540 ;
        RECT 207.530 386.340 210.150 386.480 ;
        RECT 207.530 386.280 207.850 386.340 ;
        RECT 209.830 386.280 210.150 386.340 ;
        RECT 38.250 18.260 38.570 18.320 ;
        RECT 207.530 18.260 207.850 18.320 ;
        RECT 38.250 18.120 207.850 18.260 ;
        RECT 38.250 18.060 38.570 18.120 ;
        RECT 207.530 18.060 207.850 18.120 ;
      LAYER via ;
        RECT 207.560 386.280 207.820 386.540 ;
        RECT 209.860 386.280 210.120 386.540 ;
        RECT 38.280 18.060 38.540 18.320 ;
        RECT 207.560 18.060 207.820 18.320 ;
      LAYER met2 ;
        RECT 211.130 400.250 211.410 404.000 ;
        RECT 209.920 400.110 211.410 400.250 ;
        RECT 209.920 386.570 210.060 400.110 ;
        RECT 211.130 400.000 211.410 400.110 ;
        RECT 207.560 386.250 207.820 386.570 ;
        RECT 209.860 386.250 210.120 386.570 ;
        RECT 207.620 18.350 207.760 386.250 ;
        RECT 38.280 18.030 38.540 18.350 ;
        RECT 207.560 18.030 207.820 18.350 ;
        RECT 38.340 2.400 38.480 18.030 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 239.270 15.200 239.590 15.260 ;
        RECT 270.090 15.200 270.410 15.260 ;
        RECT 239.270 15.060 270.410 15.200 ;
        RECT 239.270 15.000 239.590 15.060 ;
        RECT 270.090 15.000 270.410 15.060 ;
      LAYER via ;
        RECT 239.300 15.000 239.560 15.260 ;
        RECT 270.120 15.000 270.380 15.260 ;
      LAYER met2 ;
        RECT 273.230 400.250 273.510 404.000 ;
        RECT 272.020 400.110 273.510 400.250 ;
        RECT 272.020 324.370 272.160 400.110 ;
        RECT 273.230 400.000 273.510 400.110 ;
        RECT 270.180 324.230 272.160 324.370 ;
        RECT 270.180 15.290 270.320 324.230 ;
        RECT 239.300 14.970 239.560 15.290 ;
        RECT 270.120 14.970 270.380 15.290 ;
        RECT 239.360 2.400 239.500 14.970 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 257.670 388.520 257.990 388.580 ;
        RECT 278.830 388.520 279.150 388.580 ;
        RECT 257.670 388.380 279.150 388.520 ;
        RECT 257.670 388.320 257.990 388.380 ;
        RECT 278.830 388.320 279.150 388.380 ;
      LAYER via ;
        RECT 257.700 388.320 257.960 388.580 ;
        RECT 278.860 388.320 279.120 388.580 ;
      LAYER met2 ;
        RECT 278.750 400.180 279.030 404.000 ;
        RECT 278.750 400.000 279.060 400.180 ;
        RECT 278.920 388.610 279.060 400.000 ;
        RECT 257.700 388.290 257.960 388.610 ;
        RECT 278.860 388.290 279.120 388.610 ;
        RECT 257.760 324.370 257.900 388.290 ;
        RECT 256.840 324.230 257.900 324.370 ;
        RECT 256.840 2.400 256.980 324.230 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.690 20.640 275.010 20.700 ;
        RECT 284.350 20.640 284.670 20.700 ;
        RECT 274.690 20.500 284.670 20.640 ;
        RECT 274.690 20.440 275.010 20.500 ;
        RECT 284.350 20.440 284.670 20.500 ;
      LAYER via ;
        RECT 274.720 20.440 274.980 20.700 ;
        RECT 284.380 20.440 284.640 20.700 ;
      LAYER met2 ;
        RECT 284.270 400.250 284.550 404.000 ;
        RECT 283.980 400.110 284.550 400.250 ;
        RECT 283.980 82.870 284.120 400.110 ;
        RECT 284.270 400.000 284.550 400.110 ;
        RECT 283.980 82.730 284.580 82.870 ;
        RECT 284.440 20.730 284.580 82.730 ;
        RECT 274.720 20.410 274.980 20.730 ;
        RECT 284.380 20.410 284.640 20.730 ;
        RECT 274.780 2.400 274.920 20.410 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.790 400.180 290.070 404.000 ;
        RECT 289.790 400.000 290.100 400.180 ;
        RECT 289.960 17.410 290.100 400.000 ;
        RECT 289.960 17.270 292.400 17.410 ;
        RECT 292.260 2.400 292.400 17.270 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.790 386.480 291.110 386.540 ;
        RECT 294.010 386.480 294.330 386.540 ;
        RECT 290.790 386.340 294.330 386.480 ;
        RECT 290.790 386.280 291.110 386.340 ;
        RECT 294.010 386.280 294.330 386.340 ;
        RECT 290.790 18.600 291.110 18.660 ;
        RECT 310.110 18.600 310.430 18.660 ;
        RECT 290.790 18.460 310.430 18.600 ;
        RECT 290.790 18.400 291.110 18.460 ;
        RECT 310.110 18.400 310.430 18.460 ;
      LAYER via ;
        RECT 290.820 386.280 291.080 386.540 ;
        RECT 294.040 386.280 294.300 386.540 ;
        RECT 290.820 18.400 291.080 18.660 ;
        RECT 310.140 18.400 310.400 18.660 ;
      LAYER met2 ;
        RECT 295.310 400.250 295.590 404.000 ;
        RECT 294.100 400.110 295.590 400.250 ;
        RECT 294.100 386.570 294.240 400.110 ;
        RECT 295.310 400.000 295.590 400.110 ;
        RECT 290.820 386.250 291.080 386.570 ;
        RECT 294.040 386.250 294.300 386.570 ;
        RECT 290.880 18.690 291.020 386.250 ;
        RECT 290.820 18.370 291.080 18.690 ;
        RECT 310.140 18.370 310.400 18.690 ;
        RECT 310.200 2.400 310.340 18.370 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.450 386.480 300.770 386.540 ;
        RECT 306.890 386.480 307.210 386.540 ;
        RECT 300.450 386.340 307.210 386.480 ;
        RECT 300.450 386.280 300.770 386.340 ;
        RECT 306.890 386.280 307.210 386.340 ;
        RECT 306.890 15.200 307.210 15.260 ;
        RECT 327.590 15.200 327.910 15.260 ;
        RECT 306.890 15.060 327.910 15.200 ;
        RECT 306.890 15.000 307.210 15.060 ;
        RECT 327.590 15.000 327.910 15.060 ;
      LAYER via ;
        RECT 300.480 386.280 300.740 386.540 ;
        RECT 306.920 386.280 307.180 386.540 ;
        RECT 306.920 15.000 307.180 15.260 ;
        RECT 327.620 15.000 327.880 15.260 ;
      LAYER met2 ;
        RECT 300.370 400.180 300.650 404.000 ;
        RECT 300.370 400.000 300.680 400.180 ;
        RECT 300.540 386.570 300.680 400.000 ;
        RECT 300.480 386.250 300.740 386.570 ;
        RECT 306.920 386.250 307.180 386.570 ;
        RECT 306.980 15.290 307.120 386.250 ;
        RECT 306.920 14.970 307.180 15.290 ;
        RECT 327.620 14.970 327.880 15.290 ;
        RECT 327.680 2.400 327.820 14.970 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.130 19.280 304.450 19.340 ;
        RECT 304.130 19.140 319.540 19.280 ;
        RECT 304.130 19.080 304.450 19.140 ;
        RECT 319.400 18.260 319.540 19.140 ;
        RECT 345.530 18.260 345.850 18.320 ;
        RECT 319.400 18.120 345.850 18.260 ;
        RECT 345.530 18.060 345.850 18.120 ;
      LAYER via ;
        RECT 304.160 19.080 304.420 19.340 ;
        RECT 345.560 18.060 345.820 18.320 ;
      LAYER met2 ;
        RECT 305.890 400.250 306.170 404.000 ;
        RECT 304.680 400.110 306.170 400.250 ;
        RECT 304.680 351.970 304.820 400.110 ;
        RECT 305.890 400.000 306.170 400.110 ;
        RECT 304.220 351.830 304.820 351.970 ;
        RECT 304.220 19.370 304.360 351.830 ;
        RECT 304.160 19.050 304.420 19.370 ;
        RECT 345.560 18.030 345.820 18.350 ;
        RECT 345.620 2.400 345.760 18.030 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.570 18.600 310.890 18.660 ;
        RECT 310.570 18.460 319.080 18.600 ;
        RECT 310.570 18.400 310.890 18.460 ;
        RECT 318.940 17.920 319.080 18.460 ;
        RECT 363.010 17.920 363.330 17.980 ;
        RECT 318.940 17.780 363.330 17.920 ;
        RECT 363.010 17.720 363.330 17.780 ;
      LAYER via ;
        RECT 310.600 18.400 310.860 18.660 ;
        RECT 363.040 17.720 363.300 17.980 ;
      LAYER met2 ;
        RECT 311.410 400.250 311.690 404.000 ;
        RECT 310.660 400.110 311.690 400.250 ;
        RECT 310.660 18.690 310.800 400.110 ;
        RECT 311.410 400.000 311.690 400.110 ;
        RECT 310.600 18.370 310.860 18.690 ;
        RECT 363.040 17.690 363.300 18.010 ;
        RECT 363.100 2.400 363.240 17.690 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.570 392.260 379.890 392.320 ;
        RECT 351.830 392.120 379.890 392.260 ;
        RECT 317.010 391.920 317.330 391.980 ;
        RECT 351.830 391.920 351.970 392.120 ;
        RECT 379.570 392.060 379.890 392.120 ;
        RECT 317.010 391.780 351.970 391.920 ;
        RECT 317.010 391.720 317.330 391.780 ;
      LAYER via ;
        RECT 317.040 391.720 317.300 391.980 ;
        RECT 379.600 392.060 379.860 392.320 ;
      LAYER met2 ;
        RECT 316.930 400.180 317.210 404.000 ;
        RECT 316.930 400.000 317.240 400.180 ;
        RECT 317.100 392.010 317.240 400.000 ;
        RECT 379.600 392.030 379.860 392.350 ;
        RECT 317.040 391.690 317.300 392.010 ;
        RECT 379.660 1.770 379.800 392.030 ;
        RECT 380.830 1.770 381.390 2.400 ;
        RECT 379.660 1.630 381.390 1.770 ;
        RECT 380.830 -4.800 381.390 1.630 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.850 26.080 319.170 26.140 ;
        RECT 398.430 26.080 398.750 26.140 ;
        RECT 318.850 25.940 398.750 26.080 ;
        RECT 318.850 25.880 319.170 25.940 ;
        RECT 398.430 25.880 398.750 25.940 ;
      LAYER via ;
        RECT 318.880 25.880 319.140 26.140 ;
        RECT 398.460 25.880 398.720 26.140 ;
      LAYER met2 ;
        RECT 322.450 400.250 322.730 404.000 ;
        RECT 321.240 400.110 322.730 400.250 ;
        RECT 321.240 324.370 321.380 400.110 ;
        RECT 322.450 400.000 322.730 400.110 ;
        RECT 318.940 324.230 321.380 324.370 ;
        RECT 318.940 26.170 319.080 324.230 ;
        RECT 318.880 25.850 319.140 26.170 ;
        RECT 398.460 25.850 398.720 26.170 ;
        RECT 398.520 2.400 398.660 25.850 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 61.710 19.280 62.030 19.340 ;
        RECT 214.890 19.280 215.210 19.340 ;
        RECT 61.710 19.140 215.210 19.280 ;
        RECT 61.710 19.080 62.030 19.140 ;
        RECT 214.890 19.080 215.210 19.140 ;
      LAYER via ;
        RECT 61.740 19.080 62.000 19.340 ;
        RECT 214.920 19.080 215.180 19.340 ;
      LAYER met2 ;
        RECT 218.490 400.250 218.770 404.000 ;
        RECT 217.280 400.110 218.770 400.250 ;
        RECT 217.280 324.370 217.420 400.110 ;
        RECT 218.490 400.000 218.770 400.110 ;
        RECT 214.980 324.230 217.420 324.370 ;
        RECT 214.980 19.370 215.120 324.230 ;
        RECT 61.740 19.050 62.000 19.370 ;
        RECT 214.920 19.050 215.180 19.370 ;
        RECT 61.800 2.400 61.940 19.050 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 325.290 25.740 325.610 25.800 ;
        RECT 416.370 25.740 416.690 25.800 ;
        RECT 325.290 25.600 416.690 25.740 ;
        RECT 325.290 25.540 325.610 25.600 ;
        RECT 416.370 25.540 416.690 25.600 ;
      LAYER via ;
        RECT 325.320 25.540 325.580 25.800 ;
        RECT 416.400 25.540 416.660 25.800 ;
      LAYER met2 ;
        RECT 327.970 400.250 328.250 404.000 ;
        RECT 326.760 400.110 328.250 400.250 ;
        RECT 326.760 324.370 326.900 400.110 ;
        RECT 327.970 400.000 328.250 400.110 ;
        RECT 325.380 324.230 326.900 324.370 ;
        RECT 325.380 25.830 325.520 324.230 ;
        RECT 325.320 25.510 325.580 25.830 ;
        RECT 416.400 25.510 416.660 25.830 ;
        RECT 416.460 2.400 416.600 25.510 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 332.190 25.400 332.510 25.460 ;
        RECT 434.310 25.400 434.630 25.460 ;
        RECT 332.190 25.260 434.630 25.400 ;
        RECT 332.190 25.200 332.510 25.260 ;
        RECT 434.310 25.200 434.630 25.260 ;
      LAYER via ;
        RECT 332.220 25.200 332.480 25.460 ;
        RECT 434.340 25.200 434.600 25.460 ;
      LAYER met2 ;
        RECT 333.490 400.250 333.770 404.000 ;
        RECT 332.280 400.110 333.770 400.250 ;
        RECT 332.280 25.490 332.420 400.110 ;
        RECT 333.490 400.000 333.770 400.110 ;
        RECT 332.220 25.170 332.480 25.490 ;
        RECT 434.340 25.170 434.600 25.490 ;
        RECT 434.400 2.400 434.540 25.170 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 338.630 25.060 338.950 25.120 ;
        RECT 451.790 25.060 452.110 25.120 ;
        RECT 338.630 24.920 452.110 25.060 ;
        RECT 338.630 24.860 338.950 24.920 ;
        RECT 451.790 24.860 452.110 24.920 ;
      LAYER via ;
        RECT 338.660 24.860 338.920 25.120 ;
        RECT 451.820 24.860 452.080 25.120 ;
      LAYER met2 ;
        RECT 339.010 400.250 339.290 404.000 ;
        RECT 338.720 400.110 339.290 400.250 ;
        RECT 338.720 25.150 338.860 400.110 ;
        RECT 339.010 400.000 339.290 400.110 ;
        RECT 338.660 24.830 338.920 25.150 ;
        RECT 451.820 24.830 452.080 25.150 ;
        RECT 451.880 2.400 452.020 24.830 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 339.090 376.280 339.410 376.340 ;
        RECT 343.230 376.280 343.550 376.340 ;
        RECT 339.090 376.140 343.550 376.280 ;
        RECT 339.090 376.080 339.410 376.140 ;
        RECT 343.230 376.080 343.550 376.140 ;
        RECT 339.090 24.380 339.410 24.440 ;
        RECT 469.730 24.380 470.050 24.440 ;
        RECT 339.090 24.240 470.050 24.380 ;
        RECT 339.090 24.180 339.410 24.240 ;
        RECT 469.730 24.180 470.050 24.240 ;
      LAYER via ;
        RECT 339.120 376.080 339.380 376.340 ;
        RECT 343.260 376.080 343.520 376.340 ;
        RECT 339.120 24.180 339.380 24.440 ;
        RECT 469.760 24.180 470.020 24.440 ;
      LAYER met2 ;
        RECT 344.070 400.250 344.350 404.000 ;
        RECT 343.320 400.110 344.350 400.250 ;
        RECT 343.320 376.370 343.460 400.110 ;
        RECT 344.070 400.000 344.350 400.110 ;
        RECT 339.120 376.050 339.380 376.370 ;
        RECT 343.260 376.050 343.520 376.370 ;
        RECT 339.180 24.470 339.320 376.050 ;
        RECT 339.120 24.150 339.380 24.470 ;
        RECT 469.760 24.150 470.020 24.470 ;
        RECT 469.820 2.400 469.960 24.150 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 349.670 388.180 349.990 388.240 ;
        RECT 403.490 388.180 403.810 388.240 ;
        RECT 349.670 388.040 403.810 388.180 ;
        RECT 349.670 387.980 349.990 388.040 ;
        RECT 403.490 387.980 403.810 388.040 ;
        RECT 403.490 16.560 403.810 16.620 ;
        RECT 403.490 16.420 445.120 16.560 ;
        RECT 403.490 16.360 403.810 16.420 ;
        RECT 444.980 15.880 445.120 16.420 ;
        RECT 487.210 15.880 487.530 15.940 ;
        RECT 444.980 15.740 487.530 15.880 ;
        RECT 487.210 15.680 487.530 15.740 ;
      LAYER via ;
        RECT 349.700 387.980 349.960 388.240 ;
        RECT 403.520 387.980 403.780 388.240 ;
        RECT 403.520 16.360 403.780 16.620 ;
        RECT 487.240 15.680 487.500 15.940 ;
      LAYER met2 ;
        RECT 349.590 400.180 349.870 404.000 ;
        RECT 349.590 400.000 349.900 400.180 ;
        RECT 349.760 388.270 349.900 400.000 ;
        RECT 349.700 387.950 349.960 388.270 ;
        RECT 403.520 387.950 403.780 388.270 ;
        RECT 403.580 16.650 403.720 387.950 ;
        RECT 403.520 16.330 403.780 16.650 ;
        RECT 487.240 15.650 487.500 15.970 ;
        RECT 487.300 2.400 487.440 15.650 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 355.190 387.840 355.510 387.900 ;
        RECT 389.690 387.840 390.010 387.900 ;
        RECT 355.190 387.700 390.010 387.840 ;
        RECT 355.190 387.640 355.510 387.700 ;
        RECT 389.690 387.640 390.010 387.700 ;
        RECT 389.690 17.240 390.010 17.300 ;
        RECT 389.690 17.100 445.120 17.240 ;
        RECT 389.690 17.040 390.010 17.100 ;
        RECT 444.980 16.900 445.120 17.100 ;
        RECT 444.980 16.760 469.270 16.900 ;
        RECT 469.130 16.560 469.270 16.760 ;
        RECT 505.150 16.560 505.470 16.620 ;
        RECT 469.130 16.420 505.470 16.560 ;
        RECT 505.150 16.360 505.470 16.420 ;
      LAYER via ;
        RECT 355.220 387.640 355.480 387.900 ;
        RECT 389.720 387.640 389.980 387.900 ;
        RECT 389.720 17.040 389.980 17.300 ;
        RECT 505.180 16.360 505.440 16.620 ;
      LAYER met2 ;
        RECT 355.110 400.180 355.390 404.000 ;
        RECT 355.110 400.000 355.420 400.180 ;
        RECT 355.280 387.930 355.420 400.000 ;
        RECT 355.220 387.610 355.480 387.930 ;
        RECT 389.720 387.610 389.980 387.930 ;
        RECT 389.780 17.330 389.920 387.610 ;
        RECT 389.720 17.010 389.980 17.330 ;
        RECT 505.180 16.330 505.440 16.650 ;
        RECT 505.240 2.400 505.380 16.330 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.710 391.240 361.030 391.300 ;
        RECT 479.390 391.240 479.710 391.300 ;
        RECT 360.710 391.100 479.710 391.240 ;
        RECT 360.710 391.040 361.030 391.100 ;
        RECT 479.390 391.040 479.710 391.100 ;
        RECT 479.390 16.900 479.710 16.960 ;
        RECT 511.590 16.900 511.910 16.960 ;
        RECT 479.390 16.760 511.910 16.900 ;
        RECT 479.390 16.700 479.710 16.760 ;
        RECT 511.590 16.700 511.910 16.760 ;
        RECT 512.510 16.900 512.830 16.960 ;
        RECT 522.630 16.900 522.950 16.960 ;
        RECT 512.510 16.760 522.950 16.900 ;
        RECT 512.510 16.700 512.830 16.760 ;
        RECT 522.630 16.700 522.950 16.760 ;
      LAYER via ;
        RECT 360.740 391.040 361.000 391.300 ;
        RECT 479.420 391.040 479.680 391.300 ;
        RECT 479.420 16.700 479.680 16.960 ;
        RECT 511.620 16.700 511.880 16.960 ;
        RECT 512.540 16.700 512.800 16.960 ;
        RECT 522.660 16.700 522.920 16.960 ;
      LAYER met2 ;
        RECT 360.630 400.180 360.910 404.000 ;
        RECT 360.630 400.000 360.940 400.180 ;
        RECT 360.800 391.330 360.940 400.000 ;
        RECT 360.740 391.010 361.000 391.330 ;
        RECT 479.420 391.010 479.680 391.330 ;
        RECT 479.480 16.990 479.620 391.010 ;
        RECT 479.420 16.670 479.680 16.990 ;
        RECT 511.620 16.730 511.880 16.990 ;
        RECT 512.540 16.730 512.800 16.990 ;
        RECT 511.620 16.670 512.800 16.730 ;
        RECT 522.660 16.670 522.920 16.990 ;
        RECT 511.680 16.590 512.740 16.670 ;
        RECT 522.720 2.400 522.860 16.670 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.230 389.200 366.550 389.260 ;
        RECT 410.390 389.200 410.710 389.260 ;
        RECT 366.230 389.060 410.710 389.200 ;
        RECT 366.230 389.000 366.550 389.060 ;
        RECT 410.390 389.000 410.710 389.060 ;
        RECT 416.920 20.840 421.660 20.980 ;
        RECT 410.850 20.640 411.170 20.700 ;
        RECT 416.920 20.640 417.060 20.840 ;
        RECT 410.850 20.500 417.060 20.640 ;
        RECT 421.520 20.640 421.660 20.840 ;
        RECT 540.570 20.640 540.890 20.700 ;
        RECT 421.520 20.500 540.890 20.640 ;
        RECT 410.850 20.440 411.170 20.500 ;
        RECT 540.570 20.440 540.890 20.500 ;
      LAYER via ;
        RECT 366.260 389.000 366.520 389.260 ;
        RECT 410.420 389.000 410.680 389.260 ;
        RECT 410.880 20.440 411.140 20.700 ;
        RECT 540.600 20.440 540.860 20.700 ;
      LAYER met2 ;
        RECT 366.150 400.180 366.430 404.000 ;
        RECT 366.150 400.000 366.460 400.180 ;
        RECT 366.320 389.290 366.460 400.000 ;
        RECT 366.260 388.970 366.520 389.290 ;
        RECT 410.420 388.970 410.680 389.290 ;
        RECT 410.480 82.870 410.620 388.970 ;
        RECT 410.480 82.730 411.080 82.870 ;
        RECT 410.940 20.730 411.080 82.730 ;
        RECT 410.880 20.410 411.140 20.730 ;
        RECT 540.600 20.410 540.860 20.730 ;
        RECT 540.660 2.400 540.800 20.410 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 371.750 390.220 372.070 390.280 ;
        RECT 486.290 390.220 486.610 390.280 ;
        RECT 371.750 390.080 486.610 390.220 ;
        RECT 371.750 390.020 372.070 390.080 ;
        RECT 486.290 390.020 486.610 390.080 ;
        RECT 486.290 14.860 486.610 14.920 ;
        RECT 486.290 14.720 517.570 14.860 ;
        RECT 486.290 14.660 486.610 14.720 ;
        RECT 517.430 14.520 517.570 14.720 ;
        RECT 558.050 14.520 558.370 14.580 ;
        RECT 517.430 14.380 558.370 14.520 ;
        RECT 558.050 14.320 558.370 14.380 ;
      LAYER via ;
        RECT 371.780 390.020 372.040 390.280 ;
        RECT 486.320 390.020 486.580 390.280 ;
        RECT 486.320 14.660 486.580 14.920 ;
        RECT 558.080 14.320 558.340 14.580 ;
      LAYER met2 ;
        RECT 371.670 400.180 371.950 404.000 ;
        RECT 371.670 400.000 371.980 400.180 ;
        RECT 371.840 390.310 371.980 400.000 ;
        RECT 371.780 389.990 372.040 390.310 ;
        RECT 486.320 389.990 486.580 390.310 ;
        RECT 486.380 14.950 486.520 389.990 ;
        RECT 486.320 14.630 486.580 14.950 ;
        RECT 558.080 14.290 558.340 14.610 ;
        RECT 558.140 2.400 558.280 14.290 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 386.480 372.990 386.540 ;
        RECT 375.890 386.480 376.210 386.540 ;
        RECT 372.670 386.340 376.210 386.480 ;
        RECT 372.670 386.280 372.990 386.340 ;
        RECT 375.890 386.280 376.210 386.340 ;
        RECT 398.890 18.940 399.210 19.000 ;
        RECT 575.990 18.940 576.310 19.000 ;
        RECT 398.890 18.800 576.310 18.940 ;
        RECT 398.890 18.740 399.210 18.800 ;
        RECT 575.990 18.740 576.310 18.800 ;
        RECT 372.670 14.860 372.990 14.920 ;
        RECT 398.890 14.860 399.210 14.920 ;
        RECT 372.670 14.720 399.210 14.860 ;
        RECT 372.670 14.660 372.990 14.720 ;
        RECT 398.890 14.660 399.210 14.720 ;
      LAYER via ;
        RECT 372.700 386.280 372.960 386.540 ;
        RECT 375.920 386.280 376.180 386.540 ;
        RECT 398.920 18.740 399.180 19.000 ;
        RECT 576.020 18.740 576.280 19.000 ;
        RECT 372.700 14.660 372.960 14.920 ;
        RECT 398.920 14.660 399.180 14.920 ;
      LAYER met2 ;
        RECT 377.190 400.250 377.470 404.000 ;
        RECT 375.980 400.110 377.470 400.250 ;
        RECT 375.980 386.570 376.120 400.110 ;
        RECT 377.190 400.000 377.470 400.110 ;
        RECT 372.700 386.250 372.960 386.570 ;
        RECT 375.920 386.250 376.180 386.570 ;
        RECT 372.760 14.950 372.900 386.250 ;
        RECT 398.920 18.710 399.180 19.030 ;
        RECT 576.020 18.710 576.280 19.030 ;
        RECT 398.980 14.950 399.120 18.710 ;
        RECT 372.700 14.630 372.960 14.950 ;
        RECT 398.920 14.630 399.180 14.950 ;
        RECT 576.080 2.400 576.220 18.710 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 85.170 19.960 85.490 20.020 ;
        RECT 221.330 19.960 221.650 20.020 ;
        RECT 85.170 19.820 221.650 19.960 ;
        RECT 85.170 19.760 85.490 19.820 ;
        RECT 221.330 19.760 221.650 19.820 ;
      LAYER via ;
        RECT 85.200 19.760 85.460 20.020 ;
        RECT 221.360 19.760 221.620 20.020 ;
      LAYER met2 ;
        RECT 225.850 400.250 226.130 404.000 ;
        RECT 224.640 400.110 226.130 400.250 ;
        RECT 224.640 390.730 224.780 400.110 ;
        RECT 225.850 400.000 226.130 400.110 ;
        RECT 221.420 390.590 224.780 390.730 ;
        RECT 221.420 20.050 221.560 390.590 ;
        RECT 85.200 19.730 85.460 20.050 ;
        RECT 221.360 19.730 221.620 20.050 ;
        RECT 85.260 2.400 85.400 19.730 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.950 18.940 381.270 19.000 ;
        RECT 380.950 18.800 398.660 18.940 ;
        RECT 380.950 18.740 381.270 18.800 ;
        RECT 398.520 18.600 398.660 18.800 ;
        RECT 593.930 18.600 594.250 18.660 ;
        RECT 398.520 18.460 594.250 18.600 ;
        RECT 593.930 18.400 594.250 18.460 ;
      LAYER via ;
        RECT 380.980 18.740 381.240 19.000 ;
        RECT 593.960 18.400 594.220 18.660 ;
      LAYER met2 ;
        RECT 382.710 400.250 382.990 404.000 ;
        RECT 381.500 400.110 382.990 400.250 ;
        RECT 381.500 324.370 381.640 400.110 ;
        RECT 382.710 400.000 382.990 400.110 ;
        RECT 381.040 324.230 381.640 324.370 ;
        RECT 381.040 19.030 381.180 324.230 ;
        RECT 380.980 18.710 381.240 19.030 ;
        RECT 593.960 18.370 594.220 18.690 ;
        RECT 594.020 2.400 594.160 18.370 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 388.310 387.500 388.630 387.560 ;
        RECT 493.190 387.500 493.510 387.560 ;
        RECT 388.310 387.360 493.510 387.500 ;
        RECT 388.310 387.300 388.630 387.360 ;
        RECT 493.190 387.300 493.510 387.360 ;
        RECT 547.010 20.300 547.330 20.360 ;
        RECT 611.410 20.300 611.730 20.360 ;
        RECT 547.010 20.160 611.730 20.300 ;
        RECT 547.010 20.100 547.330 20.160 ;
        RECT 611.410 20.100 611.730 20.160 ;
        RECT 547.010 16.220 547.330 16.280 ;
        RECT 512.140 16.080 547.330 16.220 ;
        RECT 493.650 15.880 493.970 15.940 ;
        RECT 512.140 15.880 512.280 16.080 ;
        RECT 547.010 16.020 547.330 16.080 ;
        RECT 493.650 15.740 512.280 15.880 ;
        RECT 493.650 15.680 493.970 15.740 ;
      LAYER via ;
        RECT 388.340 387.300 388.600 387.560 ;
        RECT 493.220 387.300 493.480 387.560 ;
        RECT 547.040 20.100 547.300 20.360 ;
        RECT 611.440 20.100 611.700 20.360 ;
        RECT 493.680 15.680 493.940 15.940 ;
        RECT 547.040 16.020 547.300 16.280 ;
      LAYER met2 ;
        RECT 388.230 400.180 388.510 404.000 ;
        RECT 388.230 400.000 388.540 400.180 ;
        RECT 388.400 387.590 388.540 400.000 ;
        RECT 388.340 387.270 388.600 387.590 ;
        RECT 493.220 387.270 493.480 387.590 ;
        RECT 493.280 82.870 493.420 387.270 ;
        RECT 493.280 82.730 493.880 82.870 ;
        RECT 493.740 15.970 493.880 82.730 ;
        RECT 547.040 20.070 547.300 20.390 ;
        RECT 611.440 20.070 611.700 20.390 ;
        RECT 547.100 16.310 547.240 20.070 ;
        RECT 547.040 15.990 547.300 16.310 ;
        RECT 493.680 15.650 493.940 15.970 ;
        RECT 611.500 2.400 611.640 20.070 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 109.090 24.040 109.410 24.100 ;
        RECT 229.150 24.040 229.470 24.100 ;
        RECT 109.090 23.900 229.470 24.040 ;
        RECT 109.090 23.840 109.410 23.900 ;
        RECT 229.150 23.840 229.470 23.900 ;
      LAYER via ;
        RECT 109.120 23.840 109.380 24.100 ;
        RECT 229.180 23.840 229.440 24.100 ;
      LAYER met2 ;
        RECT 233.210 400.250 233.490 404.000 ;
        RECT 232.000 400.110 233.490 400.250 ;
        RECT 232.000 324.370 232.140 400.110 ;
        RECT 233.210 400.000 233.490 400.110 ;
        RECT 229.240 324.230 232.140 324.370 ;
        RECT 229.240 24.130 229.380 324.230 ;
        RECT 109.120 23.810 109.380 24.130 ;
        RECT 229.180 23.810 229.440 24.130 ;
        RECT 109.180 2.400 109.320 23.810 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.550 24.380 132.870 24.440 ;
        RECT 235.590 24.380 235.910 24.440 ;
        RECT 132.550 24.240 235.910 24.380 ;
        RECT 132.550 24.180 132.870 24.240 ;
        RECT 235.590 24.180 235.910 24.240 ;
      LAYER via ;
        RECT 132.580 24.180 132.840 24.440 ;
        RECT 235.620 24.180 235.880 24.440 ;
      LAYER met2 ;
        RECT 240.570 400.250 240.850 404.000 ;
        RECT 239.360 400.110 240.850 400.250 ;
        RECT 239.360 324.370 239.500 400.110 ;
        RECT 240.570 400.000 240.850 400.110 ;
        RECT 235.680 324.230 239.500 324.370 ;
        RECT 235.680 24.470 235.820 324.230 ;
        RECT 132.580 24.150 132.840 24.470 ;
        RECT 235.620 24.150 235.880 24.470 ;
        RECT 132.640 2.400 132.780 24.150 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.490 386.480 242.810 386.540 ;
        RECT 244.790 386.480 245.110 386.540 ;
        RECT 242.490 386.340 245.110 386.480 ;
        RECT 242.490 386.280 242.810 386.340 ;
        RECT 244.790 386.280 245.110 386.340 ;
        RECT 150.490 24.720 150.810 24.780 ;
        RECT 242.490 24.720 242.810 24.780 ;
        RECT 150.490 24.580 242.810 24.720 ;
        RECT 150.490 24.520 150.810 24.580 ;
        RECT 242.490 24.520 242.810 24.580 ;
      LAYER via ;
        RECT 242.520 386.280 242.780 386.540 ;
        RECT 244.820 386.280 245.080 386.540 ;
        RECT 150.520 24.520 150.780 24.780 ;
        RECT 242.520 24.520 242.780 24.780 ;
      LAYER met2 ;
        RECT 246.090 400.250 246.370 404.000 ;
        RECT 244.880 400.110 246.370 400.250 ;
        RECT 244.880 386.570 245.020 400.110 ;
        RECT 246.090 400.000 246.370 400.110 ;
        RECT 242.520 386.250 242.780 386.570 ;
        RECT 244.820 386.250 245.080 386.570 ;
        RECT 242.580 24.810 242.720 386.250 ;
        RECT 150.520 24.490 150.780 24.810 ;
        RECT 242.520 24.490 242.780 24.810 ;
        RECT 150.580 2.400 150.720 24.490 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 165.670 393.280 165.990 393.340 ;
        RECT 251.230 393.280 251.550 393.340 ;
        RECT 165.670 393.140 251.550 393.280 ;
        RECT 165.670 393.080 165.990 393.140 ;
        RECT 251.230 393.080 251.550 393.140 ;
      LAYER via ;
        RECT 165.700 393.080 165.960 393.340 ;
        RECT 251.260 393.080 251.520 393.340 ;
      LAYER met2 ;
        RECT 251.150 400.180 251.430 404.000 ;
        RECT 251.150 400.000 251.460 400.180 ;
        RECT 251.320 393.370 251.460 400.000 ;
        RECT 165.700 393.050 165.960 393.370 ;
        RECT 251.260 393.050 251.520 393.370 ;
        RECT 165.760 82.870 165.900 393.050 ;
        RECT 165.760 82.730 168.200 82.870 ;
        RECT 168.060 2.400 168.200 82.730 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 179.470 389.540 179.790 389.600 ;
        RECT 256.750 389.540 257.070 389.600 ;
        RECT 179.470 389.400 257.070 389.540 ;
        RECT 179.470 389.340 179.790 389.400 ;
        RECT 256.750 389.340 257.070 389.400 ;
      LAYER via ;
        RECT 179.500 389.340 179.760 389.600 ;
        RECT 256.780 389.340 257.040 389.600 ;
      LAYER met2 ;
        RECT 256.670 400.180 256.950 404.000 ;
        RECT 256.670 400.000 256.980 400.180 ;
        RECT 256.840 389.630 256.980 400.000 ;
        RECT 179.500 389.310 179.760 389.630 ;
        RECT 256.780 389.310 257.040 389.630 ;
        RECT 179.560 82.870 179.700 389.310 ;
        RECT 179.560 82.730 183.840 82.870 ;
        RECT 183.700 1.770 183.840 82.730 ;
        RECT 185.790 1.770 186.350 2.400 ;
        RECT 183.700 1.630 186.350 1.770 ;
        RECT 185.790 -4.800 186.350 1.630 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203.390 15.200 203.710 15.260 ;
        RECT 203.390 15.060 227.770 15.200 ;
        RECT 203.390 15.000 203.710 15.060 ;
        RECT 227.630 14.860 227.770 15.060 ;
        RECT 263.650 14.860 263.970 14.920 ;
        RECT 227.630 14.720 263.970 14.860 ;
        RECT 263.650 14.660 263.970 14.720 ;
      LAYER via ;
        RECT 203.420 15.000 203.680 15.260 ;
        RECT 263.680 14.660 263.940 14.920 ;
      LAYER met2 ;
        RECT 262.190 400.250 262.470 404.000 ;
        RECT 262.190 400.110 263.420 400.250 ;
        RECT 262.190 400.000 262.470 400.110 ;
        RECT 263.280 82.870 263.420 400.110 ;
        RECT 263.280 82.730 263.880 82.870 ;
        RECT 203.420 14.970 203.680 15.290 ;
        RECT 203.480 2.400 203.620 14.970 ;
        RECT 263.740 14.950 263.880 82.730 ;
        RECT 263.680 14.630 263.940 14.950 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.730 386.480 263.050 386.540 ;
        RECT 266.410 386.480 266.730 386.540 ;
        RECT 262.730 386.340 266.730 386.480 ;
        RECT 262.730 386.280 263.050 386.340 ;
        RECT 266.410 386.280 266.730 386.340 ;
        RECT 262.730 17.920 263.050 17.980 ;
        RECT 232.920 17.780 263.050 17.920 ;
        RECT 221.330 17.240 221.650 17.300 ;
        RECT 232.920 17.240 233.060 17.780 ;
        RECT 262.730 17.720 263.050 17.780 ;
        RECT 221.330 17.100 233.060 17.240 ;
        RECT 221.330 17.040 221.650 17.100 ;
      LAYER via ;
        RECT 262.760 386.280 263.020 386.540 ;
        RECT 266.440 386.280 266.700 386.540 ;
        RECT 221.360 17.040 221.620 17.300 ;
        RECT 262.760 17.720 263.020 17.980 ;
      LAYER met2 ;
        RECT 267.710 400.250 267.990 404.000 ;
        RECT 266.500 400.110 267.990 400.250 ;
        RECT 266.500 386.570 266.640 400.110 ;
        RECT 267.710 400.000 267.990 400.110 ;
        RECT 262.760 386.250 263.020 386.570 ;
        RECT 266.440 386.250 266.700 386.570 ;
        RECT 262.820 18.010 262.960 386.250 ;
        RECT 262.760 17.690 263.020 18.010 ;
        RECT 221.360 17.010 221.620 17.330 ;
        RECT 221.420 2.400 221.560 17.010 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.630 375.940 200.950 376.000 ;
        RECT 204.310 375.940 204.630 376.000 ;
        RECT 200.630 375.800 204.630 375.940 ;
        RECT 200.630 375.740 200.950 375.800 ;
        RECT 204.310 375.740 204.630 375.800 ;
        RECT 20.310 17.920 20.630 17.980 ;
        RECT 200.630 17.920 200.950 17.980 ;
        RECT 20.310 17.780 200.950 17.920 ;
        RECT 20.310 17.720 20.630 17.780 ;
        RECT 200.630 17.720 200.950 17.780 ;
      LAYER via ;
        RECT 200.660 375.740 200.920 376.000 ;
        RECT 204.340 375.740 204.600 376.000 ;
        RECT 20.340 17.720 20.600 17.980 ;
        RECT 200.660 17.720 200.920 17.980 ;
      LAYER met2 ;
        RECT 205.610 400.250 205.890 404.000 ;
        RECT 204.400 400.110 205.890 400.250 ;
        RECT 204.400 376.030 204.540 400.110 ;
        RECT 205.610 400.000 205.890 400.110 ;
        RECT 200.660 375.710 200.920 376.030 ;
        RECT 204.340 375.710 204.600 376.030 ;
        RECT 200.720 18.010 200.860 375.710 ;
        RECT 20.340 17.690 20.600 18.010 ;
        RECT 200.660 17.690 200.920 18.010 ;
        RECT 20.400 2.400 20.540 17.690 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 43.770 18.600 44.090 18.660 ;
        RECT 208.450 18.600 208.770 18.660 ;
        RECT 43.770 18.460 208.770 18.600 ;
        RECT 43.770 18.400 44.090 18.460 ;
        RECT 208.450 18.400 208.770 18.460 ;
      LAYER via ;
        RECT 43.800 18.400 44.060 18.660 ;
        RECT 208.480 18.400 208.740 18.660 ;
      LAYER met2 ;
        RECT 212.970 400.250 213.250 404.000 ;
        RECT 211.760 400.110 213.250 400.250 ;
        RECT 211.760 324.370 211.900 400.110 ;
        RECT 212.970 400.000 213.250 400.110 ;
        RECT 208.540 324.230 211.900 324.370 ;
        RECT 208.540 18.690 208.680 324.230 ;
        RECT 43.800 18.370 44.060 18.690 ;
        RECT 208.480 18.370 208.740 18.690 ;
        RECT 43.860 2.400 44.000 18.370 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.590 387.160 258.910 387.220 ;
        RECT 275.150 387.160 275.470 387.220 ;
        RECT 258.590 387.020 275.470 387.160 ;
        RECT 258.590 386.960 258.910 387.020 ;
        RECT 275.150 386.960 275.470 387.020 ;
        RECT 244.790 17.580 245.110 17.640 ;
        RECT 258.590 17.580 258.910 17.640 ;
        RECT 244.790 17.440 258.910 17.580 ;
        RECT 244.790 17.380 245.110 17.440 ;
        RECT 258.590 17.380 258.910 17.440 ;
      LAYER via ;
        RECT 258.620 386.960 258.880 387.220 ;
        RECT 275.180 386.960 275.440 387.220 ;
        RECT 244.820 17.380 245.080 17.640 ;
        RECT 258.620 17.380 258.880 17.640 ;
      LAYER met2 ;
        RECT 275.070 400.180 275.350 404.000 ;
        RECT 275.070 400.000 275.380 400.180 ;
        RECT 275.240 387.250 275.380 400.000 ;
        RECT 258.620 386.930 258.880 387.250 ;
        RECT 275.180 386.930 275.440 387.250 ;
        RECT 258.680 17.670 258.820 386.930 ;
        RECT 244.820 17.350 245.080 17.670 ;
        RECT 258.620 17.350 258.880 17.670 ;
        RECT 244.880 2.400 245.020 17.350 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.270 392.600 262.590 392.660 ;
        RECT 280.670 392.600 280.990 392.660 ;
        RECT 262.270 392.460 280.990 392.600 ;
        RECT 262.270 392.400 262.590 392.460 ;
        RECT 280.670 392.400 280.990 392.460 ;
      LAYER via ;
        RECT 262.300 392.400 262.560 392.660 ;
        RECT 280.700 392.400 280.960 392.660 ;
      LAYER met2 ;
        RECT 280.590 400.180 280.870 404.000 ;
        RECT 280.590 400.000 280.900 400.180 ;
        RECT 280.760 392.690 280.900 400.000 ;
        RECT 262.300 392.370 262.560 392.690 ;
        RECT 280.700 392.370 280.960 392.690 ;
        RECT 262.360 17.410 262.500 392.370 ;
        RECT 262.360 17.270 262.960 17.410 ;
        RECT 262.820 2.400 262.960 17.270 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 283.430 386.480 283.750 386.540 ;
        RECT 284.810 386.480 285.130 386.540 ;
        RECT 283.430 386.340 285.130 386.480 ;
        RECT 283.430 386.280 283.750 386.340 ;
        RECT 284.810 386.280 285.130 386.340 ;
      LAYER via ;
        RECT 283.460 386.280 283.720 386.540 ;
        RECT 284.840 386.280 285.100 386.540 ;
      LAYER met2 ;
        RECT 286.110 400.250 286.390 404.000 ;
        RECT 284.900 400.110 286.390 400.250 ;
        RECT 284.900 386.570 285.040 400.110 ;
        RECT 286.110 400.000 286.390 400.110 ;
        RECT 283.460 386.250 283.720 386.570 ;
        RECT 284.840 386.250 285.100 386.570 ;
        RECT 283.520 14.010 283.660 386.250 ;
        RECT 282.600 13.870 283.660 14.010 ;
        RECT 280.090 1.770 280.650 2.400 ;
        RECT 282.600 1.770 282.740 13.870 ;
        RECT 280.090 1.630 282.740 1.770 ;
        RECT 280.090 -4.800 280.650 1.630 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.330 17.920 290.650 17.980 ;
        RECT 298.150 17.920 298.470 17.980 ;
        RECT 290.330 17.780 298.470 17.920 ;
        RECT 290.330 17.720 290.650 17.780 ;
        RECT 298.150 17.720 298.470 17.780 ;
      LAYER via ;
        RECT 290.360 17.720 290.620 17.980 ;
        RECT 298.180 17.720 298.440 17.980 ;
      LAYER met2 ;
        RECT 291.630 400.250 291.910 404.000 ;
        RECT 290.420 400.110 291.910 400.250 ;
        RECT 290.420 18.010 290.560 400.110 ;
        RECT 291.630 400.000 291.910 400.110 ;
        RECT 290.360 17.690 290.620 18.010 ;
        RECT 298.180 17.690 298.440 18.010 ;
        RECT 298.240 2.400 298.380 17.690 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.770 17.580 297.090 17.640 ;
        RECT 316.090 17.580 316.410 17.640 ;
        RECT 296.770 17.440 316.410 17.580 ;
        RECT 296.770 17.380 297.090 17.440 ;
        RECT 316.090 17.380 316.410 17.440 ;
      LAYER via ;
        RECT 296.800 17.380 297.060 17.640 ;
        RECT 316.120 17.380 316.380 17.640 ;
      LAYER met2 ;
        RECT 296.690 400.180 296.970 404.000 ;
        RECT 296.690 400.000 297.000 400.180 ;
        RECT 296.860 17.670 297.000 400.000 ;
        RECT 296.800 17.350 297.060 17.670 ;
        RECT 316.120 17.350 316.380 17.670 ;
        RECT 316.180 2.400 316.320 17.350 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 297.230 14.520 297.550 14.580 ;
        RECT 333.570 14.520 333.890 14.580 ;
        RECT 297.230 14.380 333.890 14.520 ;
        RECT 297.230 14.320 297.550 14.380 ;
        RECT 333.570 14.320 333.890 14.380 ;
      LAYER via ;
        RECT 297.260 14.320 297.520 14.580 ;
        RECT 333.600 14.320 333.860 14.580 ;
      LAYER met2 ;
        RECT 302.210 400.250 302.490 404.000 ;
        RECT 301.000 400.110 302.490 400.250 ;
        RECT 301.000 324.370 301.140 400.110 ;
        RECT 302.210 400.000 302.490 400.110 ;
        RECT 297.320 324.230 301.140 324.370 ;
        RECT 297.320 14.610 297.460 324.230 ;
        RECT 297.260 14.290 297.520 14.610 ;
        RECT 333.600 14.290 333.860 14.610 ;
        RECT 333.660 2.400 333.800 14.290 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.590 19.960 304.910 20.020 ;
        RECT 304.590 19.820 320.460 19.960 ;
        RECT 304.590 19.760 304.910 19.820 ;
        RECT 320.320 18.940 320.460 19.820 ;
        RECT 351.510 18.940 351.830 19.000 ;
        RECT 320.320 18.800 351.830 18.940 ;
        RECT 351.510 18.740 351.830 18.800 ;
      LAYER via ;
        RECT 304.620 19.760 304.880 20.020 ;
        RECT 351.540 18.740 351.800 19.000 ;
      LAYER met2 ;
        RECT 307.730 400.250 308.010 404.000 ;
        RECT 306.520 400.110 308.010 400.250 ;
        RECT 306.520 324.370 306.660 400.110 ;
        RECT 307.730 400.000 308.010 400.110 ;
        RECT 304.680 324.230 306.660 324.370 ;
        RECT 304.680 20.050 304.820 324.230 ;
        RECT 304.620 19.730 304.880 20.050 ;
        RECT 351.540 18.710 351.800 19.030 ;
        RECT 351.600 2.400 351.740 18.710 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.030 18.260 311.350 18.320 ;
        RECT 311.030 18.120 318.620 18.260 ;
        RECT 311.030 18.060 311.350 18.120 ;
        RECT 318.480 17.580 318.620 18.120 ;
        RECT 368.990 17.580 369.310 17.640 ;
        RECT 318.480 17.440 369.310 17.580 ;
        RECT 368.990 17.380 369.310 17.440 ;
      LAYER via ;
        RECT 311.060 18.060 311.320 18.320 ;
        RECT 369.020 17.380 369.280 17.640 ;
      LAYER met2 ;
        RECT 313.250 400.250 313.530 404.000 ;
        RECT 312.040 400.110 313.530 400.250 ;
        RECT 312.040 324.370 312.180 400.110 ;
        RECT 313.250 400.000 313.530 400.110 ;
        RECT 311.120 324.230 312.180 324.370 ;
        RECT 311.120 18.350 311.260 324.230 ;
        RECT 311.060 18.030 311.320 18.350 ;
        RECT 369.020 17.350 369.280 17.670 ;
        RECT 369.080 2.400 369.220 17.350 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.390 20.640 318.710 20.700 ;
        RECT 322.070 20.640 322.390 20.700 ;
        RECT 318.390 20.500 322.390 20.640 ;
        RECT 318.390 20.440 318.710 20.500 ;
        RECT 322.070 20.440 322.390 20.500 ;
        RECT 322.070 15.540 322.390 15.600 ;
        RECT 386.930 15.540 387.250 15.600 ;
        RECT 322.070 15.400 387.250 15.540 ;
        RECT 322.070 15.340 322.390 15.400 ;
        RECT 386.930 15.340 387.250 15.400 ;
      LAYER via ;
        RECT 318.420 20.440 318.680 20.700 ;
        RECT 322.100 20.440 322.360 20.700 ;
        RECT 322.100 15.340 322.360 15.600 ;
        RECT 386.960 15.340 387.220 15.600 ;
      LAYER met2 ;
        RECT 318.770 400.250 319.050 404.000 ;
        RECT 318.480 400.110 319.050 400.250 ;
        RECT 318.480 20.730 318.620 400.110 ;
        RECT 318.770 400.000 319.050 400.110 ;
        RECT 318.420 20.410 318.680 20.730 ;
        RECT 322.100 20.410 322.360 20.730 ;
        RECT 322.160 15.630 322.300 20.410 ;
        RECT 322.100 15.310 322.360 15.630 ;
        RECT 386.960 15.310 387.220 15.630 ;
        RECT 387.020 2.400 387.160 15.310 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.830 17.240 325.150 17.300 ;
        RECT 358.410 17.240 358.730 17.300 ;
        RECT 324.830 17.100 358.730 17.240 ;
        RECT 324.830 17.040 325.150 17.100 ;
        RECT 358.410 17.040 358.730 17.100 ;
        RECT 358.410 15.880 358.730 15.940 ;
        RECT 404.410 15.880 404.730 15.940 ;
        RECT 358.410 15.740 404.730 15.880 ;
        RECT 358.410 15.680 358.730 15.740 ;
        RECT 404.410 15.680 404.730 15.740 ;
      LAYER via ;
        RECT 324.860 17.040 325.120 17.300 ;
        RECT 358.440 17.040 358.700 17.300 ;
        RECT 358.440 15.680 358.700 15.940 ;
        RECT 404.440 15.680 404.700 15.940 ;
      LAYER met2 ;
        RECT 324.290 400.250 324.570 404.000 ;
        RECT 324.290 400.110 325.060 400.250 ;
        RECT 324.290 400.000 324.570 400.110 ;
        RECT 324.920 17.330 325.060 400.110 ;
        RECT 324.860 17.010 325.120 17.330 ;
        RECT 358.440 17.010 358.700 17.330 ;
        RECT 358.500 15.970 358.640 17.010 ;
        RECT 358.440 15.650 358.700 15.970 ;
        RECT 404.440 15.650 404.700 15.970 ;
        RECT 404.500 2.400 404.640 15.650 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.170 390.900 62.490 390.960 ;
        RECT 220.410 390.900 220.730 390.960 ;
        RECT 62.170 390.760 220.730 390.900 ;
        RECT 62.170 390.700 62.490 390.760 ;
        RECT 220.410 390.700 220.730 390.760 ;
      LAYER via ;
        RECT 62.200 390.700 62.460 390.960 ;
        RECT 220.440 390.700 220.700 390.960 ;
      LAYER met2 ;
        RECT 220.330 400.180 220.610 404.000 ;
        RECT 220.330 400.000 220.640 400.180 ;
        RECT 220.500 390.990 220.640 400.000 ;
        RECT 62.200 390.670 62.460 390.990 ;
        RECT 220.440 390.670 220.700 390.990 ;
        RECT 62.260 82.870 62.400 390.670 ;
        RECT 62.260 82.730 67.920 82.870 ;
        RECT 67.780 2.400 67.920 82.730 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 329.890 392.600 330.210 392.660 ;
        RECT 378.650 392.600 378.970 392.660 ;
        RECT 329.890 392.460 378.970 392.600 ;
        RECT 329.890 392.400 330.210 392.460 ;
        RECT 378.650 392.400 378.970 392.460 ;
        RECT 378.650 386.820 378.970 386.880 ;
        RECT 417.290 386.820 417.610 386.880 ;
        RECT 378.650 386.680 417.610 386.820 ;
        RECT 378.650 386.620 378.970 386.680 ;
        RECT 417.290 386.620 417.610 386.680 ;
        RECT 417.290 20.640 417.610 20.700 ;
        RECT 420.970 20.640 421.290 20.700 ;
        RECT 417.290 20.500 421.290 20.640 ;
        RECT 417.290 20.440 417.610 20.500 ;
        RECT 420.970 20.440 421.290 20.500 ;
      LAYER via ;
        RECT 329.920 392.400 330.180 392.660 ;
        RECT 378.680 392.400 378.940 392.660 ;
        RECT 378.680 386.620 378.940 386.880 ;
        RECT 417.320 386.620 417.580 386.880 ;
        RECT 417.320 20.440 417.580 20.700 ;
        RECT 421.000 20.440 421.260 20.700 ;
      LAYER met2 ;
        RECT 329.810 400.180 330.090 404.000 ;
        RECT 329.810 400.000 330.120 400.180 ;
        RECT 329.980 392.690 330.120 400.000 ;
        RECT 329.920 392.370 330.180 392.690 ;
        RECT 378.680 392.370 378.940 392.690 ;
        RECT 378.740 386.910 378.880 392.370 ;
        RECT 378.680 386.590 378.940 386.910 ;
        RECT 417.320 386.590 417.580 386.910 ;
        RECT 417.380 20.730 417.520 386.590 ;
        RECT 417.320 20.410 417.580 20.730 ;
        RECT 421.000 20.410 421.260 20.730 ;
        RECT 421.060 1.770 421.200 20.410 ;
        RECT 422.230 1.770 422.790 2.400 ;
        RECT 421.060 1.630 422.790 1.770 ;
        RECT 422.230 -4.800 422.790 1.630 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 335.410 393.280 335.730 393.340 ;
        RECT 335.410 393.140 379.340 393.280 ;
        RECT 335.410 393.080 335.730 393.140 ;
        RECT 379.200 392.940 379.340 393.140 ;
        RECT 424.190 392.940 424.510 393.000 ;
        RECT 379.200 392.800 424.510 392.940 ;
        RECT 424.190 392.740 424.510 392.800 ;
        RECT 424.190 16.900 424.510 16.960 ;
        RECT 439.830 16.900 440.150 16.960 ;
        RECT 424.190 16.760 440.150 16.900 ;
        RECT 424.190 16.700 424.510 16.760 ;
        RECT 439.830 16.700 440.150 16.760 ;
      LAYER via ;
        RECT 335.440 393.080 335.700 393.340 ;
        RECT 424.220 392.740 424.480 393.000 ;
        RECT 424.220 16.700 424.480 16.960 ;
        RECT 439.860 16.700 440.120 16.960 ;
      LAYER met2 ;
        RECT 335.330 400.180 335.610 404.000 ;
        RECT 335.330 400.000 335.640 400.180 ;
        RECT 335.500 393.370 335.640 400.000 ;
        RECT 335.440 393.050 335.700 393.370 ;
        RECT 424.220 392.710 424.480 393.030 ;
        RECT 424.280 16.990 424.420 392.710 ;
        RECT 424.220 16.670 424.480 16.990 ;
        RECT 439.860 16.670 440.120 16.990 ;
        RECT 439.920 2.400 440.060 16.670 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 339.550 24.720 339.870 24.780 ;
        RECT 457.770 24.720 458.090 24.780 ;
        RECT 339.550 24.580 458.090 24.720 ;
        RECT 339.550 24.520 339.870 24.580 ;
        RECT 457.770 24.520 458.090 24.580 ;
      LAYER via ;
        RECT 339.580 24.520 339.840 24.780 ;
        RECT 457.800 24.520 458.060 24.780 ;
      LAYER met2 ;
        RECT 340.850 400.250 341.130 404.000 ;
        RECT 339.640 400.110 341.130 400.250 ;
        RECT 339.640 24.810 339.780 400.110 ;
        RECT 340.850 400.000 341.130 400.110 ;
        RECT 339.580 24.490 339.840 24.810 ;
        RECT 457.800 24.490 458.060 24.810 ;
        RECT 457.860 2.400 458.000 24.490 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 397.050 391.920 397.370 391.980 ;
        RECT 465.590 391.920 465.910 391.980 ;
        RECT 397.050 391.780 465.910 391.920 ;
        RECT 397.050 391.720 397.370 391.780 ;
        RECT 465.590 391.720 465.910 391.780 ;
        RECT 345.990 389.540 346.310 389.600 ;
        RECT 397.050 389.540 397.370 389.600 ;
        RECT 345.990 389.400 397.370 389.540 ;
        RECT 345.990 389.340 346.310 389.400 ;
        RECT 397.050 389.340 397.370 389.400 ;
        RECT 465.590 20.300 465.910 20.360 ;
        RECT 475.710 20.300 476.030 20.360 ;
        RECT 465.590 20.160 476.030 20.300 ;
        RECT 465.590 20.100 465.910 20.160 ;
        RECT 475.710 20.100 476.030 20.160 ;
      LAYER via ;
        RECT 397.080 391.720 397.340 391.980 ;
        RECT 465.620 391.720 465.880 391.980 ;
        RECT 346.020 389.340 346.280 389.600 ;
        RECT 397.080 389.340 397.340 389.600 ;
        RECT 465.620 20.100 465.880 20.360 ;
        RECT 475.740 20.100 476.000 20.360 ;
      LAYER met2 ;
        RECT 345.910 400.180 346.190 404.000 ;
        RECT 345.910 400.000 346.220 400.180 ;
        RECT 346.080 389.630 346.220 400.000 ;
        RECT 397.080 391.690 397.340 392.010 ;
        RECT 465.620 391.690 465.880 392.010 ;
        RECT 397.140 389.630 397.280 391.690 ;
        RECT 346.020 389.310 346.280 389.630 ;
        RECT 397.080 389.310 397.340 389.630 ;
        RECT 465.680 20.390 465.820 391.690 ;
        RECT 465.620 20.070 465.880 20.390 ;
        RECT 475.740 20.070 476.000 20.390 ;
        RECT 475.800 2.400 475.940 20.070 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 376.280 345.390 376.340 ;
        RECT 350.130 376.280 350.450 376.340 ;
        RECT 345.070 376.140 350.450 376.280 ;
        RECT 345.070 376.080 345.390 376.140 ;
        RECT 350.130 376.080 350.450 376.140 ;
        RECT 397.050 19.960 397.370 20.020 ;
        RECT 493.190 19.960 493.510 20.020 ;
        RECT 397.050 19.820 493.510 19.960 ;
        RECT 397.050 19.760 397.370 19.820 ;
        RECT 493.190 19.760 493.510 19.820 ;
        RECT 345.070 18.600 345.390 18.660 ;
        RECT 397.050 18.600 397.370 18.660 ;
        RECT 345.070 18.460 397.370 18.600 ;
        RECT 345.070 18.400 345.390 18.460 ;
        RECT 397.050 18.400 397.370 18.460 ;
      LAYER via ;
        RECT 345.100 376.080 345.360 376.340 ;
        RECT 350.160 376.080 350.420 376.340 ;
        RECT 397.080 19.760 397.340 20.020 ;
        RECT 493.220 19.760 493.480 20.020 ;
        RECT 345.100 18.400 345.360 18.660 ;
        RECT 397.080 18.400 397.340 18.660 ;
      LAYER met2 ;
        RECT 351.430 400.250 351.710 404.000 ;
        RECT 350.220 400.110 351.710 400.250 ;
        RECT 350.220 376.370 350.360 400.110 ;
        RECT 351.430 400.000 351.710 400.110 ;
        RECT 345.100 376.050 345.360 376.370 ;
        RECT 350.160 376.050 350.420 376.370 ;
        RECT 345.160 18.690 345.300 376.050 ;
        RECT 397.080 19.730 397.340 20.050 ;
        RECT 493.220 19.730 493.480 20.050 ;
        RECT 397.140 18.690 397.280 19.730 ;
        RECT 345.100 18.370 345.360 18.690 ;
        RECT 397.080 18.370 397.340 18.690 ;
        RECT 493.280 2.400 493.420 19.730 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.090 391.580 500.410 391.640 ;
        RECT 479.940 391.440 500.410 391.580 ;
        RECT 357.030 390.900 357.350 390.960 ;
        RECT 479.940 390.900 480.080 391.440 ;
        RECT 500.090 391.380 500.410 391.440 ;
        RECT 357.030 390.760 480.080 390.900 ;
        RECT 357.030 390.700 357.350 390.760 ;
        RECT 500.090 17.240 500.410 17.300 ;
        RECT 511.130 17.240 511.450 17.300 ;
        RECT 500.090 17.100 511.450 17.240 ;
        RECT 500.090 17.040 500.410 17.100 ;
        RECT 511.130 17.040 511.450 17.100 ;
      LAYER via ;
        RECT 357.060 390.700 357.320 390.960 ;
        RECT 500.120 391.380 500.380 391.640 ;
        RECT 500.120 17.040 500.380 17.300 ;
        RECT 511.160 17.040 511.420 17.300 ;
      LAYER met2 ;
        RECT 356.950 400.180 357.230 404.000 ;
        RECT 356.950 400.000 357.260 400.180 ;
        RECT 357.120 390.990 357.260 400.000 ;
        RECT 500.120 391.350 500.380 391.670 ;
        RECT 357.060 390.670 357.320 390.990 ;
        RECT 500.180 17.330 500.320 391.350 ;
        RECT 500.120 17.010 500.380 17.330 ;
        RECT 511.160 17.010 511.420 17.330 ;
        RECT 511.220 2.400 511.360 17.010 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.330 19.280 359.650 19.340 ;
        RECT 528.610 19.280 528.930 19.340 ;
        RECT 359.330 19.140 528.930 19.280 ;
        RECT 359.330 19.080 359.650 19.140 ;
        RECT 528.610 19.080 528.930 19.140 ;
      LAYER via ;
        RECT 359.360 19.080 359.620 19.340 ;
        RECT 528.640 19.080 528.900 19.340 ;
      LAYER met2 ;
        RECT 362.470 400.250 362.750 404.000 ;
        RECT 361.260 400.110 362.750 400.250 ;
        RECT 361.260 324.370 361.400 400.110 ;
        RECT 362.470 400.000 362.750 400.110 ;
        RECT 359.420 324.230 361.400 324.370 ;
        RECT 359.420 19.370 359.560 324.230 ;
        RECT 359.360 19.050 359.620 19.370 ;
        RECT 528.640 19.050 528.900 19.370 ;
        RECT 528.700 2.400 528.840 19.050 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 368.070 388.860 368.390 388.920 ;
        RECT 506.530 388.860 506.850 388.920 ;
        RECT 368.070 388.720 506.850 388.860 ;
        RECT 368.070 388.660 368.390 388.720 ;
        RECT 506.530 388.660 506.850 388.720 ;
        RECT 507.450 20.300 507.770 20.360 ;
        RECT 546.550 20.300 546.870 20.360 ;
        RECT 507.450 20.160 546.870 20.300 ;
        RECT 507.450 20.100 507.770 20.160 ;
        RECT 546.550 20.100 546.870 20.160 ;
      LAYER via ;
        RECT 368.100 388.660 368.360 388.920 ;
        RECT 506.560 388.660 506.820 388.920 ;
        RECT 507.480 20.100 507.740 20.360 ;
        RECT 546.580 20.100 546.840 20.360 ;
      LAYER met2 ;
        RECT 367.990 400.180 368.270 404.000 ;
        RECT 367.990 400.000 368.300 400.180 ;
        RECT 368.160 388.950 368.300 400.000 ;
        RECT 368.100 388.630 368.360 388.950 ;
        RECT 506.560 388.630 506.820 388.950 ;
        RECT 506.620 372.670 506.760 388.630 ;
        RECT 506.620 372.530 507.220 372.670 ;
        RECT 507.080 82.870 507.220 372.530 ;
        RECT 507.080 82.730 507.680 82.870 ;
        RECT 507.540 20.390 507.680 82.730 ;
        RECT 507.480 20.070 507.740 20.390 ;
        RECT 546.580 20.070 546.840 20.390 ;
        RECT 546.640 2.400 546.780 20.070 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 373.130 24.040 373.450 24.100 ;
        RECT 503.770 24.040 504.090 24.100 ;
        RECT 373.130 23.900 504.090 24.040 ;
        RECT 373.130 23.840 373.450 23.900 ;
        RECT 503.770 23.840 504.090 23.900 ;
        RECT 503.770 15.540 504.090 15.600 ;
        RECT 564.030 15.540 564.350 15.600 ;
        RECT 503.770 15.400 564.350 15.540 ;
        RECT 503.770 15.340 504.090 15.400 ;
        RECT 564.030 15.340 564.350 15.400 ;
      LAYER via ;
        RECT 373.160 23.840 373.420 24.100 ;
        RECT 503.800 23.840 504.060 24.100 ;
        RECT 503.800 15.340 504.060 15.600 ;
        RECT 564.060 15.340 564.320 15.600 ;
      LAYER met2 ;
        RECT 373.510 400.250 373.790 404.000 ;
        RECT 373.220 400.110 373.790 400.250 ;
        RECT 373.220 24.130 373.360 400.110 ;
        RECT 373.510 400.000 373.790 400.110 ;
        RECT 373.160 23.810 373.420 24.130 ;
        RECT 503.800 23.810 504.060 24.130 ;
        RECT 503.860 15.630 504.000 23.810 ;
        RECT 503.800 15.310 504.060 15.630 ;
        RECT 564.060 15.310 564.320 15.630 ;
        RECT 564.120 2.400 564.260 15.310 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.110 392.600 379.430 392.660 ;
        RECT 424.650 392.600 424.970 392.660 ;
        RECT 379.110 392.460 424.970 392.600 ;
        RECT 379.110 392.400 379.430 392.460 ;
        RECT 424.650 392.400 424.970 392.460 ;
        RECT 424.650 388.520 424.970 388.580 ;
        RECT 514.810 388.520 515.130 388.580 ;
        RECT 424.650 388.380 515.130 388.520 ;
        RECT 424.650 388.320 424.970 388.380 ;
        RECT 514.810 388.320 515.130 388.380 ;
        RECT 513.890 15.880 514.210 15.940 ;
        RECT 581.970 15.880 582.290 15.940 ;
        RECT 513.890 15.740 582.290 15.880 ;
        RECT 513.890 15.680 514.210 15.740 ;
        RECT 581.970 15.680 582.290 15.740 ;
      LAYER via ;
        RECT 379.140 392.400 379.400 392.660 ;
        RECT 424.680 392.400 424.940 392.660 ;
        RECT 424.680 388.320 424.940 388.580 ;
        RECT 514.840 388.320 515.100 388.580 ;
        RECT 513.920 15.680 514.180 15.940 ;
        RECT 582.000 15.680 582.260 15.940 ;
      LAYER met2 ;
        RECT 379.030 400.180 379.310 404.000 ;
        RECT 379.030 400.000 379.340 400.180 ;
        RECT 379.200 392.690 379.340 400.000 ;
        RECT 379.140 392.370 379.400 392.690 ;
        RECT 424.680 392.370 424.940 392.690 ;
        RECT 424.740 388.610 424.880 392.370 ;
        RECT 424.680 388.290 424.940 388.610 ;
        RECT 514.840 388.290 515.100 388.610 ;
        RECT 514.900 381.890 515.040 388.290 ;
        RECT 513.980 381.750 515.040 381.890 ;
        RECT 513.980 15.970 514.120 381.750 ;
        RECT 513.920 15.650 514.180 15.970 ;
        RECT 582.000 15.650 582.260 15.970 ;
        RECT 582.060 2.400 582.200 15.650 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 91.150 19.620 91.470 19.680 ;
        RECT 228.690 19.620 229.010 19.680 ;
        RECT 91.150 19.480 229.010 19.620 ;
        RECT 91.150 19.420 91.470 19.480 ;
        RECT 228.690 19.420 229.010 19.480 ;
      LAYER via ;
        RECT 91.180 19.420 91.440 19.680 ;
        RECT 228.720 19.420 228.980 19.680 ;
      LAYER met2 ;
        RECT 227.690 400.250 227.970 404.000 ;
        RECT 227.690 400.110 228.920 400.250 ;
        RECT 227.690 400.000 227.970 400.110 ;
        RECT 228.780 19.710 228.920 400.110 ;
        RECT 91.180 19.390 91.440 19.710 ;
        RECT 228.720 19.390 228.980 19.710 ;
        RECT 91.240 2.400 91.380 19.390 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.490 386.480 380.810 386.540 ;
        RECT 383.250 386.480 383.570 386.540 ;
        RECT 380.490 386.340 383.570 386.480 ;
        RECT 380.490 386.280 380.810 386.340 ;
        RECT 383.250 386.280 383.570 386.340 ;
        RECT 380.490 17.920 380.810 17.980 ;
        RECT 599.450 17.920 599.770 17.980 ;
        RECT 380.490 17.780 599.770 17.920 ;
        RECT 380.490 17.720 380.810 17.780 ;
        RECT 599.450 17.720 599.770 17.780 ;
      LAYER via ;
        RECT 380.520 386.280 380.780 386.540 ;
        RECT 383.280 386.280 383.540 386.540 ;
        RECT 380.520 17.720 380.780 17.980 ;
        RECT 599.480 17.720 599.740 17.980 ;
      LAYER met2 ;
        RECT 384.550 400.250 384.830 404.000 ;
        RECT 383.340 400.110 384.830 400.250 ;
        RECT 383.340 386.570 383.480 400.110 ;
        RECT 384.550 400.000 384.830 400.110 ;
        RECT 380.520 386.250 380.780 386.570 ;
        RECT 383.280 386.250 383.540 386.570 ;
        RECT 380.580 18.010 380.720 386.250 ;
        RECT 380.520 17.690 380.780 18.010 ;
        RECT 599.480 17.690 599.740 18.010 ;
        RECT 599.540 2.400 599.680 17.690 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 390.150 388.520 390.470 388.580 ;
        RECT 390.150 388.380 424.420 388.520 ;
        RECT 390.150 388.320 390.470 388.380 ;
        RECT 424.280 388.180 424.420 388.380 ;
        RECT 520.790 388.180 521.110 388.240 ;
        RECT 424.280 388.040 521.110 388.180 ;
        RECT 520.790 387.980 521.110 388.040 ;
        RECT 520.790 19.960 521.110 20.020 ;
        RECT 520.790 19.820 530.220 19.960 ;
        RECT 520.790 19.760 521.110 19.820 ;
        RECT 530.080 19.620 530.220 19.820 ;
        RECT 617.390 19.620 617.710 19.680 ;
        RECT 530.080 19.480 617.710 19.620 ;
        RECT 617.390 19.420 617.710 19.480 ;
      LAYER via ;
        RECT 390.180 388.320 390.440 388.580 ;
        RECT 520.820 387.980 521.080 388.240 ;
        RECT 520.820 19.760 521.080 20.020 ;
        RECT 617.420 19.420 617.680 19.680 ;
      LAYER met2 ;
        RECT 390.070 400.180 390.350 404.000 ;
        RECT 390.070 400.000 390.380 400.180 ;
        RECT 390.240 388.610 390.380 400.000 ;
        RECT 390.180 388.290 390.440 388.610 ;
        RECT 520.820 387.950 521.080 388.270 ;
        RECT 520.880 20.050 521.020 387.950 ;
        RECT 520.820 19.730 521.080 20.050 ;
        RECT 617.420 19.390 617.680 19.710 ;
        RECT 617.480 2.400 617.620 19.390 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 110.470 391.580 110.790 391.640 ;
        RECT 235.130 391.580 235.450 391.640 ;
        RECT 110.470 391.440 235.450 391.580 ;
        RECT 110.470 391.380 110.790 391.440 ;
        RECT 235.130 391.380 235.450 391.440 ;
      LAYER via ;
        RECT 110.500 391.380 110.760 391.640 ;
        RECT 235.160 391.380 235.420 391.640 ;
      LAYER met2 ;
        RECT 235.050 400.180 235.330 404.000 ;
        RECT 235.050 400.000 235.360 400.180 ;
        RECT 235.220 391.670 235.360 400.000 ;
        RECT 110.500 391.350 110.760 391.670 ;
        RECT 235.160 391.350 235.420 391.670 ;
        RECT 110.560 82.870 110.700 391.350 ;
        RECT 110.560 82.730 113.000 82.870 ;
        RECT 112.860 1.770 113.000 82.730 ;
        RECT 114.950 1.770 115.510 2.400 ;
        RECT 112.860 1.630 115.510 1.770 ;
        RECT 114.950 -4.800 115.510 1.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.530 16.900 138.850 16.960 ;
        RECT 242.030 16.900 242.350 16.960 ;
        RECT 138.530 16.760 242.350 16.900 ;
        RECT 138.530 16.700 138.850 16.760 ;
        RECT 242.030 16.700 242.350 16.760 ;
      LAYER via ;
        RECT 138.560 16.700 138.820 16.960 ;
        RECT 242.060 16.700 242.320 16.960 ;
      LAYER met2 ;
        RECT 242.410 400.250 242.690 404.000 ;
        RECT 242.120 400.110 242.690 400.250 ;
        RECT 242.120 16.990 242.260 400.110 ;
        RECT 242.410 400.000 242.690 400.110 ;
        RECT 138.560 16.670 138.820 16.990 ;
        RECT 242.060 16.670 242.320 16.990 ;
        RECT 138.620 2.400 138.760 16.670 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 151.870 392.940 152.190 393.000 ;
        RECT 248.010 392.940 248.330 393.000 ;
        RECT 151.870 392.800 248.330 392.940 ;
        RECT 151.870 392.740 152.190 392.800 ;
        RECT 248.010 392.740 248.330 392.800 ;
      LAYER via ;
        RECT 151.900 392.740 152.160 393.000 ;
        RECT 248.040 392.740 248.300 393.000 ;
      LAYER met2 ;
        RECT 247.930 400.180 248.210 404.000 ;
        RECT 247.930 400.000 248.240 400.180 ;
        RECT 248.100 393.030 248.240 400.000 ;
        RECT 151.900 392.710 152.160 393.030 ;
        RECT 248.040 392.710 248.300 393.030 ;
        RECT 151.960 82.870 152.100 392.710 ;
        RECT 151.960 82.730 154.400 82.870 ;
        RECT 154.260 1.770 154.400 82.730 ;
        RECT 156.350 1.770 156.910 2.400 ;
        RECT 154.260 1.630 156.910 1.770 ;
        RECT 156.350 -4.800 156.910 1.630 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 173.950 16.220 174.270 16.280 ;
        RECT 249.390 16.220 249.710 16.280 ;
        RECT 173.950 16.080 249.710 16.220 ;
        RECT 173.950 16.020 174.270 16.080 ;
        RECT 249.390 16.020 249.710 16.080 ;
      LAYER via ;
        RECT 173.980 16.020 174.240 16.280 ;
        RECT 249.420 16.020 249.680 16.280 ;
      LAYER met2 ;
        RECT 252.990 400.250 253.270 404.000 ;
        RECT 251.780 400.110 253.270 400.250 ;
        RECT 251.780 386.650 251.920 400.110 ;
        RECT 252.990 400.000 253.270 400.110 ;
        RECT 249.480 386.510 251.920 386.650 ;
        RECT 249.480 16.310 249.620 386.510 ;
        RECT 173.980 15.990 174.240 16.310 ;
        RECT 249.420 15.990 249.680 16.310 ;
        RECT 174.040 2.400 174.180 15.990 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 191.890 15.880 192.210 15.940 ;
        RECT 255.830 15.880 256.150 15.940 ;
        RECT 191.890 15.740 256.150 15.880 ;
        RECT 191.890 15.680 192.210 15.740 ;
        RECT 255.830 15.680 256.150 15.740 ;
      LAYER via ;
        RECT 191.920 15.680 192.180 15.940 ;
        RECT 255.860 15.680 256.120 15.940 ;
      LAYER met2 ;
        RECT 258.510 400.250 258.790 404.000 ;
        RECT 257.300 400.110 258.790 400.250 ;
        RECT 257.300 386.650 257.440 400.110 ;
        RECT 258.510 400.000 258.790 400.110 ;
        RECT 255.920 386.510 257.440 386.650 ;
        RECT 255.920 15.970 256.060 386.510 ;
        RECT 191.920 15.650 192.180 15.970 ;
        RECT 255.860 15.650 256.120 15.970 ;
        RECT 191.980 2.400 192.120 15.650 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 252.150 386.820 252.470 386.880 ;
        RECT 264.110 386.820 264.430 386.880 ;
        RECT 252.150 386.680 264.430 386.820 ;
        RECT 252.150 386.620 252.470 386.680 ;
        RECT 264.110 386.620 264.430 386.680 ;
        RECT 251.690 18.260 252.010 18.320 ;
        RECT 228.320 18.120 252.010 18.260 ;
        RECT 209.370 17.920 209.690 17.980 ;
        RECT 209.370 17.780 227.770 17.920 ;
        RECT 209.370 17.720 209.690 17.780 ;
        RECT 227.630 17.580 227.770 17.780 ;
        RECT 228.320 17.580 228.460 18.120 ;
        RECT 251.690 18.060 252.010 18.120 ;
        RECT 227.630 17.440 228.460 17.580 ;
      LAYER via ;
        RECT 252.180 386.620 252.440 386.880 ;
        RECT 264.140 386.620 264.400 386.880 ;
        RECT 209.400 17.720 209.660 17.980 ;
        RECT 251.720 18.060 251.980 18.320 ;
      LAYER met2 ;
        RECT 264.030 400.180 264.310 404.000 ;
        RECT 264.030 400.000 264.340 400.180 ;
        RECT 264.200 386.910 264.340 400.000 ;
        RECT 252.180 386.590 252.440 386.910 ;
        RECT 264.140 386.590 264.400 386.910 ;
        RECT 252.240 324.370 252.380 386.590 ;
        RECT 251.780 324.230 252.380 324.370 ;
        RECT 251.780 18.350 251.920 324.230 ;
        RECT 251.720 18.030 251.980 18.350 ;
        RECT 209.400 17.690 209.660 18.010 ;
        RECT 209.460 2.400 209.600 17.690 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.870 389.880 221.190 389.940 ;
        RECT 269.630 389.880 269.950 389.940 ;
        RECT 220.870 389.740 269.950 389.880 ;
        RECT 220.870 389.680 221.190 389.740 ;
        RECT 269.630 389.680 269.950 389.740 ;
      LAYER via ;
        RECT 220.900 389.680 221.160 389.940 ;
        RECT 269.660 389.680 269.920 389.940 ;
      LAYER met2 ;
        RECT 269.550 400.180 269.830 404.000 ;
        RECT 269.550 400.000 269.860 400.180 ;
        RECT 269.720 389.970 269.860 400.000 ;
        RECT 220.900 389.650 221.160 389.970 ;
        RECT 269.660 389.650 269.920 389.970 ;
        RECT 220.960 18.090 221.100 389.650 ;
        RECT 220.960 17.950 223.860 18.090 ;
        RECT 223.720 2.450 223.860 17.950 ;
        RECT 223.720 2.310 225.240 2.450 ;
        RECT 225.100 1.770 225.240 2.310 ;
        RECT 227.190 1.770 227.750 2.400 ;
        RECT 225.100 1.630 227.750 1.770 ;
        RECT 227.190 -4.800 227.750 1.630 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 48.370 390.220 48.690 390.280 ;
        RECT 214.890 390.220 215.210 390.280 ;
        RECT 48.370 390.080 215.210 390.220 ;
        RECT 48.370 390.020 48.690 390.080 ;
        RECT 214.890 390.020 215.210 390.080 ;
      LAYER via ;
        RECT 48.400 390.020 48.660 390.280 ;
        RECT 214.920 390.020 215.180 390.280 ;
      LAYER met2 ;
        RECT 214.810 400.180 215.090 404.000 ;
        RECT 214.810 400.000 215.120 400.180 ;
        RECT 214.980 390.310 215.120 400.000 ;
        RECT 48.400 389.990 48.660 390.310 ;
        RECT 214.920 389.990 215.180 390.310 ;
        RECT 48.460 1.770 48.600 389.990 ;
        RECT 49.630 1.770 50.190 2.400 ;
        RECT 48.460 1.630 50.190 1.770 ;
        RECT 49.630 -4.800 50.190 1.630 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.470 391.580 248.790 391.640 ;
        RECT 276.990 391.580 277.310 391.640 ;
        RECT 248.470 391.440 277.310 391.580 ;
        RECT 248.470 391.380 248.790 391.440 ;
        RECT 276.990 391.380 277.310 391.440 ;
      LAYER via ;
        RECT 248.500 391.380 248.760 391.640 ;
        RECT 277.020 391.380 277.280 391.640 ;
      LAYER met2 ;
        RECT 276.910 400.180 277.190 404.000 ;
        RECT 276.910 400.000 277.220 400.180 ;
        RECT 277.080 391.670 277.220 400.000 ;
        RECT 248.500 391.350 248.760 391.670 ;
        RECT 277.020 391.350 277.280 391.670 ;
        RECT 248.560 14.690 248.700 391.350 ;
        RECT 248.560 14.550 251.000 14.690 ;
        RECT 250.860 2.400 251.000 14.550 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 272.390 393.280 272.710 393.340 ;
        RECT 282.510 393.280 282.830 393.340 ;
        RECT 272.390 393.140 282.830 393.280 ;
        RECT 272.390 393.080 272.710 393.140 ;
        RECT 282.510 393.080 282.830 393.140 ;
        RECT 268.710 16.560 269.030 16.620 ;
        RECT 272.390 16.560 272.710 16.620 ;
        RECT 268.710 16.420 272.710 16.560 ;
        RECT 268.710 16.360 269.030 16.420 ;
        RECT 272.390 16.360 272.710 16.420 ;
      LAYER via ;
        RECT 272.420 393.080 272.680 393.340 ;
        RECT 282.540 393.080 282.800 393.340 ;
        RECT 268.740 16.360 269.000 16.620 ;
        RECT 272.420 16.360 272.680 16.620 ;
      LAYER met2 ;
        RECT 282.430 400.180 282.710 404.000 ;
        RECT 282.430 400.000 282.740 400.180 ;
        RECT 282.600 393.370 282.740 400.000 ;
        RECT 272.420 393.050 272.680 393.370 ;
        RECT 282.540 393.050 282.800 393.370 ;
        RECT 272.480 16.650 272.620 393.050 ;
        RECT 268.740 16.330 269.000 16.650 ;
        RECT 272.420 16.330 272.680 16.650 ;
        RECT 268.800 2.400 268.940 16.330 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.970 386.140 283.290 386.200 ;
        RECT 286.650 386.140 286.970 386.200 ;
        RECT 282.970 386.000 286.970 386.140 ;
        RECT 282.970 385.940 283.290 386.000 ;
        RECT 286.650 385.940 286.970 386.000 ;
        RECT 282.970 17.580 283.290 17.640 ;
        RECT 284.350 17.580 284.670 17.640 ;
        RECT 282.970 17.440 284.670 17.580 ;
        RECT 282.970 17.380 283.290 17.440 ;
        RECT 284.350 17.380 284.670 17.440 ;
      LAYER via ;
        RECT 283.000 385.940 283.260 386.200 ;
        RECT 286.680 385.940 286.940 386.200 ;
        RECT 283.000 17.380 283.260 17.640 ;
        RECT 284.380 17.380 284.640 17.640 ;
      LAYER met2 ;
        RECT 287.950 400.250 288.230 404.000 ;
        RECT 286.740 400.110 288.230 400.250 ;
        RECT 286.740 386.230 286.880 400.110 ;
        RECT 287.950 400.000 288.230 400.110 ;
        RECT 283.000 385.910 283.260 386.230 ;
        RECT 286.680 385.910 286.940 386.230 ;
        RECT 283.060 17.670 283.200 385.910 ;
        RECT 283.000 17.350 283.260 17.670 ;
        RECT 284.380 17.350 284.640 17.670 ;
        RECT 284.440 1.770 284.580 17.350 ;
        RECT 286.070 1.770 286.630 2.400 ;
        RECT 284.440 1.630 286.630 1.770 ;
        RECT 286.070 -4.800 286.630 1.630 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 291.250 18.260 291.570 18.320 ;
        RECT 304.130 18.260 304.450 18.320 ;
        RECT 291.250 18.120 304.450 18.260 ;
        RECT 291.250 18.060 291.570 18.120 ;
        RECT 304.130 18.060 304.450 18.120 ;
      LAYER via ;
        RECT 291.280 18.060 291.540 18.320 ;
        RECT 304.160 18.060 304.420 18.320 ;
      LAYER met2 ;
        RECT 293.470 400.250 293.750 404.000 ;
        RECT 292.260 400.110 293.750 400.250 ;
        RECT 292.260 324.370 292.400 400.110 ;
        RECT 293.470 400.000 293.750 400.110 ;
        RECT 291.340 324.230 292.400 324.370 ;
        RECT 291.340 18.350 291.480 324.230 ;
        RECT 291.280 18.030 291.540 18.350 ;
        RECT 304.160 18.030 304.420 18.350 ;
        RECT 304.220 2.400 304.360 18.030 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.610 386.820 298.930 386.880 ;
        RECT 317.470 386.820 317.790 386.880 ;
        RECT 298.610 386.680 317.790 386.820 ;
        RECT 298.610 386.620 298.930 386.680 ;
        RECT 317.470 386.620 317.790 386.680 ;
      LAYER via ;
        RECT 298.640 386.620 298.900 386.880 ;
        RECT 317.500 386.620 317.760 386.880 ;
      LAYER met2 ;
        RECT 298.530 400.180 298.810 404.000 ;
        RECT 298.530 400.000 298.840 400.180 ;
        RECT 298.700 386.910 298.840 400.000 ;
        RECT 298.640 386.590 298.900 386.910 ;
        RECT 317.500 386.590 317.760 386.910 ;
        RECT 317.560 17.410 317.700 386.590 ;
        RECT 317.560 17.270 321.840 17.410 ;
        RECT 321.700 2.400 321.840 17.270 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.670 19.620 303.990 19.680 ;
        RECT 303.670 19.480 320.000 19.620 ;
        RECT 303.670 19.420 303.990 19.480 ;
        RECT 319.860 18.600 320.000 19.480 ;
        RECT 339.550 18.600 339.870 18.660 ;
        RECT 319.860 18.460 339.870 18.600 ;
        RECT 339.550 18.400 339.870 18.460 ;
      LAYER via ;
        RECT 303.700 19.420 303.960 19.680 ;
        RECT 339.580 18.400 339.840 18.660 ;
      LAYER met2 ;
        RECT 304.050 400.250 304.330 404.000 ;
        RECT 303.760 400.110 304.330 400.250 ;
        RECT 303.760 19.710 303.900 400.110 ;
        RECT 304.050 400.000 304.330 400.110 ;
        RECT 303.700 19.390 303.960 19.710 ;
        RECT 339.580 18.370 339.840 18.690 ;
        RECT 339.640 2.400 339.780 18.370 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 309.650 389.540 309.970 389.600 ;
        RECT 341.390 389.540 341.710 389.600 ;
        RECT 309.650 389.400 341.710 389.540 ;
        RECT 309.650 389.340 309.970 389.400 ;
        RECT 341.390 389.340 341.710 389.400 ;
        RECT 341.390 16.220 341.710 16.280 ;
        RECT 357.490 16.220 357.810 16.280 ;
        RECT 341.390 16.080 357.810 16.220 ;
        RECT 341.390 16.020 341.710 16.080 ;
        RECT 357.490 16.020 357.810 16.080 ;
      LAYER via ;
        RECT 309.680 389.340 309.940 389.600 ;
        RECT 341.420 389.340 341.680 389.600 ;
        RECT 341.420 16.020 341.680 16.280 ;
        RECT 357.520 16.020 357.780 16.280 ;
      LAYER met2 ;
        RECT 309.570 400.180 309.850 404.000 ;
        RECT 309.570 400.000 309.880 400.180 ;
        RECT 309.740 389.630 309.880 400.000 ;
        RECT 309.680 389.310 309.940 389.630 ;
        RECT 341.420 389.310 341.680 389.630 ;
        RECT 341.480 16.310 341.620 389.310 ;
        RECT 341.420 15.990 341.680 16.310 ;
        RECT 357.520 15.990 357.780 16.310 ;
        RECT 357.580 2.400 357.720 15.990 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 315.170 386.480 315.490 386.540 ;
        RECT 348.290 386.480 348.610 386.540 ;
        RECT 315.170 386.340 348.610 386.480 ;
        RECT 315.170 386.280 315.490 386.340 ;
        RECT 348.290 386.280 348.610 386.340 ;
        RECT 348.290 20.300 348.610 20.360 ;
        RECT 374.970 20.300 375.290 20.360 ;
        RECT 348.290 20.160 375.290 20.300 ;
        RECT 348.290 20.100 348.610 20.160 ;
        RECT 374.970 20.100 375.290 20.160 ;
      LAYER via ;
        RECT 315.200 386.280 315.460 386.540 ;
        RECT 348.320 386.280 348.580 386.540 ;
        RECT 348.320 20.100 348.580 20.360 ;
        RECT 375.000 20.100 375.260 20.360 ;
      LAYER met2 ;
        RECT 315.090 400.180 315.370 404.000 ;
        RECT 315.090 400.000 315.400 400.180 ;
        RECT 315.260 386.570 315.400 400.000 ;
        RECT 315.200 386.250 315.460 386.570 ;
        RECT 348.320 386.250 348.580 386.570 ;
        RECT 348.380 20.390 348.520 386.250 ;
        RECT 348.320 20.070 348.580 20.390 ;
        RECT 375.000 20.070 375.260 20.390 ;
        RECT 375.060 2.400 375.200 20.070 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.930 376.280 318.250 376.340 ;
        RECT 319.310 376.280 319.630 376.340 ;
        RECT 317.930 376.140 319.630 376.280 ;
        RECT 317.930 376.080 318.250 376.140 ;
        RECT 319.310 376.080 319.630 376.140 ;
        RECT 317.930 17.720 318.250 17.980 ;
        RECT 318.020 16.560 318.160 17.720 ;
        RECT 392.910 16.560 393.230 16.620 ;
        RECT 318.020 16.420 393.230 16.560 ;
        RECT 392.910 16.360 393.230 16.420 ;
      LAYER via ;
        RECT 317.960 376.080 318.220 376.340 ;
        RECT 319.340 376.080 319.600 376.340 ;
        RECT 317.960 17.720 318.220 17.980 ;
        RECT 392.940 16.360 393.200 16.620 ;
      LAYER met2 ;
        RECT 320.610 400.250 320.890 404.000 ;
        RECT 319.400 400.110 320.890 400.250 ;
        RECT 319.400 376.370 319.540 400.110 ;
        RECT 320.610 400.000 320.890 400.110 ;
        RECT 317.960 376.050 318.220 376.370 ;
        RECT 319.340 376.050 319.600 376.370 ;
        RECT 318.020 18.010 318.160 376.050 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 392.940 16.330 393.200 16.650 ;
        RECT 393.000 2.400 393.140 16.330 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 376.280 324.690 376.340 ;
        RECT 325.290 376.280 325.610 376.340 ;
        RECT 324.370 376.140 325.610 376.280 ;
        RECT 324.370 376.080 324.690 376.140 ;
        RECT 325.290 376.080 325.610 376.140 ;
        RECT 324.370 20.640 324.690 20.700 ;
        RECT 410.390 20.640 410.710 20.700 ;
        RECT 324.370 20.500 410.710 20.640 ;
        RECT 324.370 20.440 324.690 20.500 ;
        RECT 410.390 20.440 410.710 20.500 ;
      LAYER via ;
        RECT 324.400 376.080 324.660 376.340 ;
        RECT 325.320 376.080 325.580 376.340 ;
        RECT 324.400 20.440 324.660 20.700 ;
        RECT 410.420 20.440 410.680 20.700 ;
      LAYER met2 ;
        RECT 326.130 400.250 326.410 404.000 ;
        RECT 325.380 400.110 326.410 400.250 ;
        RECT 325.380 376.370 325.520 400.110 ;
        RECT 326.130 400.000 326.410 400.110 ;
        RECT 324.400 376.050 324.660 376.370 ;
        RECT 325.320 376.050 325.580 376.370 ;
        RECT 324.460 20.730 324.600 376.050 ;
        RECT 324.400 20.410 324.660 20.730 ;
        RECT 410.420 20.410 410.680 20.730 ;
        RECT 410.480 2.400 410.620 20.410 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 69.070 390.560 69.390 390.620 ;
        RECT 220.870 390.560 221.190 390.620 ;
        RECT 69.070 390.420 221.190 390.560 ;
        RECT 69.070 390.360 69.390 390.420 ;
        RECT 220.870 390.360 221.190 390.420 ;
      LAYER via ;
        RECT 69.100 390.360 69.360 390.620 ;
        RECT 220.900 390.360 221.160 390.620 ;
      LAYER met2 ;
        RECT 222.170 400.250 222.450 404.000 ;
        RECT 220.960 400.110 222.450 400.250 ;
        RECT 220.960 390.650 221.100 400.110 ;
        RECT 222.170 400.000 222.450 400.110 ;
        RECT 69.100 390.330 69.360 390.650 ;
        RECT 220.900 390.330 221.160 390.650 ;
        RECT 69.160 82.870 69.300 390.330 ;
        RECT 69.160 82.730 71.600 82.870 ;
        RECT 71.460 1.770 71.600 82.730 ;
        RECT 73.550 1.770 74.110 2.400 ;
        RECT 71.460 1.630 74.110 1.770 ;
        RECT 73.550 -4.800 74.110 1.630 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.330 16.220 428.650 16.280 ;
        RECT 358.040 16.080 428.650 16.220 ;
        RECT 331.270 15.880 331.590 15.940 ;
        RECT 358.040 15.880 358.180 16.080 ;
        RECT 428.330 16.020 428.650 16.080 ;
        RECT 331.270 15.740 358.180 15.880 ;
        RECT 331.270 15.680 331.590 15.740 ;
      LAYER via ;
        RECT 331.300 15.680 331.560 15.940 ;
        RECT 428.360 16.020 428.620 16.280 ;
      LAYER met2 ;
        RECT 331.650 400.250 331.930 404.000 ;
        RECT 331.360 400.110 331.930 400.250 ;
        RECT 331.360 15.970 331.500 400.110 ;
        RECT 331.650 400.000 331.930 400.110 ;
        RECT 428.360 15.990 428.620 16.310 ;
        RECT 331.300 15.650 331.560 15.970 ;
        RECT 428.420 2.400 428.560 15.990 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.730 376.280 332.050 376.340 ;
        RECT 335.870 376.280 336.190 376.340 ;
        RECT 331.730 376.140 336.190 376.280 ;
        RECT 331.730 376.080 332.050 376.140 ;
        RECT 335.870 376.080 336.190 376.140 ;
        RECT 331.730 15.200 332.050 15.260 ;
        RECT 445.810 15.200 446.130 15.260 ;
        RECT 331.730 15.060 446.130 15.200 ;
        RECT 331.730 15.000 332.050 15.060 ;
        RECT 445.810 15.000 446.130 15.060 ;
      LAYER via ;
        RECT 331.760 376.080 332.020 376.340 ;
        RECT 335.900 376.080 336.160 376.340 ;
        RECT 331.760 15.000 332.020 15.260 ;
        RECT 445.840 15.000 446.100 15.260 ;
      LAYER met2 ;
        RECT 337.170 400.250 337.450 404.000 ;
        RECT 335.960 400.110 337.450 400.250 ;
        RECT 335.960 376.370 336.100 400.110 ;
        RECT 337.170 400.000 337.450 400.110 ;
        RECT 331.760 376.050 332.020 376.370 ;
        RECT 335.900 376.050 336.160 376.370 ;
        RECT 331.820 15.290 331.960 376.050 ;
        RECT 331.760 14.970 332.020 15.290 ;
        RECT 445.840 14.970 446.100 15.290 ;
        RECT 445.900 2.400 446.040 14.970 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 338.170 392.260 338.490 392.320 ;
        RECT 341.390 392.260 341.710 392.320 ;
        RECT 338.170 392.120 341.710 392.260 ;
        RECT 338.170 392.060 338.490 392.120 ;
        RECT 341.390 392.060 341.710 392.120 ;
        RECT 338.170 16.900 338.490 16.960 ;
        RECT 423.730 16.900 424.050 16.960 ;
        RECT 338.170 16.760 424.050 16.900 ;
        RECT 338.170 16.700 338.490 16.760 ;
        RECT 423.730 16.700 424.050 16.760 ;
        RECT 423.730 15.540 424.050 15.600 ;
        RECT 463.750 15.540 464.070 15.600 ;
        RECT 423.730 15.400 464.070 15.540 ;
        RECT 423.730 15.340 424.050 15.400 ;
        RECT 463.750 15.340 464.070 15.400 ;
      LAYER via ;
        RECT 338.200 392.060 338.460 392.320 ;
        RECT 341.420 392.060 341.680 392.320 ;
        RECT 338.200 16.700 338.460 16.960 ;
        RECT 423.760 16.700 424.020 16.960 ;
        RECT 423.760 15.340 424.020 15.600 ;
        RECT 463.780 15.340 464.040 15.600 ;
      LAYER met2 ;
        RECT 342.690 400.250 342.970 404.000 ;
        RECT 341.480 400.110 342.970 400.250 ;
        RECT 341.480 392.350 341.620 400.110 ;
        RECT 342.690 400.000 342.970 400.110 ;
        RECT 338.200 392.030 338.460 392.350 ;
        RECT 341.420 392.030 341.680 392.350 ;
        RECT 338.260 16.990 338.400 392.030 ;
        RECT 338.200 16.670 338.460 16.990 ;
        RECT 423.760 16.670 424.020 16.990 ;
        RECT 423.820 15.630 423.960 16.670 ;
        RECT 423.760 15.310 424.020 15.630 ;
        RECT 463.780 15.310 464.040 15.630 ;
        RECT 463.840 2.400 463.980 15.310 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.350 20.300 445.670 20.360 ;
        RECT 396.680 20.160 445.670 20.300 ;
        RECT 345.530 19.960 345.850 20.020 ;
        RECT 396.680 19.960 396.820 20.160 ;
        RECT 445.350 20.100 445.670 20.160 ;
        RECT 345.530 19.820 396.820 19.960 ;
        RECT 345.530 19.760 345.850 19.820 ;
        RECT 445.350 17.240 445.670 17.300 ;
        RECT 481.230 17.240 481.550 17.300 ;
        RECT 445.350 17.100 481.550 17.240 ;
        RECT 445.350 17.040 445.670 17.100 ;
        RECT 481.230 17.040 481.550 17.100 ;
      LAYER via ;
        RECT 345.560 19.760 345.820 20.020 ;
        RECT 445.380 20.100 445.640 20.360 ;
        RECT 445.380 17.040 445.640 17.300 ;
        RECT 481.260 17.040 481.520 17.300 ;
      LAYER met2 ;
        RECT 347.750 400.250 348.030 404.000 ;
        RECT 346.540 400.110 348.030 400.250 ;
        RECT 346.540 324.370 346.680 400.110 ;
        RECT 347.750 400.000 348.030 400.110 ;
        RECT 345.620 324.230 346.680 324.370 ;
        RECT 345.620 20.050 345.760 324.230 ;
        RECT 445.380 20.070 445.640 20.390 ;
        RECT 345.560 19.730 345.820 20.050 ;
        RECT 445.440 17.330 445.580 20.070 ;
        RECT 445.380 17.010 445.640 17.330 ;
        RECT 481.260 17.010 481.520 17.330 ;
        RECT 481.320 2.400 481.460 17.010 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 466.050 392.260 466.370 392.320 ;
        RECT 396.680 392.120 466.370 392.260 ;
        RECT 353.350 391.920 353.670 391.980 ;
        RECT 396.680 391.920 396.820 392.120 ;
        RECT 466.050 392.060 466.370 392.120 ;
        RECT 353.350 391.780 396.820 391.920 ;
        RECT 353.350 391.720 353.670 391.780 ;
        RECT 466.050 15.540 466.370 15.600 ;
        RECT 499.170 15.540 499.490 15.600 ;
        RECT 466.050 15.400 499.490 15.540 ;
        RECT 466.050 15.340 466.370 15.400 ;
        RECT 499.170 15.340 499.490 15.400 ;
      LAYER via ;
        RECT 353.380 391.720 353.640 391.980 ;
        RECT 466.080 392.060 466.340 392.320 ;
        RECT 466.080 15.340 466.340 15.600 ;
        RECT 499.200 15.340 499.460 15.600 ;
      LAYER met2 ;
        RECT 353.270 400.180 353.550 404.000 ;
        RECT 353.270 400.000 353.580 400.180 ;
        RECT 353.440 392.010 353.580 400.000 ;
        RECT 466.080 392.030 466.340 392.350 ;
        RECT 353.380 391.690 353.640 392.010 ;
        RECT 466.140 15.630 466.280 392.030 ;
        RECT 466.080 15.310 466.340 15.630 ;
        RECT 499.200 15.310 499.460 15.630 ;
        RECT 499.260 2.400 499.400 15.310 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 19.620 359.190 19.680 ;
        RECT 516.650 19.620 516.970 19.680 ;
        RECT 358.870 19.480 516.970 19.620 ;
        RECT 358.870 19.420 359.190 19.480 ;
        RECT 516.650 19.420 516.970 19.480 ;
      LAYER via ;
        RECT 358.900 19.420 359.160 19.680 ;
        RECT 516.680 19.420 516.940 19.680 ;
      LAYER met2 ;
        RECT 358.790 400.180 359.070 404.000 ;
        RECT 358.790 400.000 359.100 400.180 ;
        RECT 358.960 19.710 359.100 400.000 ;
        RECT 358.900 19.390 359.160 19.710 ;
        RECT 516.680 19.390 516.940 19.710 ;
        RECT 516.740 2.400 516.880 19.390 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.390 389.880 364.710 389.940 ;
        RECT 364.390 389.740 400.270 389.880 ;
        RECT 364.390 389.680 364.710 389.740 ;
        RECT 400.130 389.540 400.270 389.740 ;
        RECT 517.570 389.540 517.890 389.600 ;
        RECT 400.130 389.400 517.890 389.540 ;
        RECT 517.570 389.340 517.890 389.400 ;
        RECT 517.570 388.860 517.890 388.920 ;
        RECT 521.250 388.860 521.570 388.920 ;
        RECT 517.570 388.720 521.570 388.860 ;
        RECT 517.570 388.660 517.890 388.720 ;
        RECT 521.250 388.660 521.570 388.720 ;
        RECT 521.250 15.200 521.570 15.260 ;
        RECT 534.590 15.200 534.910 15.260 ;
        RECT 521.250 15.060 534.910 15.200 ;
        RECT 521.250 15.000 521.570 15.060 ;
        RECT 534.590 15.000 534.910 15.060 ;
      LAYER via ;
        RECT 364.420 389.680 364.680 389.940 ;
        RECT 517.600 389.340 517.860 389.600 ;
        RECT 517.600 388.660 517.860 388.920 ;
        RECT 521.280 388.660 521.540 388.920 ;
        RECT 521.280 15.000 521.540 15.260 ;
        RECT 534.620 15.000 534.880 15.260 ;
      LAYER met2 ;
        RECT 364.310 400.180 364.590 404.000 ;
        RECT 364.310 400.000 364.620 400.180 ;
        RECT 364.480 389.970 364.620 400.000 ;
        RECT 364.420 389.650 364.680 389.970 ;
        RECT 517.600 389.310 517.860 389.630 ;
        RECT 517.660 388.950 517.800 389.310 ;
        RECT 517.600 388.630 517.860 388.950 ;
        RECT 521.280 388.630 521.540 388.950 ;
        RECT 521.340 15.290 521.480 388.630 ;
        RECT 521.280 14.970 521.540 15.290 ;
        RECT 534.620 14.970 534.880 15.290 ;
        RECT 534.680 2.400 534.820 14.970 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 369.910 391.580 370.230 391.640 ;
        RECT 449.030 391.580 449.350 391.640 ;
        RECT 369.910 391.440 449.350 391.580 ;
        RECT 369.910 391.380 370.230 391.440 ;
        RECT 449.030 391.380 449.350 391.440 ;
        RECT 449.490 389.880 449.810 389.940 ;
        RECT 515.270 389.880 515.590 389.940 ;
        RECT 449.490 389.740 515.590 389.880 ;
        RECT 449.490 389.680 449.810 389.740 ;
        RECT 515.270 389.680 515.590 389.740 ;
        RECT 514.350 15.200 514.670 15.260 ;
        RECT 514.350 15.060 521.020 15.200 ;
        RECT 514.350 15.000 514.670 15.060 ;
        RECT 520.880 14.860 521.020 15.060 ;
        RECT 552.530 14.860 552.850 14.920 ;
        RECT 520.880 14.720 552.850 14.860 ;
        RECT 552.530 14.660 552.850 14.720 ;
      LAYER via ;
        RECT 369.940 391.380 370.200 391.640 ;
        RECT 449.060 391.380 449.320 391.640 ;
        RECT 449.520 389.680 449.780 389.940 ;
        RECT 515.300 389.680 515.560 389.940 ;
        RECT 514.380 15.000 514.640 15.260 ;
        RECT 552.560 14.660 552.820 14.920 ;
      LAYER met2 ;
        RECT 369.830 400.180 370.110 404.000 ;
        RECT 369.830 400.000 370.140 400.180 ;
        RECT 370.000 391.670 370.140 400.000 ;
        RECT 369.940 391.350 370.200 391.670 ;
        RECT 449.060 391.410 449.320 391.670 ;
        RECT 449.060 391.350 449.720 391.410 ;
        RECT 449.120 391.270 449.720 391.350 ;
        RECT 449.580 389.970 449.720 391.270 ;
        RECT 449.520 389.650 449.780 389.970 ;
        RECT 515.300 389.650 515.560 389.970 ;
        RECT 515.360 324.370 515.500 389.650 ;
        RECT 514.440 324.230 515.500 324.370 ;
        RECT 514.440 15.290 514.580 324.230 ;
        RECT 514.380 14.970 514.640 15.290 ;
        RECT 552.560 14.630 552.820 14.950 ;
        RECT 552.620 2.400 552.760 14.630 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 375.430 390.560 375.750 390.620 ;
        RECT 449.030 390.560 449.350 390.620 ;
        RECT 375.430 390.420 449.350 390.560 ;
        RECT 375.430 390.360 375.750 390.420 ;
        RECT 449.030 390.360 449.350 390.420 ;
        RECT 449.030 387.160 449.350 387.220 ;
        RECT 449.030 387.020 527.920 387.160 ;
        RECT 449.030 386.960 449.350 387.020 ;
        RECT 527.780 386.200 527.920 387.020 ;
        RECT 527.690 385.940 528.010 386.200 ;
        RECT 527.690 19.620 528.010 19.680 ;
        RECT 527.690 19.480 529.300 19.620 ;
        RECT 527.690 19.420 528.010 19.480 ;
        RECT 529.160 19.280 529.300 19.480 ;
        RECT 570.010 19.280 570.330 19.340 ;
        RECT 529.160 19.140 570.330 19.280 ;
        RECT 570.010 19.080 570.330 19.140 ;
      LAYER via ;
        RECT 375.460 390.360 375.720 390.620 ;
        RECT 449.060 390.360 449.320 390.620 ;
        RECT 449.060 386.960 449.320 387.220 ;
        RECT 527.720 385.940 527.980 386.200 ;
        RECT 527.720 19.420 527.980 19.680 ;
        RECT 570.040 19.080 570.300 19.340 ;
      LAYER met2 ;
        RECT 375.350 400.180 375.630 404.000 ;
        RECT 375.350 400.000 375.660 400.180 ;
        RECT 375.520 390.650 375.660 400.000 ;
        RECT 375.460 390.330 375.720 390.650 ;
        RECT 449.060 390.330 449.320 390.650 ;
        RECT 449.120 387.250 449.260 390.330 ;
        RECT 449.060 386.930 449.320 387.250 ;
        RECT 527.720 385.910 527.980 386.230 ;
        RECT 527.780 19.710 527.920 385.910 ;
        RECT 527.720 19.390 527.980 19.710 ;
        RECT 570.040 19.050 570.300 19.370 ;
        RECT 570.100 2.400 570.240 19.050 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.030 18.260 380.350 18.320 ;
        RECT 587.950 18.260 588.270 18.320 ;
        RECT 380.030 18.120 588.270 18.260 ;
        RECT 380.030 18.060 380.350 18.120 ;
        RECT 587.950 18.060 588.270 18.120 ;
      LAYER via ;
        RECT 380.060 18.060 380.320 18.320 ;
        RECT 587.980 18.060 588.240 18.320 ;
      LAYER met2 ;
        RECT 380.870 400.250 381.150 404.000 ;
        RECT 380.120 400.110 381.150 400.250 ;
        RECT 380.120 18.350 380.260 400.110 ;
        RECT 380.870 400.000 381.150 400.110 ;
        RECT 380.060 18.030 380.320 18.350 ;
        RECT 587.980 18.030 588.240 18.350 ;
        RECT 588.040 2.400 588.180 18.030 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 227.770 386.140 228.090 386.200 ;
        RECT 229.150 386.140 229.470 386.200 ;
        RECT 227.770 386.000 229.470 386.140 ;
        RECT 227.770 385.940 228.090 386.000 ;
        RECT 229.150 385.940 229.470 386.000 ;
        RECT 97.130 20.640 97.450 20.700 ;
        RECT 227.770 20.640 228.090 20.700 ;
        RECT 97.130 20.500 228.090 20.640 ;
        RECT 97.130 20.440 97.450 20.500 ;
        RECT 227.770 20.440 228.090 20.500 ;
      LAYER via ;
        RECT 227.800 385.940 228.060 386.200 ;
        RECT 229.180 385.940 229.440 386.200 ;
        RECT 97.160 20.440 97.420 20.700 ;
        RECT 227.800 20.440 228.060 20.700 ;
      LAYER met2 ;
        RECT 229.530 400.250 229.810 404.000 ;
        RECT 229.240 400.110 229.810 400.250 ;
        RECT 229.240 386.230 229.380 400.110 ;
        RECT 229.530 400.000 229.810 400.110 ;
        RECT 227.800 385.910 228.060 386.230 ;
        RECT 229.180 385.910 229.440 386.230 ;
        RECT 227.860 20.730 228.000 385.910 ;
        RECT 97.160 20.410 97.420 20.730 ;
        RECT 227.800 20.410 228.060 20.730 ;
        RECT 97.220 2.400 97.360 20.410 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.470 17.580 386.790 17.640 ;
        RECT 605.430 17.580 605.750 17.640 ;
        RECT 386.470 17.440 605.750 17.580 ;
        RECT 386.470 17.380 386.790 17.440 ;
        RECT 605.430 17.380 605.750 17.440 ;
      LAYER via ;
        RECT 386.500 17.380 386.760 17.640 ;
        RECT 605.460 17.380 605.720 17.640 ;
      LAYER met2 ;
        RECT 386.390 400.180 386.670 404.000 ;
        RECT 386.390 400.000 386.700 400.180 ;
        RECT 386.560 17.670 386.700 400.000 ;
        RECT 386.500 17.350 386.760 17.670 ;
        RECT 605.460 17.350 605.720 17.670 ;
        RECT 605.520 2.400 605.660 17.350 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.050 16.900 535.370 16.960 ;
        RECT 623.370 16.900 623.690 16.960 ;
        RECT 535.050 16.760 623.690 16.900 ;
        RECT 535.050 16.700 535.370 16.760 ;
        RECT 623.370 16.700 623.690 16.760 ;
      LAYER via ;
        RECT 535.080 16.700 535.340 16.960 ;
        RECT 623.400 16.700 623.660 16.960 ;
      LAYER met2 ;
        RECT 391.450 400.180 391.730 404.000 ;
        RECT 391.450 400.000 391.760 400.180 ;
        RECT 391.620 389.485 391.760 400.000 ;
        RECT 391.550 389.115 391.830 389.485 ;
        RECT 534.610 389.115 534.890 389.485 ;
        RECT 534.680 82.870 534.820 389.115 ;
        RECT 534.680 82.730 535.280 82.870 ;
        RECT 535.140 16.990 535.280 82.730 ;
        RECT 535.080 16.670 535.340 16.990 ;
        RECT 623.400 16.670 623.660 16.990 ;
        RECT 623.460 2.400 623.600 16.670 ;
        RECT 623.250 -4.800 623.810 2.400 ;
      LAYER via2 ;
        RECT 391.550 389.160 391.830 389.440 ;
        RECT 534.610 389.160 534.890 389.440 ;
      LAYER met3 ;
        RECT 391.525 389.450 391.855 389.465 ;
        RECT 534.585 389.450 534.915 389.465 ;
        RECT 391.525 389.150 534.915 389.450 ;
        RECT 391.525 389.135 391.855 389.150 ;
        RECT 534.585 389.135 534.915 389.150 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 117.370 391.920 117.690 391.980 ;
        RECT 236.970 391.920 237.290 391.980 ;
        RECT 117.370 391.780 237.290 391.920 ;
        RECT 117.370 391.720 117.690 391.780 ;
        RECT 236.970 391.720 237.290 391.780 ;
      LAYER via ;
        RECT 117.400 391.720 117.660 391.980 ;
        RECT 237.000 391.720 237.260 391.980 ;
      LAYER met2 ;
        RECT 236.890 400.180 237.170 404.000 ;
        RECT 236.890 400.000 237.200 400.180 ;
        RECT 237.060 392.010 237.200 400.000 ;
        RECT 117.400 391.690 117.660 392.010 ;
        RECT 237.000 391.690 237.260 392.010 ;
        RECT 117.460 82.870 117.600 391.690 ;
        RECT 117.460 82.730 121.280 82.870 ;
        RECT 121.140 2.400 121.280 82.730 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 144.510 16.560 144.830 16.620 ;
        RECT 242.950 16.560 243.270 16.620 ;
        RECT 144.510 16.420 243.270 16.560 ;
        RECT 144.510 16.360 144.830 16.420 ;
        RECT 242.950 16.360 243.270 16.420 ;
      LAYER via ;
        RECT 144.540 16.360 144.800 16.620 ;
        RECT 242.980 16.360 243.240 16.620 ;
      LAYER met2 ;
        RECT 244.250 400.250 244.530 404.000 ;
        RECT 243.040 400.110 244.530 400.250 ;
        RECT 243.040 16.650 243.180 400.110 ;
        RECT 244.250 400.000 244.530 400.110 ;
        RECT 144.540 16.330 144.800 16.650 ;
        RECT 242.980 16.330 243.240 16.650 ;
        RECT 144.600 2.400 144.740 16.330 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.770 392.600 159.090 392.660 ;
        RECT 249.390 392.600 249.710 392.660 ;
        RECT 158.770 392.460 249.710 392.600 ;
        RECT 158.770 392.400 159.090 392.460 ;
        RECT 249.390 392.400 249.710 392.460 ;
      LAYER via ;
        RECT 158.800 392.400 159.060 392.660 ;
        RECT 249.420 392.400 249.680 392.660 ;
      LAYER met2 ;
        RECT 249.310 400.180 249.590 404.000 ;
        RECT 249.310 400.000 249.620 400.180 ;
        RECT 249.480 392.690 249.620 400.000 ;
        RECT 158.800 392.370 159.060 392.690 ;
        RECT 249.420 392.370 249.680 392.690 ;
        RECT 158.860 82.870 159.000 392.370 ;
        RECT 158.860 82.730 159.920 82.870 ;
        RECT 159.780 1.770 159.920 82.730 ;
        RECT 161.870 1.770 162.430 2.400 ;
        RECT 159.780 1.630 162.430 1.770 ;
        RECT 161.870 -4.800 162.430 1.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.930 386.480 249.250 386.540 ;
        RECT 253.530 386.480 253.850 386.540 ;
        RECT 248.930 386.340 253.850 386.480 ;
        RECT 248.930 386.280 249.250 386.340 ;
        RECT 253.530 386.280 253.850 386.340 ;
        RECT 179.930 15.540 180.250 15.600 ;
        RECT 248.930 15.540 249.250 15.600 ;
        RECT 179.930 15.400 249.250 15.540 ;
        RECT 179.930 15.340 180.250 15.400 ;
        RECT 248.930 15.340 249.250 15.400 ;
      LAYER via ;
        RECT 248.960 386.280 249.220 386.540 ;
        RECT 253.560 386.280 253.820 386.540 ;
        RECT 179.960 15.340 180.220 15.600 ;
        RECT 248.960 15.340 249.220 15.600 ;
      LAYER met2 ;
        RECT 254.830 400.250 255.110 404.000 ;
        RECT 253.620 400.110 255.110 400.250 ;
        RECT 253.620 386.570 253.760 400.110 ;
        RECT 254.830 400.000 255.110 400.110 ;
        RECT 248.960 386.250 249.220 386.570 ;
        RECT 253.560 386.250 253.820 386.570 ;
        RECT 249.020 15.630 249.160 386.250 ;
        RECT 179.960 15.310 180.220 15.630 ;
        RECT 248.960 15.310 249.220 15.630 ;
        RECT 180.020 2.400 180.160 15.310 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 193.270 388.860 193.590 388.920 ;
        RECT 260.430 388.860 260.750 388.920 ;
        RECT 193.270 388.720 260.750 388.860 ;
        RECT 193.270 388.660 193.590 388.720 ;
        RECT 260.430 388.660 260.750 388.720 ;
      LAYER via ;
        RECT 193.300 388.660 193.560 388.920 ;
        RECT 260.460 388.660 260.720 388.920 ;
      LAYER met2 ;
        RECT 260.350 400.180 260.630 404.000 ;
        RECT 260.350 400.000 260.660 400.180 ;
        RECT 260.520 388.950 260.660 400.000 ;
        RECT 193.300 388.630 193.560 388.950 ;
        RECT 260.460 388.630 260.720 388.950 ;
        RECT 193.360 82.870 193.500 388.630 ;
        RECT 193.360 82.730 195.800 82.870 ;
        RECT 195.660 1.770 195.800 82.730 ;
        RECT 197.750 1.770 198.310 2.400 ;
        RECT 195.660 1.630 198.310 1.770 ;
        RECT 197.750 -4.800 198.310 1.630 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 224.090 390.220 224.410 390.280 ;
        RECT 265.950 390.220 266.270 390.280 ;
        RECT 224.090 390.080 266.270 390.220 ;
        RECT 224.090 390.020 224.410 390.080 ;
        RECT 265.950 390.020 266.270 390.080 ;
        RECT 215.350 17.580 215.670 17.640 ;
        RECT 224.090 17.580 224.410 17.640 ;
        RECT 215.350 17.440 224.410 17.580 ;
        RECT 215.350 17.380 215.670 17.440 ;
        RECT 224.090 17.380 224.410 17.440 ;
      LAYER via ;
        RECT 224.120 390.020 224.380 390.280 ;
        RECT 265.980 390.020 266.240 390.280 ;
        RECT 215.380 17.380 215.640 17.640 ;
        RECT 224.120 17.380 224.380 17.640 ;
      LAYER met2 ;
        RECT 265.870 400.180 266.150 404.000 ;
        RECT 265.870 400.000 266.180 400.180 ;
        RECT 266.040 390.310 266.180 400.000 ;
        RECT 224.120 389.990 224.380 390.310 ;
        RECT 265.980 389.990 266.240 390.310 ;
        RECT 224.180 17.670 224.320 389.990 ;
        RECT 215.380 17.350 215.640 17.670 ;
        RECT 224.120 17.350 224.380 17.670 ;
        RECT 215.440 2.400 215.580 17.350 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 265.490 386.820 265.810 386.880 ;
        RECT 271.470 386.820 271.790 386.880 ;
        RECT 265.490 386.680 271.790 386.820 ;
        RECT 265.490 386.620 265.810 386.680 ;
        RECT 271.470 386.620 271.790 386.680 ;
        RECT 233.290 17.240 233.610 17.300 ;
        RECT 265.490 17.240 265.810 17.300 ;
        RECT 233.290 17.100 265.810 17.240 ;
        RECT 233.290 17.040 233.610 17.100 ;
        RECT 265.490 17.040 265.810 17.100 ;
      LAYER via ;
        RECT 265.520 386.620 265.780 386.880 ;
        RECT 271.500 386.620 271.760 386.880 ;
        RECT 233.320 17.040 233.580 17.300 ;
        RECT 265.520 17.040 265.780 17.300 ;
      LAYER met2 ;
        RECT 271.390 400.180 271.670 404.000 ;
        RECT 271.390 400.000 271.700 400.180 ;
        RECT 271.560 386.910 271.700 400.000 ;
        RECT 265.520 386.590 265.780 386.910 ;
        RECT 271.500 386.590 271.760 386.910 ;
        RECT 265.580 17.330 265.720 386.590 ;
        RECT 233.320 17.010 233.580 17.330 ;
        RECT 265.520 17.010 265.780 17.330 ;
        RECT 233.380 2.400 233.520 17.010 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 55.730 18.940 56.050 19.000 ;
        RECT 214.430 18.940 214.750 19.000 ;
        RECT 55.730 18.800 214.750 18.940 ;
        RECT 55.730 18.740 56.050 18.800 ;
        RECT 214.430 18.740 214.750 18.800 ;
      LAYER via ;
        RECT 55.760 18.740 56.020 19.000 ;
        RECT 214.460 18.740 214.720 19.000 ;
      LAYER met2 ;
        RECT 216.650 400.250 216.930 404.000 ;
        RECT 215.440 400.110 216.930 400.250 ;
        RECT 215.440 386.470 215.580 400.110 ;
        RECT 216.650 400.000 216.930 400.110 ;
        RECT 214.520 386.330 215.580 386.470 ;
        RECT 214.520 19.030 214.660 386.330 ;
        RECT 55.760 18.710 56.020 19.030 ;
        RECT 214.460 18.710 214.720 19.030 ;
        RECT 55.820 2.400 55.960 18.710 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 75.970 391.240 76.290 391.300 ;
        RECT 224.090 391.240 224.410 391.300 ;
        RECT 75.970 391.100 224.410 391.240 ;
        RECT 75.970 391.040 76.290 391.100 ;
        RECT 224.090 391.040 224.410 391.100 ;
      LAYER via ;
        RECT 76.000 391.040 76.260 391.300 ;
        RECT 224.120 391.040 224.380 391.300 ;
      LAYER met2 ;
        RECT 224.010 400.180 224.290 404.000 ;
        RECT 224.010 400.000 224.320 400.180 ;
        RECT 224.180 391.330 224.320 400.000 ;
        RECT 76.000 391.010 76.260 391.330 ;
        RECT 224.120 391.010 224.380 391.330 ;
        RECT 76.060 82.870 76.200 391.010 ;
        RECT 76.060 82.730 79.880 82.870 ;
        RECT 79.740 2.400 79.880 82.730 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.230 386.480 228.550 386.540 ;
        RECT 230.070 386.480 230.390 386.540 ;
        RECT 228.230 386.340 230.390 386.480 ;
        RECT 228.230 386.280 228.550 386.340 ;
        RECT 230.070 386.280 230.390 386.340 ;
        RECT 103.110 20.300 103.430 20.360 ;
        RECT 228.230 20.300 228.550 20.360 ;
        RECT 103.110 20.160 228.550 20.300 ;
        RECT 103.110 20.100 103.430 20.160 ;
        RECT 228.230 20.100 228.550 20.160 ;
      LAYER via ;
        RECT 228.260 386.280 228.520 386.540 ;
        RECT 230.100 386.280 230.360 386.540 ;
        RECT 103.140 20.100 103.400 20.360 ;
        RECT 228.260 20.100 228.520 20.360 ;
      LAYER met2 ;
        RECT 231.370 400.250 231.650 404.000 ;
        RECT 230.160 400.110 231.650 400.250 ;
        RECT 230.160 386.570 230.300 400.110 ;
        RECT 231.370 400.000 231.650 400.110 ;
        RECT 228.260 386.250 228.520 386.570 ;
        RECT 230.100 386.250 230.360 386.570 ;
        RECT 228.320 20.390 228.460 386.250 ;
        RECT 103.140 20.070 103.400 20.390 ;
        RECT 228.260 20.070 228.520 20.390 ;
        RECT 103.200 2.400 103.340 20.070 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.270 392.260 124.590 392.320 ;
        RECT 238.810 392.260 239.130 392.320 ;
        RECT 124.270 392.120 239.130 392.260 ;
        RECT 124.270 392.060 124.590 392.120 ;
        RECT 238.810 392.060 239.130 392.120 ;
      LAYER via ;
        RECT 124.300 392.060 124.560 392.320 ;
        RECT 238.840 392.060 239.100 392.320 ;
      LAYER met2 ;
        RECT 238.730 400.180 239.010 404.000 ;
        RECT 238.730 400.000 239.040 400.180 ;
        RECT 238.900 392.350 239.040 400.000 ;
        RECT 124.300 392.030 124.560 392.350 ;
        RECT 238.840 392.030 239.100 392.350 ;
        RECT 124.360 82.870 124.500 392.030 ;
        RECT 124.360 82.730 126.800 82.870 ;
        RECT 126.660 2.400 126.800 82.730 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 207.990 17.240 208.310 17.300 ;
        RECT 26.290 17.100 208.310 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 207.990 17.040 208.310 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 208.020 17.040 208.280 17.300 ;
      LAYER met2 ;
        RECT 207.450 400.250 207.730 404.000 ;
        RECT 207.450 400.110 208.220 400.250 ;
        RECT 207.450 400.000 207.730 400.110 ;
        RECT 208.080 17.330 208.220 400.110 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 208.020 17.010 208.280 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.670 389.880 27.990 389.940 ;
        RECT 209.370 389.880 209.690 389.940 ;
        RECT 27.670 389.740 209.690 389.880 ;
        RECT 27.670 389.680 27.990 389.740 ;
        RECT 209.370 389.680 209.690 389.740 ;
      LAYER via ;
        RECT 27.700 389.680 27.960 389.940 ;
        RECT 209.400 389.680 209.660 389.940 ;
      LAYER met2 ;
        RECT 209.290 400.180 209.570 404.000 ;
        RECT 209.290 400.000 209.600 400.180 ;
        RECT 209.460 389.970 209.600 400.000 ;
        RECT 27.700 389.650 27.960 389.970 ;
        RECT 209.400 389.650 209.660 389.970 ;
        RECT 27.760 82.870 27.900 389.650 ;
        RECT 27.760 82.730 30.200 82.870 ;
        RECT 30.060 1.770 30.200 82.730 ;
        RECT 32.150 1.770 32.710 2.400 ;
        RECT 30.060 1.630 32.710 1.770 ;
        RECT 32.150 -4.800 32.710 1.630 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 205.520 410.795 1094.240 987.605 ;
      LAYER met1 ;
        RECT 203.290 410.640 1094.240 993.600 ;
      LAYER met2 ;
        RECT 203.870 995.720 209.930 996.770 ;
        RECT 210.770 995.720 216.830 996.770 ;
        RECT 217.670 995.720 224.190 996.770 ;
        RECT 225.030 995.720 231.090 996.770 ;
        RECT 231.930 995.720 238.450 996.770 ;
        RECT 239.290 995.720 245.350 996.770 ;
        RECT 246.190 995.720 252.250 996.770 ;
        RECT 253.090 995.720 259.610 996.770 ;
        RECT 260.450 995.720 266.510 996.770 ;
        RECT 267.350 995.720 273.870 996.770 ;
        RECT 274.710 995.720 280.770 996.770 ;
        RECT 281.610 995.720 287.670 996.770 ;
        RECT 288.510 995.720 295.030 996.770 ;
        RECT 295.870 995.720 301.930 996.770 ;
        RECT 302.770 995.720 309.290 996.770 ;
        RECT 310.130 995.720 316.190 996.770 ;
        RECT 317.030 995.720 323.090 996.770 ;
        RECT 323.930 995.720 330.450 996.770 ;
        RECT 331.290 995.720 337.350 996.770 ;
        RECT 338.190 995.720 344.710 996.770 ;
        RECT 345.550 995.720 351.610 996.770 ;
        RECT 352.450 995.720 358.970 996.770 ;
        RECT 359.810 995.720 365.870 996.770 ;
        RECT 366.710 995.720 372.770 996.770 ;
        RECT 373.610 995.720 380.130 996.770 ;
        RECT 380.970 995.720 387.030 996.770 ;
        RECT 387.870 995.720 394.390 996.770 ;
        RECT 395.230 995.720 401.290 996.770 ;
        RECT 402.130 995.720 408.190 996.770 ;
        RECT 409.030 995.720 415.550 996.770 ;
        RECT 416.390 995.720 422.450 996.770 ;
        RECT 423.290 995.720 429.810 996.770 ;
        RECT 430.650 995.720 436.710 996.770 ;
        RECT 437.550 995.720 443.610 996.770 ;
        RECT 444.450 995.720 450.970 996.770 ;
        RECT 451.810 995.720 457.870 996.770 ;
        RECT 458.710 995.720 465.230 996.770 ;
        RECT 466.070 995.720 472.130 996.770 ;
        RECT 472.970 995.720 479.030 996.770 ;
        RECT 479.870 995.720 486.390 996.770 ;
        RECT 487.230 995.720 493.290 996.770 ;
        RECT 494.130 995.720 500.650 996.770 ;
        RECT 501.490 995.720 507.550 996.770 ;
        RECT 508.390 995.720 514.910 996.770 ;
        RECT 515.750 995.720 521.810 996.770 ;
        RECT 522.650 995.720 528.710 996.770 ;
        RECT 529.550 995.720 536.070 996.770 ;
        RECT 536.910 995.720 542.970 996.770 ;
        RECT 543.810 995.720 550.330 996.770 ;
        RECT 551.170 995.720 557.230 996.770 ;
        RECT 558.070 995.720 564.130 996.770 ;
        RECT 564.970 995.720 571.490 996.770 ;
        RECT 572.330 995.720 578.390 996.770 ;
        RECT 579.230 995.720 585.750 996.770 ;
        RECT 586.590 995.720 592.650 996.770 ;
        RECT 593.490 995.720 599.550 996.770 ;
        RECT 600.390 995.720 606.910 996.770 ;
        RECT 607.750 995.720 613.810 996.770 ;
        RECT 614.650 995.720 621.170 996.770 ;
        RECT 622.010 995.720 628.070 996.770 ;
        RECT 628.910 995.720 634.970 996.770 ;
        RECT 635.810 995.720 642.330 996.770 ;
        RECT 643.170 995.720 649.230 996.770 ;
        RECT 650.070 995.720 656.590 996.770 ;
        RECT 657.430 995.720 663.490 996.770 ;
        RECT 664.330 995.720 670.850 996.770 ;
        RECT 671.690 995.720 677.750 996.770 ;
        RECT 678.590 995.720 684.650 996.770 ;
        RECT 685.490 995.720 692.010 996.770 ;
        RECT 692.850 995.720 698.910 996.770 ;
        RECT 699.750 995.720 706.270 996.770 ;
        RECT 707.110 995.720 713.170 996.770 ;
        RECT 714.010 995.720 720.070 996.770 ;
        RECT 720.910 995.720 727.430 996.770 ;
        RECT 728.270 995.720 734.330 996.770 ;
        RECT 735.170 995.720 741.690 996.770 ;
        RECT 742.530 995.720 748.590 996.770 ;
        RECT 749.430 995.720 755.490 996.770 ;
        RECT 756.330 995.720 762.850 996.770 ;
        RECT 763.690 995.720 769.750 996.770 ;
        RECT 770.590 995.720 777.110 996.770 ;
        RECT 777.950 995.720 784.010 996.770 ;
        RECT 784.850 995.720 790.910 996.770 ;
        RECT 791.750 995.720 798.270 996.770 ;
        RECT 799.110 995.720 805.170 996.770 ;
        RECT 806.010 995.720 812.530 996.770 ;
        RECT 813.370 995.720 819.430 996.770 ;
        RECT 820.270 995.720 826.790 996.770 ;
        RECT 827.630 995.720 833.690 996.770 ;
        RECT 834.530 995.720 840.590 996.770 ;
        RECT 841.430 995.720 847.950 996.770 ;
        RECT 848.790 995.720 854.850 996.770 ;
        RECT 855.690 995.720 862.210 996.770 ;
        RECT 863.050 995.720 869.110 996.770 ;
        RECT 869.950 995.720 876.010 996.770 ;
        RECT 876.850 995.720 883.370 996.770 ;
        RECT 884.210 995.720 890.270 996.770 ;
        RECT 891.110 995.720 897.630 996.770 ;
        RECT 898.470 995.720 904.530 996.770 ;
        RECT 905.370 995.720 911.430 996.770 ;
        RECT 912.270 995.720 918.790 996.770 ;
        RECT 919.630 995.720 925.690 996.770 ;
        RECT 926.530 995.720 933.050 996.770 ;
        RECT 933.890 995.720 939.950 996.770 ;
        RECT 940.790 995.720 946.850 996.770 ;
        RECT 947.690 995.720 954.210 996.770 ;
        RECT 955.050 995.720 961.110 996.770 ;
        RECT 961.950 995.720 968.470 996.770 ;
        RECT 969.310 995.720 975.370 996.770 ;
        RECT 976.210 995.720 982.730 996.770 ;
        RECT 983.570 995.720 989.630 996.770 ;
        RECT 990.470 995.720 996.530 996.770 ;
        RECT 997.370 995.720 1003.890 996.770 ;
        RECT 1004.730 995.720 1010.790 996.770 ;
        RECT 1011.630 995.720 1018.150 996.770 ;
        RECT 1018.990 995.720 1025.050 996.770 ;
        RECT 1025.890 995.720 1031.950 996.770 ;
        RECT 1032.790 995.720 1039.310 996.770 ;
        RECT 1040.150 995.720 1046.210 996.770 ;
        RECT 1047.050 995.720 1053.570 996.770 ;
        RECT 1054.410 995.720 1060.470 996.770 ;
        RECT 1061.310 995.720 1067.370 996.770 ;
        RECT 1068.210 995.720 1074.730 996.770 ;
        RECT 1075.570 995.720 1081.630 996.770 ;
        RECT 1082.470 995.720 1088.990 996.770 ;
        RECT 1089.830 995.720 1090.930 996.770 ;
        RECT 203.320 404.280 1090.930 995.720 ;
      LAYER met2 ;
        RECT 200.550 400.000 200.830 404.000 ;
      LAYER met2 ;
        RECT 203.320 403.670 203.490 404.280 ;
        RECT 204.330 403.670 205.330 404.280 ;
        RECT 206.170 403.670 207.170 404.280 ;
        RECT 208.010 403.670 209.010 404.280 ;
        RECT 209.850 403.670 210.850 404.280 ;
        RECT 211.690 403.670 212.690 404.280 ;
        RECT 213.530 403.670 214.530 404.280 ;
        RECT 215.370 403.670 216.370 404.280 ;
        RECT 217.210 403.670 218.210 404.280 ;
        RECT 219.050 403.670 220.050 404.280 ;
        RECT 220.890 403.670 221.890 404.280 ;
        RECT 222.730 403.670 223.730 404.280 ;
        RECT 224.570 403.670 225.570 404.280 ;
        RECT 226.410 403.670 227.410 404.280 ;
        RECT 228.250 403.670 229.250 404.280 ;
        RECT 230.090 403.670 231.090 404.280 ;
        RECT 231.930 403.670 232.930 404.280 ;
        RECT 233.770 403.670 234.770 404.280 ;
        RECT 235.610 403.670 236.610 404.280 ;
        RECT 237.450 403.670 238.450 404.280 ;
        RECT 239.290 403.670 240.290 404.280 ;
        RECT 241.130 403.670 242.130 404.280 ;
        RECT 242.970 403.670 243.970 404.280 ;
        RECT 244.810 403.670 245.810 404.280 ;
        RECT 246.650 403.670 247.650 404.280 ;
        RECT 248.490 403.670 249.030 404.280 ;
        RECT 249.870 403.670 250.870 404.280 ;
        RECT 251.710 403.670 252.710 404.280 ;
        RECT 253.550 403.670 254.550 404.280 ;
        RECT 255.390 403.670 256.390 404.280 ;
        RECT 257.230 403.670 258.230 404.280 ;
        RECT 259.070 403.670 260.070 404.280 ;
        RECT 260.910 403.670 261.910 404.280 ;
        RECT 262.750 403.670 263.750 404.280 ;
        RECT 264.590 403.670 265.590 404.280 ;
        RECT 266.430 403.670 267.430 404.280 ;
        RECT 268.270 403.670 269.270 404.280 ;
        RECT 270.110 403.670 271.110 404.280 ;
        RECT 271.950 403.670 272.950 404.280 ;
        RECT 273.790 403.670 274.790 404.280 ;
        RECT 275.630 403.670 276.630 404.280 ;
        RECT 277.470 403.670 278.470 404.280 ;
        RECT 279.310 403.670 280.310 404.280 ;
        RECT 281.150 403.670 282.150 404.280 ;
        RECT 282.990 403.670 283.990 404.280 ;
        RECT 284.830 403.670 285.830 404.280 ;
        RECT 286.670 403.670 287.670 404.280 ;
        RECT 288.510 403.670 289.510 404.280 ;
        RECT 290.350 403.670 291.350 404.280 ;
        RECT 292.190 403.670 293.190 404.280 ;
        RECT 294.030 403.670 295.030 404.280 ;
        RECT 295.870 403.670 296.410 404.280 ;
        RECT 297.250 403.670 298.250 404.280 ;
        RECT 299.090 403.670 300.090 404.280 ;
        RECT 300.930 403.670 301.930 404.280 ;
        RECT 302.770 403.670 303.770 404.280 ;
        RECT 304.610 403.670 305.610 404.280 ;
        RECT 306.450 403.670 307.450 404.280 ;
        RECT 308.290 403.670 309.290 404.280 ;
        RECT 310.130 403.670 311.130 404.280 ;
        RECT 311.970 403.670 312.970 404.280 ;
        RECT 313.810 403.670 314.810 404.280 ;
        RECT 315.650 403.670 316.650 404.280 ;
        RECT 317.490 403.670 318.490 404.280 ;
        RECT 319.330 403.670 320.330 404.280 ;
        RECT 321.170 403.670 322.170 404.280 ;
        RECT 323.010 403.670 324.010 404.280 ;
        RECT 324.850 403.670 325.850 404.280 ;
        RECT 326.690 403.670 327.690 404.280 ;
        RECT 328.530 403.670 329.530 404.280 ;
        RECT 330.370 403.670 331.370 404.280 ;
        RECT 332.210 403.670 333.210 404.280 ;
        RECT 334.050 403.670 335.050 404.280 ;
        RECT 335.890 403.670 336.890 404.280 ;
        RECT 337.730 403.670 338.730 404.280 ;
        RECT 339.570 403.670 340.570 404.280 ;
        RECT 341.410 403.670 342.410 404.280 ;
        RECT 343.250 403.670 343.790 404.280 ;
        RECT 344.630 403.670 345.630 404.280 ;
        RECT 346.470 403.670 347.470 404.280 ;
        RECT 348.310 403.670 349.310 404.280 ;
        RECT 350.150 403.670 351.150 404.280 ;
        RECT 351.990 403.670 352.990 404.280 ;
        RECT 353.830 403.670 354.830 404.280 ;
        RECT 355.670 403.670 356.670 404.280 ;
        RECT 357.510 403.670 358.510 404.280 ;
        RECT 359.350 403.670 360.350 404.280 ;
        RECT 361.190 403.670 362.190 404.280 ;
        RECT 363.030 403.670 364.030 404.280 ;
        RECT 364.870 403.670 365.870 404.280 ;
        RECT 366.710 403.670 367.710 404.280 ;
        RECT 368.550 403.670 369.550 404.280 ;
        RECT 370.390 403.670 371.390 404.280 ;
        RECT 372.230 403.670 373.230 404.280 ;
        RECT 374.070 403.670 375.070 404.280 ;
        RECT 375.910 403.670 376.910 404.280 ;
        RECT 377.750 403.670 378.750 404.280 ;
        RECT 379.590 403.670 380.590 404.280 ;
        RECT 381.430 403.670 382.430 404.280 ;
        RECT 383.270 403.670 384.270 404.280 ;
        RECT 385.110 403.670 386.110 404.280 ;
        RECT 386.950 403.670 387.950 404.280 ;
        RECT 388.790 403.670 389.790 404.280 ;
        RECT 390.630 403.670 391.170 404.280 ;
        RECT 392.010 403.670 393.010 404.280 ;
        RECT 393.850 403.670 394.850 404.280 ;
        RECT 395.690 403.670 396.690 404.280 ;
        RECT 397.530 403.670 398.530 404.280 ;
        RECT 399.370 403.670 400.370 404.280 ;
        RECT 401.210 403.670 402.210 404.280 ;
        RECT 403.050 403.670 404.050 404.280 ;
        RECT 404.890 403.670 405.890 404.280 ;
        RECT 406.730 403.670 407.730 404.280 ;
        RECT 408.570 403.670 409.570 404.280 ;
        RECT 410.410 403.670 411.410 404.280 ;
        RECT 412.250 403.670 413.250 404.280 ;
        RECT 414.090 403.670 415.090 404.280 ;
        RECT 415.930 403.670 416.930 404.280 ;
        RECT 417.770 403.670 418.770 404.280 ;
        RECT 419.610 403.670 420.610 404.280 ;
        RECT 421.450 403.670 422.450 404.280 ;
        RECT 423.290 403.670 424.290 404.280 ;
        RECT 425.130 403.670 426.130 404.280 ;
        RECT 426.970 403.670 427.970 404.280 ;
        RECT 428.810 403.670 429.810 404.280 ;
        RECT 430.650 403.670 431.650 404.280 ;
        RECT 432.490 403.670 433.490 404.280 ;
        RECT 434.330 403.670 435.330 404.280 ;
        RECT 436.170 403.670 437.170 404.280 ;
        RECT 438.010 403.670 438.550 404.280 ;
        RECT 439.390 403.670 440.390 404.280 ;
        RECT 441.230 403.670 442.230 404.280 ;
        RECT 443.070 403.670 444.070 404.280 ;
        RECT 444.910 403.670 445.910 404.280 ;
        RECT 446.750 403.670 447.750 404.280 ;
        RECT 448.590 403.670 449.590 404.280 ;
        RECT 450.430 403.670 451.430 404.280 ;
        RECT 452.270 403.670 453.270 404.280 ;
        RECT 454.110 403.670 455.110 404.280 ;
        RECT 455.950 403.670 456.950 404.280 ;
        RECT 457.790 403.670 458.790 404.280 ;
        RECT 459.630 403.670 460.630 404.280 ;
        RECT 461.470 403.670 462.470 404.280 ;
        RECT 463.310 403.670 464.310 404.280 ;
        RECT 465.150 403.670 466.150 404.280 ;
        RECT 466.990 403.670 467.990 404.280 ;
        RECT 468.830 403.670 469.830 404.280 ;
        RECT 470.670 403.670 471.670 404.280 ;
        RECT 472.510 403.670 473.510 404.280 ;
        RECT 474.350 403.670 475.350 404.280 ;
        RECT 476.190 403.670 477.190 404.280 ;
        RECT 478.030 403.670 479.030 404.280 ;
        RECT 479.870 403.670 480.870 404.280 ;
        RECT 481.710 403.670 482.710 404.280 ;
        RECT 483.550 403.670 484.550 404.280 ;
        RECT 485.390 403.670 485.930 404.280 ;
        RECT 486.770 403.670 487.770 404.280 ;
        RECT 488.610 403.670 489.610 404.280 ;
        RECT 490.450 403.670 491.450 404.280 ;
        RECT 492.290 403.670 493.290 404.280 ;
        RECT 494.130 403.670 495.130 404.280 ;
        RECT 495.970 403.670 496.970 404.280 ;
        RECT 497.810 403.670 498.810 404.280 ;
        RECT 499.650 403.670 500.650 404.280 ;
        RECT 501.490 403.670 502.490 404.280 ;
        RECT 503.330 403.670 504.330 404.280 ;
        RECT 505.170 403.670 506.170 404.280 ;
        RECT 507.010 403.670 508.010 404.280 ;
        RECT 508.850 403.670 509.850 404.280 ;
        RECT 510.690 403.670 511.690 404.280 ;
        RECT 512.530 403.670 513.530 404.280 ;
        RECT 514.370 403.670 515.370 404.280 ;
        RECT 516.210 403.670 517.210 404.280 ;
        RECT 518.050 403.670 519.050 404.280 ;
        RECT 519.890 403.670 520.890 404.280 ;
        RECT 521.730 403.670 522.730 404.280 ;
        RECT 523.570 403.670 524.570 404.280 ;
        RECT 525.410 403.670 526.410 404.280 ;
        RECT 527.250 403.670 528.250 404.280 ;
        RECT 529.090 403.670 530.090 404.280 ;
        RECT 530.930 403.670 531.930 404.280 ;
        RECT 532.770 403.670 533.310 404.280 ;
        RECT 534.150 403.670 535.150 404.280 ;
        RECT 535.990 403.670 536.990 404.280 ;
        RECT 537.830 403.670 538.830 404.280 ;
        RECT 539.670 403.670 540.670 404.280 ;
        RECT 541.510 403.670 542.510 404.280 ;
        RECT 543.350 403.670 544.350 404.280 ;
        RECT 545.190 403.670 546.190 404.280 ;
        RECT 547.030 403.670 548.030 404.280 ;
        RECT 548.870 403.670 549.870 404.280 ;
        RECT 550.710 403.670 551.710 404.280 ;
        RECT 552.550 403.670 553.550 404.280 ;
        RECT 554.390 403.670 555.390 404.280 ;
        RECT 556.230 403.670 557.230 404.280 ;
        RECT 558.070 403.670 559.070 404.280 ;
        RECT 559.910 403.670 560.910 404.280 ;
        RECT 561.750 403.670 562.750 404.280 ;
        RECT 563.590 403.670 564.590 404.280 ;
        RECT 565.430 403.670 566.430 404.280 ;
        RECT 567.270 403.670 568.270 404.280 ;
        RECT 569.110 403.670 570.110 404.280 ;
        RECT 570.950 403.670 571.950 404.280 ;
        RECT 572.790 403.670 573.790 404.280 ;
        RECT 574.630 403.670 575.630 404.280 ;
        RECT 576.470 403.670 577.470 404.280 ;
        RECT 578.310 403.670 579.310 404.280 ;
        RECT 580.150 403.670 580.690 404.280 ;
        RECT 581.530 403.670 582.530 404.280 ;
        RECT 583.370 403.670 584.370 404.280 ;
        RECT 585.210 403.670 586.210 404.280 ;
        RECT 587.050 403.670 588.050 404.280 ;
        RECT 588.890 403.670 589.890 404.280 ;
        RECT 590.730 403.670 591.730 404.280 ;
        RECT 592.570 403.670 593.570 404.280 ;
        RECT 594.410 403.670 595.410 404.280 ;
        RECT 596.250 403.670 597.250 404.280 ;
        RECT 598.090 403.670 599.090 404.280 ;
        RECT 599.930 403.670 600.930 404.280 ;
        RECT 601.770 403.670 602.770 404.280 ;
        RECT 603.610 403.670 604.610 404.280 ;
        RECT 605.450 403.670 606.450 404.280 ;
        RECT 607.290 403.670 608.290 404.280 ;
        RECT 609.130 403.670 610.130 404.280 ;
        RECT 610.970 403.670 611.970 404.280 ;
        RECT 612.810 403.670 613.810 404.280 ;
        RECT 614.650 403.670 615.650 404.280 ;
        RECT 616.490 403.670 617.490 404.280 ;
        RECT 618.330 403.670 619.330 404.280 ;
        RECT 620.170 403.670 621.170 404.280 ;
        RECT 622.010 403.670 623.010 404.280 ;
        RECT 623.850 403.670 624.850 404.280 ;
        RECT 625.690 403.670 626.690 404.280 ;
        RECT 627.530 403.670 628.070 404.280 ;
        RECT 628.910 403.670 629.910 404.280 ;
        RECT 630.750 403.670 631.750 404.280 ;
        RECT 632.590 403.670 633.590 404.280 ;
        RECT 634.430 403.670 635.430 404.280 ;
        RECT 636.270 403.670 637.270 404.280 ;
        RECT 638.110 403.670 639.110 404.280 ;
        RECT 639.950 403.670 640.950 404.280 ;
        RECT 641.790 403.670 642.790 404.280 ;
        RECT 643.630 403.670 644.630 404.280 ;
        RECT 645.470 403.670 646.470 404.280 ;
        RECT 647.310 403.670 648.310 404.280 ;
        RECT 649.150 403.670 650.150 404.280 ;
        RECT 650.990 403.670 651.990 404.280 ;
        RECT 652.830 403.670 653.830 404.280 ;
        RECT 654.670 403.670 655.670 404.280 ;
        RECT 656.510 403.670 657.510 404.280 ;
        RECT 658.350 403.670 659.350 404.280 ;
        RECT 660.190 403.670 661.190 404.280 ;
        RECT 662.030 403.670 663.030 404.280 ;
        RECT 663.870 403.670 664.870 404.280 ;
        RECT 665.710 403.670 666.710 404.280 ;
        RECT 667.550 403.670 668.550 404.280 ;
        RECT 669.390 403.670 670.390 404.280 ;
        RECT 671.230 403.670 672.230 404.280 ;
        RECT 673.070 403.670 674.070 404.280 ;
        RECT 674.910 403.670 675.450 404.280 ;
        RECT 676.290 403.670 677.290 404.280 ;
        RECT 678.130 403.670 679.130 404.280 ;
        RECT 679.970 403.670 680.970 404.280 ;
        RECT 681.810 403.670 682.810 404.280 ;
        RECT 683.650 403.670 684.650 404.280 ;
        RECT 685.490 403.670 686.490 404.280 ;
        RECT 687.330 403.670 688.330 404.280 ;
        RECT 689.170 403.670 690.170 404.280 ;
        RECT 691.010 403.670 692.010 404.280 ;
        RECT 692.850 403.670 693.850 404.280 ;
        RECT 694.690 403.670 695.690 404.280 ;
        RECT 696.530 403.670 697.530 404.280 ;
        RECT 698.370 403.670 699.370 404.280 ;
        RECT 700.210 403.670 701.210 404.280 ;
        RECT 702.050 403.670 703.050 404.280 ;
        RECT 703.890 403.670 704.890 404.280 ;
        RECT 705.730 403.670 706.730 404.280 ;
        RECT 707.570 403.670 708.570 404.280 ;
        RECT 709.410 403.670 710.410 404.280 ;
        RECT 711.250 403.670 712.250 404.280 ;
        RECT 713.090 403.670 714.090 404.280 ;
        RECT 714.930 403.670 715.930 404.280 ;
        RECT 716.770 403.670 717.770 404.280 ;
        RECT 718.610 403.670 719.610 404.280 ;
        RECT 720.450 403.670 721.450 404.280 ;
        RECT 722.290 403.670 722.830 404.280 ;
        RECT 723.670 403.670 724.670 404.280 ;
        RECT 725.510 403.670 726.510 404.280 ;
        RECT 727.350 403.670 728.350 404.280 ;
        RECT 729.190 403.670 730.190 404.280 ;
        RECT 731.030 403.670 732.030 404.280 ;
        RECT 732.870 403.670 733.870 404.280 ;
        RECT 734.710 403.670 735.710 404.280 ;
        RECT 736.550 403.670 737.550 404.280 ;
        RECT 738.390 403.670 739.390 404.280 ;
        RECT 740.230 403.670 741.230 404.280 ;
        RECT 742.070 403.670 743.070 404.280 ;
        RECT 743.910 403.670 744.910 404.280 ;
        RECT 745.750 403.670 746.750 404.280 ;
        RECT 747.590 403.670 748.590 404.280 ;
        RECT 749.430 403.670 750.430 404.280 ;
        RECT 751.270 403.670 752.270 404.280 ;
        RECT 753.110 403.670 754.110 404.280 ;
        RECT 754.950 403.670 755.950 404.280 ;
        RECT 756.790 403.670 757.790 404.280 ;
        RECT 758.630 403.670 759.630 404.280 ;
        RECT 760.470 403.670 761.470 404.280 ;
        RECT 762.310 403.670 763.310 404.280 ;
        RECT 764.150 403.670 765.150 404.280 ;
        RECT 765.990 403.670 766.990 404.280 ;
        RECT 767.830 403.670 768.830 404.280 ;
        RECT 769.670 403.670 770.210 404.280 ;
        RECT 771.050 403.670 772.050 404.280 ;
        RECT 772.890 403.670 773.890 404.280 ;
        RECT 774.730 403.670 775.730 404.280 ;
        RECT 776.570 403.670 777.570 404.280 ;
        RECT 778.410 403.670 779.410 404.280 ;
        RECT 780.250 403.670 781.250 404.280 ;
        RECT 782.090 403.670 783.090 404.280 ;
        RECT 783.930 403.670 784.930 404.280 ;
        RECT 785.770 403.670 786.770 404.280 ;
        RECT 787.610 403.670 788.610 404.280 ;
        RECT 789.450 403.670 790.450 404.280 ;
        RECT 791.290 403.670 792.290 404.280 ;
        RECT 793.130 403.670 794.130 404.280 ;
        RECT 794.970 403.670 795.970 404.280 ;
        RECT 796.810 403.670 797.810 404.280 ;
        RECT 798.650 403.670 799.650 404.280 ;
        RECT 800.490 403.670 801.490 404.280 ;
        RECT 802.330 403.670 803.330 404.280 ;
        RECT 804.170 403.670 805.170 404.280 ;
        RECT 806.010 403.670 807.010 404.280 ;
        RECT 807.850 403.670 808.850 404.280 ;
        RECT 809.690 403.670 810.690 404.280 ;
        RECT 811.530 403.670 812.530 404.280 ;
        RECT 813.370 403.670 814.370 404.280 ;
        RECT 815.210 403.670 816.210 404.280 ;
        RECT 817.050 403.670 817.590 404.280 ;
        RECT 818.430 403.670 819.430 404.280 ;
        RECT 820.270 403.670 821.270 404.280 ;
        RECT 822.110 403.670 823.110 404.280 ;
        RECT 823.950 403.670 824.950 404.280 ;
        RECT 825.790 403.670 826.790 404.280 ;
        RECT 827.630 403.670 828.630 404.280 ;
        RECT 829.470 403.670 830.470 404.280 ;
        RECT 831.310 403.670 832.310 404.280 ;
        RECT 833.150 403.670 834.150 404.280 ;
        RECT 834.990 403.670 835.990 404.280 ;
        RECT 836.830 403.670 837.830 404.280 ;
        RECT 838.670 403.670 839.670 404.280 ;
        RECT 840.510 403.670 841.510 404.280 ;
        RECT 842.350 403.670 843.350 404.280 ;
        RECT 844.190 403.670 845.190 404.280 ;
        RECT 846.030 403.670 847.030 404.280 ;
        RECT 847.870 403.670 848.870 404.280 ;
        RECT 849.710 403.670 850.710 404.280 ;
        RECT 851.550 403.670 852.550 404.280 ;
        RECT 853.390 403.670 854.390 404.280 ;
        RECT 855.230 403.670 856.230 404.280 ;
        RECT 857.070 403.670 858.070 404.280 ;
        RECT 858.910 403.670 859.910 404.280 ;
        RECT 860.750 403.670 861.750 404.280 ;
        RECT 862.590 403.670 863.590 404.280 ;
        RECT 864.430 403.670 864.970 404.280 ;
        RECT 865.810 403.670 866.810 404.280 ;
        RECT 867.650 403.670 868.650 404.280 ;
        RECT 869.490 403.670 870.490 404.280 ;
        RECT 871.330 403.670 872.330 404.280 ;
        RECT 873.170 403.670 874.170 404.280 ;
        RECT 875.010 403.670 876.010 404.280 ;
        RECT 876.850 403.670 877.850 404.280 ;
        RECT 878.690 403.670 879.690 404.280 ;
        RECT 880.530 403.670 881.530 404.280 ;
        RECT 882.370 403.670 883.370 404.280 ;
        RECT 884.210 403.670 885.210 404.280 ;
        RECT 886.050 403.670 887.050 404.280 ;
        RECT 887.890 403.670 888.890 404.280 ;
        RECT 889.730 403.670 890.730 404.280 ;
        RECT 891.570 403.670 892.570 404.280 ;
        RECT 893.410 403.670 894.410 404.280 ;
        RECT 895.250 403.670 896.250 404.280 ;
        RECT 897.090 403.670 898.090 404.280 ;
        RECT 898.930 403.670 899.930 404.280 ;
        RECT 900.770 403.670 901.770 404.280 ;
        RECT 902.610 403.670 903.610 404.280 ;
        RECT 904.450 403.670 905.450 404.280 ;
        RECT 906.290 403.670 907.290 404.280 ;
        RECT 908.130 403.670 909.130 404.280 ;
        RECT 909.970 403.670 910.970 404.280 ;
        RECT 911.810 403.670 912.350 404.280 ;
        RECT 913.190 403.670 914.190 404.280 ;
        RECT 915.030 403.670 916.030 404.280 ;
        RECT 916.870 403.670 917.870 404.280 ;
        RECT 918.710 403.670 919.710 404.280 ;
        RECT 920.550 403.670 921.550 404.280 ;
        RECT 922.390 403.670 923.390 404.280 ;
        RECT 924.230 403.670 925.230 404.280 ;
        RECT 926.070 403.670 927.070 404.280 ;
        RECT 927.910 403.670 928.910 404.280 ;
        RECT 929.750 403.670 930.750 404.280 ;
        RECT 931.590 403.670 932.590 404.280 ;
        RECT 933.430 403.670 934.430 404.280 ;
        RECT 935.270 403.670 936.270 404.280 ;
        RECT 937.110 403.670 938.110 404.280 ;
        RECT 938.950 403.670 939.950 404.280 ;
        RECT 940.790 403.670 941.790 404.280 ;
        RECT 942.630 403.670 943.630 404.280 ;
        RECT 944.470 403.670 945.470 404.280 ;
        RECT 946.310 403.670 947.310 404.280 ;
        RECT 948.150 403.670 949.150 404.280 ;
        RECT 949.990 403.670 950.990 404.280 ;
        RECT 951.830 403.670 952.830 404.280 ;
        RECT 953.670 403.670 954.670 404.280 ;
        RECT 955.510 403.670 956.510 404.280 ;
        RECT 957.350 403.670 958.350 404.280 ;
        RECT 959.190 403.670 959.730 404.280 ;
        RECT 960.570 403.670 961.570 404.280 ;
        RECT 962.410 403.670 963.410 404.280 ;
        RECT 964.250 403.670 965.250 404.280 ;
        RECT 966.090 403.670 967.090 404.280 ;
        RECT 967.930 403.670 968.930 404.280 ;
        RECT 969.770 403.670 970.770 404.280 ;
        RECT 971.610 403.670 972.610 404.280 ;
        RECT 973.450 403.670 974.450 404.280 ;
        RECT 975.290 403.670 976.290 404.280 ;
        RECT 977.130 403.670 978.130 404.280 ;
        RECT 978.970 403.670 979.970 404.280 ;
        RECT 980.810 403.670 981.810 404.280 ;
        RECT 982.650 403.670 983.650 404.280 ;
        RECT 984.490 403.670 985.490 404.280 ;
        RECT 986.330 403.670 987.330 404.280 ;
        RECT 988.170 403.670 989.170 404.280 ;
        RECT 990.010 403.670 991.010 404.280 ;
        RECT 991.850 403.670 992.850 404.280 ;
        RECT 993.690 403.670 994.690 404.280 ;
        RECT 995.530 403.670 996.530 404.280 ;
        RECT 997.370 403.670 998.370 404.280 ;
        RECT 999.210 403.670 1000.210 404.280 ;
        RECT 1001.050 403.670 1002.050 404.280 ;
        RECT 1002.890 403.670 1003.890 404.280 ;
        RECT 1004.730 403.670 1005.730 404.280 ;
        RECT 1006.570 403.670 1007.110 404.280 ;
        RECT 1007.950 403.670 1008.950 404.280 ;
        RECT 1009.790 403.670 1010.790 404.280 ;
        RECT 1011.630 403.670 1012.630 404.280 ;
        RECT 1013.470 403.670 1014.470 404.280 ;
        RECT 1015.310 403.670 1016.310 404.280 ;
        RECT 1017.150 403.670 1018.150 404.280 ;
        RECT 1018.990 403.670 1019.990 404.280 ;
        RECT 1020.830 403.670 1021.830 404.280 ;
        RECT 1022.670 403.670 1023.670 404.280 ;
        RECT 1024.510 403.670 1025.510 404.280 ;
        RECT 1026.350 403.670 1027.350 404.280 ;
        RECT 1028.190 403.670 1029.190 404.280 ;
        RECT 1030.030 403.670 1031.030 404.280 ;
        RECT 1031.870 403.670 1032.870 404.280 ;
        RECT 1033.710 403.670 1034.710 404.280 ;
        RECT 1035.550 403.670 1036.550 404.280 ;
        RECT 1037.390 403.670 1038.390 404.280 ;
        RECT 1039.230 403.670 1040.230 404.280 ;
        RECT 1041.070 403.670 1042.070 404.280 ;
        RECT 1042.910 403.670 1043.910 404.280 ;
        RECT 1044.750 403.670 1045.750 404.280 ;
        RECT 1046.590 403.670 1047.590 404.280 ;
        RECT 1048.430 403.670 1049.430 404.280 ;
        RECT 1050.270 403.670 1051.270 404.280 ;
        RECT 1052.110 403.670 1053.110 404.280 ;
        RECT 1053.950 403.670 1054.490 404.280 ;
        RECT 1055.330 403.670 1056.330 404.280 ;
        RECT 1057.170 403.670 1058.170 404.280 ;
        RECT 1059.010 403.670 1060.010 404.280 ;
        RECT 1060.850 403.670 1061.850 404.280 ;
        RECT 1062.690 403.670 1063.690 404.280 ;
        RECT 1064.530 403.670 1065.530 404.280 ;
        RECT 1066.370 403.670 1067.370 404.280 ;
        RECT 1068.210 403.670 1069.210 404.280 ;
        RECT 1070.050 403.670 1071.050 404.280 ;
        RECT 1071.890 403.670 1072.890 404.280 ;
        RECT 1073.730 403.670 1074.730 404.280 ;
        RECT 1075.570 403.670 1076.570 404.280 ;
        RECT 1077.410 403.670 1078.410 404.280 ;
        RECT 1079.250 403.670 1080.250 404.280 ;
        RECT 1081.090 403.670 1082.090 404.280 ;
        RECT 1082.930 403.670 1083.930 404.280 ;
        RECT 1084.770 403.670 1085.770 404.280 ;
        RECT 1086.610 403.670 1087.610 404.280 ;
        RECT 1088.450 403.670 1089.450 404.280 ;
        RECT 1090.290 403.670 1090.930 404.280 ;
      LAYER met3 ;
        RECT 204.000 970.200 1096.000 988.705 ;
        RECT 204.000 968.800 1095.600 970.200 ;
        RECT 204.000 957.960 1096.000 968.800 ;
        RECT 204.400 956.560 1096.000 957.960 ;
        RECT 204.000 910.360 1096.000 956.560 ;
        RECT 204.000 908.960 1095.600 910.360 ;
        RECT 204.000 872.280 1096.000 908.960 ;
        RECT 204.400 870.880 1096.000 872.280 ;
        RECT 204.000 850.520 1096.000 870.880 ;
        RECT 204.000 849.120 1095.600 850.520 ;
        RECT 204.000 790.680 1096.000 849.120 ;
        RECT 204.000 789.280 1095.600 790.680 ;
        RECT 204.000 786.600 1096.000 789.280 ;
        RECT 204.400 785.200 1096.000 786.600 ;
        RECT 204.000 730.840 1096.000 785.200 ;
        RECT 204.000 729.440 1095.600 730.840 ;
        RECT 204.000 700.920 1096.000 729.440 ;
        RECT 204.400 699.520 1096.000 700.920 ;
        RECT 204.000 670.320 1096.000 699.520 ;
        RECT 204.000 668.920 1095.600 670.320 ;
        RECT 204.000 615.240 1096.000 668.920 ;
        RECT 204.400 613.840 1096.000 615.240 ;
        RECT 204.000 610.480 1096.000 613.840 ;
        RECT 204.000 609.080 1095.600 610.480 ;
        RECT 204.000 550.640 1096.000 609.080 ;
        RECT 204.000 549.240 1095.600 550.640 ;
        RECT 204.000 529.560 1096.000 549.240 ;
        RECT 204.400 528.160 1096.000 529.560 ;
        RECT 204.000 490.800 1096.000 528.160 ;
        RECT 204.000 489.400 1095.600 490.800 ;
        RECT 204.000 443.880 1096.000 489.400 ;
        RECT 204.400 442.480 1096.000 443.880 ;
        RECT 204.000 430.960 1096.000 442.480 ;
        RECT 204.000 429.560 1095.600 430.960 ;
        RECT 204.000 410.715 1096.000 429.560 ;
      LAYER met4 ;
        RECT 515.855 951.655 527.840 988.025 ;
        RECT 530.240 951.655 604.640 988.025 ;
        RECT 607.040 951.655 680.865 988.025 ;
  END
END user_project_wrapper
END LIBRARY

