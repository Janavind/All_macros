magic
tech sky130A
magscale 1 2
timestamp 1654286010
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 117836
<< metal2 >>
rect 662 119200 718 120000
rect 2042 119200 2098 120000
rect 3514 119200 3570 120000
rect 4986 119200 5042 120000
rect 6458 119200 6514 120000
rect 7930 119200 7986 120000
rect 9402 119200 9458 120000
rect 10874 119200 10930 120000
rect 12346 119200 12402 120000
rect 13818 119200 13874 120000
rect 15290 119200 15346 120000
rect 16762 119200 16818 120000
rect 18142 119200 18198 120000
rect 19614 119200 19670 120000
rect 21086 119200 21142 120000
rect 22558 119200 22614 120000
rect 24030 119200 24086 120000
rect 25502 119200 25558 120000
rect 26974 119200 27030 120000
rect 28446 119200 28502 120000
rect 29918 119200 29974 120000
rect 31390 119200 31446 120000
rect 32862 119200 32918 120000
rect 34242 119200 34298 120000
rect 35714 119200 35770 120000
rect 37186 119200 37242 120000
rect 38658 119200 38714 120000
rect 40130 119200 40186 120000
rect 41602 119200 41658 120000
rect 43074 119200 43130 120000
rect 44546 119200 44602 120000
rect 46018 119200 46074 120000
rect 47490 119200 47546 120000
rect 48962 119200 49018 120000
rect 50342 119200 50398 120000
rect 51814 119200 51870 120000
rect 53286 119200 53342 120000
rect 54758 119200 54814 120000
rect 56230 119200 56286 120000
rect 57702 119200 57758 120000
rect 59174 119200 59230 120000
rect 60646 119200 60702 120000
rect 62118 119200 62174 120000
rect 63590 119200 63646 120000
rect 65062 119200 65118 120000
rect 66442 119200 66498 120000
rect 67914 119200 67970 120000
rect 69386 119200 69442 120000
rect 70858 119200 70914 120000
rect 72330 119200 72386 120000
rect 73802 119200 73858 120000
rect 75274 119200 75330 120000
rect 76746 119200 76802 120000
rect 78218 119200 78274 120000
rect 79690 119200 79746 120000
rect 81162 119200 81218 120000
rect 82542 119200 82598 120000
rect 84014 119200 84070 120000
rect 85486 119200 85542 120000
rect 86958 119200 87014 120000
rect 88430 119200 88486 120000
rect 89902 119200 89958 120000
rect 91374 119200 91430 120000
rect 92846 119200 92902 120000
rect 94318 119200 94374 120000
rect 95790 119200 95846 120000
rect 97262 119200 97318 120000
rect 98734 119200 98790 120000
rect 100114 119200 100170 120000
rect 101586 119200 101642 120000
rect 103058 119200 103114 120000
rect 104530 119200 104586 120000
rect 106002 119200 106058 120000
rect 107474 119200 107530 120000
rect 108946 119200 109002 120000
rect 110418 119200 110474 120000
rect 111890 119200 111946 120000
rect 113362 119200 113418 120000
rect 114834 119200 114890 120000
rect 116214 119200 116270 120000
rect 117686 119200 117742 120000
rect 119158 119200 119214 120000
rect 120630 119200 120686 120000
rect 122102 119200 122158 120000
rect 123574 119200 123630 120000
rect 125046 119200 125102 120000
rect 126518 119200 126574 120000
rect 127990 119200 128046 120000
rect 129462 119200 129518 120000
rect 130934 119200 130990 120000
rect 132314 119200 132370 120000
rect 133786 119200 133842 120000
rect 135258 119200 135314 120000
rect 136730 119200 136786 120000
rect 138202 119200 138258 120000
rect 139674 119200 139730 120000
rect 141146 119200 141202 120000
rect 142618 119200 142674 120000
rect 144090 119200 144146 120000
rect 145562 119200 145618 120000
rect 147034 119200 147090 120000
rect 148414 119200 148470 120000
rect 149886 119200 149942 120000
rect 151358 119200 151414 120000
rect 152830 119200 152886 120000
rect 154302 119200 154358 120000
rect 155774 119200 155830 120000
rect 157246 119200 157302 120000
rect 158718 119200 158774 120000
rect 160190 119200 160246 120000
rect 161662 119200 161718 120000
rect 163134 119200 163190 120000
rect 164514 119200 164570 120000
rect 165986 119200 166042 120000
rect 167458 119200 167514 120000
rect 168930 119200 168986 120000
rect 170402 119200 170458 120000
rect 171874 119200 171930 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21270 0 21326 800
rect 21638 0 21694 800
rect 22006 0 22062 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24214 0 24270 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58438 0 58494 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67362 0 67418 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 69938 0 69994 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 71042 0 71098 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74262 0 74318 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76746 0 76802 800
rect 77114 0 77170 800
rect 77482 0 77538 800
rect 77850 0 77906 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100850 0 100906 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102690 0 102746 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104162 0 104218 800
rect 104530 0 104586 800
rect 104806 0 104862 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105910 0 105966 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107750 0 107806 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 110970 0 111026 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112810 0 112866 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116766 0 116822 800
rect 117134 0 117190 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122470 0 122526 800
rect 122838 0 122894 800
rect 123206 0 123262 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127162 0 127218 800
rect 127530 0 127586 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143722 0 143778 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145194 0 145250 800
rect 145562 0 145618 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 150898 0 150954 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155222 0 155278 800
rect 155590 0 155646 800
rect 155958 0 156014 800
rect 156326 0 156382 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159178 0 159234 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162122 0 162178 800
rect 162490 0 162546 800
rect 162858 0 162914 800
rect 163226 0 163282 800
rect 163502 0 163558 800
rect 163870 0 163926 800
rect 164238 0 164294 800
rect 164606 0 164662 800
rect 164974 0 165030 800
rect 165342 0 165398 800
rect 165710 0 165766 800
rect 166078 0 166134 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 167826 0 167882 800
rect 168194 0 168250 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 170034 0 170090 800
rect 170402 0 170458 800
rect 170770 0 170826 800
rect 171138 0 171194 800
rect 171506 0 171562 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 774 119144 1986 119354
rect 2154 119144 3458 119354
rect 3626 119144 4930 119354
rect 5098 119144 6402 119354
rect 6570 119144 7874 119354
rect 8042 119144 9346 119354
rect 9514 119144 10818 119354
rect 10986 119144 12290 119354
rect 12458 119144 13762 119354
rect 13930 119144 15234 119354
rect 15402 119144 16706 119354
rect 16874 119144 18086 119354
rect 18254 119144 19558 119354
rect 19726 119144 21030 119354
rect 21198 119144 22502 119354
rect 22670 119144 23974 119354
rect 24142 119144 25446 119354
rect 25614 119144 26918 119354
rect 27086 119144 28390 119354
rect 28558 119144 29862 119354
rect 30030 119144 31334 119354
rect 31502 119144 32806 119354
rect 32974 119144 34186 119354
rect 34354 119144 35658 119354
rect 35826 119144 37130 119354
rect 37298 119144 38602 119354
rect 38770 119144 40074 119354
rect 40242 119144 41546 119354
rect 41714 119144 43018 119354
rect 43186 119144 44490 119354
rect 44658 119144 45962 119354
rect 46130 119144 47434 119354
rect 47602 119144 48906 119354
rect 49074 119144 50286 119354
rect 50454 119144 51758 119354
rect 51926 119144 53230 119354
rect 53398 119144 54702 119354
rect 54870 119144 56174 119354
rect 56342 119144 57646 119354
rect 57814 119144 59118 119354
rect 59286 119144 60590 119354
rect 60758 119144 62062 119354
rect 62230 119144 63534 119354
rect 63702 119144 65006 119354
rect 65174 119144 66386 119354
rect 66554 119144 67858 119354
rect 68026 119144 69330 119354
rect 69498 119144 70802 119354
rect 70970 119144 72274 119354
rect 72442 119144 73746 119354
rect 73914 119144 75218 119354
rect 75386 119144 76690 119354
rect 76858 119144 78162 119354
rect 78330 119144 79634 119354
rect 79802 119144 81106 119354
rect 81274 119144 82486 119354
rect 82654 119144 83958 119354
rect 84126 119144 85430 119354
rect 85598 119144 86902 119354
rect 87070 119144 88374 119354
rect 88542 119144 89846 119354
rect 90014 119144 91318 119354
rect 91486 119144 92790 119354
rect 92958 119144 94262 119354
rect 94430 119144 95734 119354
rect 95902 119144 97206 119354
rect 97374 119144 98678 119354
rect 98846 119144 100058 119354
rect 100226 119144 101530 119354
rect 101698 119144 103002 119354
rect 103170 119144 104474 119354
rect 104642 119144 105946 119354
rect 106114 119144 107418 119354
rect 107586 119144 108890 119354
rect 109058 119144 110362 119354
rect 110530 119144 111834 119354
rect 112002 119144 113306 119354
rect 113474 119144 114778 119354
rect 114946 119144 116158 119354
rect 116326 119144 117630 119354
rect 117798 119144 119102 119354
rect 119270 119144 120574 119354
rect 120742 119144 122046 119354
rect 122214 119144 123518 119354
rect 123686 119144 124990 119354
rect 125158 119144 126462 119354
rect 126630 119144 127934 119354
rect 128102 119144 129406 119354
rect 129574 119144 130878 119354
rect 131046 119144 132258 119354
rect 132426 119144 133730 119354
rect 133898 119144 135202 119354
rect 135370 119144 136674 119354
rect 136842 119144 138146 119354
rect 138314 119144 139618 119354
rect 139786 119144 141090 119354
rect 141258 119144 142562 119354
rect 142730 119144 144034 119354
rect 144202 119144 145506 119354
rect 145674 119144 146978 119354
rect 147146 119144 148358 119354
rect 148526 119144 149830 119354
rect 149998 119144 151302 119354
rect 151470 119144 152774 119354
rect 152942 119144 154246 119354
rect 154414 119144 155718 119354
rect 155886 119144 157190 119354
rect 157358 119144 158662 119354
rect 158830 119144 160134 119354
rect 160302 119144 161606 119354
rect 161774 119144 163078 119354
rect 163246 119144 164458 119354
rect 164626 119144 165930 119354
rect 166098 119144 167402 119354
rect 167570 119144 168874 119354
rect 169042 119144 170346 119354
rect 170514 119144 171818 119354
rect 171986 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3274 856
rect 3442 800 3642 856
rect 3810 800 4010 856
rect 4178 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6494 856
rect 6662 800 6862 856
rect 7030 800 7230 856
rect 7398 800 7598 856
rect 7766 800 7966 856
rect 8134 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9346 856
rect 9514 800 9714 856
rect 9882 800 10082 856
rect 10250 800 10450 856
rect 10618 800 10818 856
rect 10986 800 11186 856
rect 11354 800 11554 856
rect 11722 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12566 856
rect 12734 800 12934 856
rect 13102 800 13302 856
rect 13470 800 13670 856
rect 13838 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15878 856
rect 16046 800 16246 856
rect 16414 800 16614 856
rect 16782 800 16890 856
rect 17058 800 17258 856
rect 17426 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18730 856
rect 18898 800 19098 856
rect 19266 800 19466 856
rect 19634 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21214 856
rect 21382 800 21582 856
rect 21750 800 21950 856
rect 22118 800 22318 856
rect 22486 800 22686 856
rect 22854 800 23054 856
rect 23222 800 23422 856
rect 23590 800 23790 856
rect 23958 800 24158 856
rect 24326 800 24526 856
rect 24694 800 24894 856
rect 25062 800 25170 856
rect 25338 800 25538 856
rect 25706 800 25906 856
rect 26074 800 26274 856
rect 26442 800 26642 856
rect 26810 800 27010 856
rect 27178 800 27378 856
rect 27546 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28482 856
rect 28650 800 28850 856
rect 29018 800 29218 856
rect 29386 800 29494 856
rect 29662 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31334 856
rect 31502 800 31702 856
rect 31870 800 32070 856
rect 32238 800 32438 856
rect 32606 800 32806 856
rect 32974 800 33174 856
rect 33342 800 33542 856
rect 33710 800 33818 856
rect 33986 800 34186 856
rect 34354 800 34554 856
rect 34722 800 34922 856
rect 35090 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37774 856
rect 37942 800 38142 856
rect 38310 800 38510 856
rect 38678 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39614 856
rect 39782 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42098 856
rect 42266 800 42466 856
rect 42634 800 42834 856
rect 43002 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43938 856
rect 44106 800 44306 856
rect 44474 800 44674 856
rect 44842 800 45042 856
rect 45210 800 45410 856
rect 45578 800 45778 856
rect 45946 800 46054 856
rect 46222 800 46422 856
rect 46590 800 46790 856
rect 46958 800 47158 856
rect 47326 800 47526 856
rect 47694 800 47894 856
rect 48062 800 48262 856
rect 48430 800 48630 856
rect 48798 800 48998 856
rect 49166 800 49366 856
rect 49534 800 49734 856
rect 49902 800 50102 856
rect 50270 800 50378 856
rect 50546 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51482 856
rect 51650 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52586 856
rect 52754 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53690 856
rect 53858 800 54058 856
rect 54226 800 54426 856
rect 54594 800 54702 856
rect 54870 800 55070 856
rect 55238 800 55438 856
rect 55606 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56542 856
rect 56710 800 56910 856
rect 57078 800 57278 856
rect 57446 800 57646 856
rect 57814 800 58014 856
rect 58182 800 58382 856
rect 58550 800 58658 856
rect 58826 800 59026 856
rect 59194 800 59394 856
rect 59562 800 59762 856
rect 59930 800 60130 856
rect 60298 800 60498 856
rect 60666 800 60866 856
rect 61034 800 61234 856
rect 61402 800 61602 856
rect 61770 800 61970 856
rect 62138 800 62338 856
rect 62506 800 62706 856
rect 62874 800 62982 856
rect 63150 800 63350 856
rect 63518 800 63718 856
rect 63886 800 64086 856
rect 64254 800 64454 856
rect 64622 800 64822 856
rect 64990 800 65190 856
rect 65358 800 65558 856
rect 65726 800 65926 856
rect 66094 800 66294 856
rect 66462 800 66662 856
rect 66830 800 67030 856
rect 67198 800 67306 856
rect 67474 800 67674 856
rect 67842 800 68042 856
rect 68210 800 68410 856
rect 68578 800 68778 856
rect 68946 800 69146 856
rect 69314 800 69514 856
rect 69682 800 69882 856
rect 70050 800 70250 856
rect 70418 800 70618 856
rect 70786 800 70986 856
rect 71154 800 71262 856
rect 71430 800 71630 856
rect 71798 800 71998 856
rect 72166 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73838 856
rect 74006 800 74206 856
rect 74374 800 74574 856
rect 74742 800 74942 856
rect 75110 800 75310 856
rect 75478 800 75586 856
rect 75754 800 75954 856
rect 76122 800 76322 856
rect 76490 800 76690 856
rect 76858 800 77058 856
rect 77226 800 77426 856
rect 77594 800 77794 856
rect 77962 800 78162 856
rect 78330 800 78530 856
rect 78698 800 78898 856
rect 79066 800 79266 856
rect 79434 800 79542 856
rect 79710 800 79910 856
rect 80078 800 80278 856
rect 80446 800 80646 856
rect 80814 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81750 856
rect 81918 800 82118 856
rect 82286 800 82486 856
rect 82654 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84602 856
rect 84770 800 84970 856
rect 85138 800 85338 856
rect 85506 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88190 856
rect 88358 800 88558 856
rect 88726 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90398 856
rect 90566 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91870 856
rect 92038 800 92146 856
rect 92314 800 92514 856
rect 92682 800 92882 856
rect 93050 800 93250 856
rect 93418 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95458 856
rect 95626 800 95826 856
rect 95994 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97206 856
rect 97374 800 97574 856
rect 97742 800 97942 856
rect 98110 800 98310 856
rect 98478 800 98678 856
rect 98846 800 99046 856
rect 99214 800 99414 856
rect 99582 800 99782 856
rect 99950 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100794 856
rect 100962 800 101162 856
rect 101330 800 101530 856
rect 101698 800 101898 856
rect 102066 800 102266 856
rect 102434 800 102634 856
rect 102802 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104106 856
rect 104274 800 104474 856
rect 104642 800 104750 856
rect 104918 800 105118 856
rect 105286 800 105486 856
rect 105654 800 105854 856
rect 106022 800 106222 856
rect 106390 800 106590 856
rect 106758 800 106958 856
rect 107126 800 107326 856
rect 107494 800 107694 856
rect 107862 800 108062 856
rect 108230 800 108430 856
rect 108598 800 108798 856
rect 108966 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110546 856
rect 110714 800 110914 856
rect 111082 800 111282 856
rect 111450 800 111650 856
rect 111818 800 112018 856
rect 112186 800 112386 856
rect 112554 800 112754 856
rect 112922 800 113030 856
rect 113198 800 113398 856
rect 113566 800 113766 856
rect 113934 800 114134 856
rect 114302 800 114502 856
rect 114670 800 114870 856
rect 115038 800 115238 856
rect 115406 800 115606 856
rect 115774 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116710 856
rect 116878 800 117078 856
rect 117246 800 117354 856
rect 117522 800 117722 856
rect 117890 800 118090 856
rect 118258 800 118458 856
rect 118626 800 118826 856
rect 118994 800 119194 856
rect 119362 800 119562 856
rect 119730 800 119930 856
rect 120098 800 120298 856
rect 120466 800 120666 856
rect 120834 800 121034 856
rect 121202 800 121402 856
rect 121570 800 121678 856
rect 121846 800 122046 856
rect 122214 800 122414 856
rect 122582 800 122782 856
rect 122950 800 123150 856
rect 123318 800 123518 856
rect 123686 800 123886 856
rect 124054 800 124254 856
rect 124422 800 124622 856
rect 124790 800 124990 856
rect 125158 800 125358 856
rect 125526 800 125634 856
rect 125802 800 126002 856
rect 126170 800 126370 856
rect 126538 800 126738 856
rect 126906 800 127106 856
rect 127274 800 127474 856
rect 127642 800 127842 856
rect 128010 800 128210 856
rect 128378 800 128578 856
rect 128746 800 128946 856
rect 129114 800 129314 856
rect 129482 800 129682 856
rect 129850 800 129958 856
rect 130126 800 130326 856
rect 130494 800 130694 856
rect 130862 800 131062 856
rect 131230 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132166 856
rect 132334 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133270 856
rect 133438 800 133638 856
rect 133806 800 134006 856
rect 134174 800 134282 856
rect 134450 800 134650 856
rect 134818 800 135018 856
rect 135186 800 135386 856
rect 135554 800 135754 856
rect 135922 800 136122 856
rect 136290 800 136490 856
rect 136658 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137594 856
rect 137762 800 137962 856
rect 138130 800 138238 856
rect 138406 800 138606 856
rect 138774 800 138974 856
rect 139142 800 139342 856
rect 139510 800 139710 856
rect 139878 800 140078 856
rect 140246 800 140446 856
rect 140614 800 140814 856
rect 140982 800 141182 856
rect 141350 800 141550 856
rect 141718 800 141918 856
rect 142086 800 142286 856
rect 142454 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143298 856
rect 143466 800 143666 856
rect 143834 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144770 856
rect 144938 800 145138 856
rect 145306 800 145506 856
rect 145674 800 145874 856
rect 146042 800 146242 856
rect 146410 800 146518 856
rect 146686 800 146886 856
rect 147054 800 147254 856
rect 147422 800 147622 856
rect 147790 800 147990 856
rect 148158 800 148358 856
rect 148526 800 148726 856
rect 148894 800 149094 856
rect 149262 800 149462 856
rect 149630 800 149830 856
rect 149998 800 150198 856
rect 150366 800 150566 856
rect 150734 800 150842 856
rect 151010 800 151210 856
rect 151378 800 151578 856
rect 151746 800 151946 856
rect 152114 800 152314 856
rect 152482 800 152682 856
rect 152850 800 153050 856
rect 153218 800 153418 856
rect 153586 800 153786 856
rect 153954 800 154154 856
rect 154322 800 154522 856
rect 154690 800 154890 856
rect 155058 800 155166 856
rect 155334 800 155534 856
rect 155702 800 155902 856
rect 156070 800 156270 856
rect 156438 800 156638 856
rect 156806 800 157006 856
rect 157174 800 157374 856
rect 157542 800 157742 856
rect 157910 800 158110 856
rect 158278 800 158478 856
rect 158646 800 158846 856
rect 159014 800 159122 856
rect 159290 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160594 856
rect 160762 800 160962 856
rect 161130 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162066 856
rect 162234 800 162434 856
rect 162602 800 162802 856
rect 162970 800 163170 856
rect 163338 800 163446 856
rect 163614 800 163814 856
rect 163982 800 164182 856
rect 164350 800 164550 856
rect 164718 800 164918 856
rect 165086 800 165286 856
rect 165454 800 165654 856
rect 165822 800 166022 856
rect 166190 800 166390 856
rect 166558 800 166758 856
rect 166926 800 167126 856
rect 167294 800 167494 856
rect 167662 800 167770 856
rect 167938 800 168138 856
rect 168306 800 168506 856
rect 168674 800 168874 856
rect 169042 800 169242 856
rect 169410 800 169610 856
rect 169778 800 169978 856
rect 170146 800 170346 856
rect 170514 800 170714 856
rect 170882 800 171082 856
rect 171250 800 171450 856
rect 171618 800 171726 856
rect 171894 800 172094 856
rect 172262 800 172462 856
rect 172630 800 172830 856
rect 172998 800 173198 856
rect 173366 800 173566 856
rect 173734 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
rect 175574 800 175774 856
rect 175942 800 176050 856
rect 176218 800 176418 856
rect 176586 800 176786 856
rect 176954 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178186 856
<< metal3 >>
rect 179200 113296 180000 113416
rect 0 109896 800 110016
rect 179200 99968 180000 100088
rect 0 89904 800 90024
rect 179200 86640 180000 86760
rect 179200 73312 180000 73432
rect 0 69912 800 70032
rect 179200 59984 180000 60104
rect 0 49920 800 50040
rect 179200 46656 180000 46776
rect 179200 33328 180000 33448
rect 0 29928 800 30048
rect 179200 20000 180000 20120
rect 0 9936 800 10056
rect 179200 6672 180000 6792
<< obsm3 >>
rect 800 113496 179200 117537
rect 800 113216 179120 113496
rect 800 110096 179200 113216
rect 880 109816 179200 110096
rect 800 100168 179200 109816
rect 800 99888 179120 100168
rect 800 90104 179200 99888
rect 880 89824 179200 90104
rect 800 86840 179200 89824
rect 800 86560 179120 86840
rect 800 73512 179200 86560
rect 800 73232 179120 73512
rect 800 70112 179200 73232
rect 880 69832 179200 70112
rect 800 60184 179200 69832
rect 800 59904 179120 60184
rect 800 50120 179200 59904
rect 880 49840 179200 50120
rect 800 46856 179200 49840
rect 800 46576 179120 46856
rect 800 33528 179200 46576
rect 800 33248 179120 33528
rect 800 30128 179200 33248
rect 880 29848 179200 30128
rect 800 20200 179200 29848
rect 800 19920 179120 20200
rect 800 10136 179200 19920
rect 880 9856 179200 10136
rect 800 6872 179200 9856
rect 800 6592 179120 6872
rect 800 2143 179200 6592
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 84883 3299 91021 116381
<< labels >>
rlabel metal3 s 0 9936 800 10056 6 active
port 1 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 0 69912 800 70032 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 0 89904 800 90024 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 179200 73312 180000 73432 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 171874 119200 171930 120000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal3 s 0 109896 800 110016 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 179200 86640 180000 86760 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 179200 33328 180000 33448 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal3 s 179200 99968 180000 100088 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 179200 113296 180000 113416 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal2 s 167458 119200 167514 120000 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 0 29928 800 30048 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 0 49920 800 50040 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 179200 46656 180000 46776 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal2 s 168930 119200 168986 120000 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal2 s 170402 119200 170458 120000 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 179200 59984 180000 60104 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 44546 119200 44602 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 48962 119200 49018 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 53286 119200 53342 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 57702 119200 57758 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 62118 119200 62174 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 66442 119200 66498 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 70858 119200 70914 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 75274 119200 75330 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 79690 119200 79746 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 84014 119200 84070 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 4986 119200 5042 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 88430 119200 88486 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 92846 119200 92902 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 97262 119200 97318 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 101586 119200 101642 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 106002 119200 106058 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 110418 119200 110474 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 114834 119200 114890 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 123574 119200 123630 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 127990 119200 128046 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9402 119200 9458 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 132314 119200 132370 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 136730 119200 136786 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 141146 119200 141202 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 145562 119200 145618 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 149886 119200 149942 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 154302 119200 154358 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 158718 119200 158774 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 163134 119200 163190 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 13818 119200 13874 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18142 119200 18198 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 22558 119200 22614 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 26974 119200 27030 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31390 119200 31446 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 35714 119200 35770 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 40130 119200 40186 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2042 119200 2098 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 46018 119200 46074 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 50342 119200 50398 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 54758 119200 54814 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 59174 119200 59230 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 63590 119200 63646 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 67914 119200 67970 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 72330 119200 72386 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 76746 119200 76802 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 81162 119200 81218 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 85486 119200 85542 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6458 119200 6514 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 94318 119200 94374 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 98734 119200 98790 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 103058 119200 103114 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 107474 119200 107530 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 116214 119200 116270 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 120630 119200 120686 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 125046 119200 125102 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 129462 119200 129518 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 10874 119200 10930 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 133786 119200 133842 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 138202 119200 138258 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 142618 119200 142674 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 147034 119200 147090 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 151358 119200 151414 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 155774 119200 155830 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 160190 119200 160246 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 164514 119200 164570 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15290 119200 15346 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 19614 119200 19670 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24030 119200 24086 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28446 119200 28502 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 32862 119200 32918 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 37186 119200 37242 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 41602 119200 41658 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3514 119200 3570 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 47490 119200 47546 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 51814 119200 51870 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 56230 119200 56286 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 60646 119200 60702 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 65062 119200 65118 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 69386 119200 69442 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 73802 119200 73858 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 78218 119200 78274 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 86958 119200 87014 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 7930 119200 7986 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 91374 119200 91430 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 95790 119200 95846 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 100114 119200 100170 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 104530 119200 104586 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 108946 119200 109002 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 113362 119200 113418 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 117686 119200 117742 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 122102 119200 122158 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 126518 119200 126574 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 130934 119200 130990 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12346 119200 12402 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 135258 119200 135314 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 139674 119200 139730 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 144090 119200 144146 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 148414 119200 148470 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 152830 119200 152886 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 157246 119200 157302 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 161662 119200 161718 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 165986 119200 166042 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 16762 119200 16818 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21086 119200 21142 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25502 119200 25558 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 29918 119200 29974 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 34242 119200 34298 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 38658 119200 38714 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 43074 119200 43130 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 164606 0 164662 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 161754 0 161810 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 167182 0 167238 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 168194 0 168250 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86130 0 86186 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 179200 6672 180000 6792 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 179200 20000 180000 20120 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 user_irq[1]
port 531 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6507630
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_no_fill.magic.gds
string GDS_START 297240
<< end >>

