magic
tech sky130A
magscale 1 2
timestamp 1653457307
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 658 2128 178848 118720
<< metal2 >>
rect 662 119200 718 120000
rect 2042 119200 2098 120000
rect 3422 119200 3478 120000
rect 4894 119200 4950 120000
rect 6274 119200 6330 120000
rect 7746 119200 7802 120000
rect 9126 119200 9182 120000
rect 10506 119200 10562 120000
rect 11978 119200 12034 120000
rect 13358 119200 13414 120000
rect 14830 119200 14886 120000
rect 16210 119200 16266 120000
rect 17590 119200 17646 120000
rect 19062 119200 19118 120000
rect 20442 119200 20498 120000
rect 21914 119200 21970 120000
rect 23294 119200 23350 120000
rect 24674 119200 24730 120000
rect 26146 119200 26202 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30378 119200 30434 120000
rect 31850 119200 31906 120000
rect 33230 119200 33286 120000
rect 34610 119200 34666 120000
rect 36082 119200 36138 120000
rect 37462 119200 37518 120000
rect 38934 119200 38990 120000
rect 40314 119200 40370 120000
rect 41694 119200 41750 120000
rect 43166 119200 43222 120000
rect 44546 119200 44602 120000
rect 46018 119200 46074 120000
rect 47398 119200 47454 120000
rect 48778 119200 48834 120000
rect 50250 119200 50306 120000
rect 51630 119200 51686 120000
rect 53102 119200 53158 120000
rect 54482 119200 54538 120000
rect 55862 119200 55918 120000
rect 57334 119200 57390 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61566 119200 61622 120000
rect 63038 119200 63094 120000
rect 64418 119200 64474 120000
rect 65798 119200 65854 120000
rect 67270 119200 67326 120000
rect 68650 119200 68706 120000
rect 70122 119200 70178 120000
rect 71502 119200 71558 120000
rect 72882 119200 72938 120000
rect 74354 119200 74410 120000
rect 75734 119200 75790 120000
rect 77206 119200 77262 120000
rect 78586 119200 78642 120000
rect 79966 119200 80022 120000
rect 81438 119200 81494 120000
rect 82818 119200 82874 120000
rect 84290 119200 84346 120000
rect 85670 119200 85726 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89902 119200 89958 120000
rect 91374 119200 91430 120000
rect 92754 119200 92810 120000
rect 94226 119200 94282 120000
rect 95606 119200 95662 120000
rect 96986 119200 97042 120000
rect 98458 119200 98514 120000
rect 99838 119200 99894 120000
rect 101310 119200 101366 120000
rect 102690 119200 102746 120000
rect 104070 119200 104126 120000
rect 105542 119200 105598 120000
rect 106922 119200 106978 120000
rect 108394 119200 108450 120000
rect 109774 119200 109830 120000
rect 111154 119200 111210 120000
rect 112626 119200 112682 120000
rect 114006 119200 114062 120000
rect 115478 119200 115534 120000
rect 116858 119200 116914 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121090 119200 121146 120000
rect 122562 119200 122618 120000
rect 123942 119200 123998 120000
rect 125414 119200 125470 120000
rect 126794 119200 126850 120000
rect 128174 119200 128230 120000
rect 129646 119200 129702 120000
rect 131026 119200 131082 120000
rect 132498 119200 132554 120000
rect 133878 119200 133934 120000
rect 135258 119200 135314 120000
rect 136730 119200 136786 120000
rect 138110 119200 138166 120000
rect 139582 119200 139638 120000
rect 140962 119200 141018 120000
rect 142342 119200 142398 120000
rect 143814 119200 143870 120000
rect 145194 119200 145250 120000
rect 146666 119200 146722 120000
rect 148046 119200 148102 120000
rect 149426 119200 149482 120000
rect 150898 119200 150954 120000
rect 152278 119200 152334 120000
rect 153750 119200 153806 120000
rect 155130 119200 155186 120000
rect 156602 119200 156658 120000
rect 157982 119200 158038 120000
rect 159362 119200 159418 120000
rect 160834 119200 160890 120000
rect 162214 119200 162270 120000
rect 163686 119200 163742 120000
rect 165066 119200 165122 120000
rect 166446 119200 166502 120000
rect 167918 119200 167974 120000
rect 169298 119200 169354 120000
rect 170770 119200 170826 120000
rect 172150 119200 172206 120000
rect 173530 119200 173586 120000
rect 175002 119200 175058 120000
rect 176382 119200 176438 120000
rect 177854 119200 177910 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40130 0 40186 800
rect 40498 0 40554 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46018 0 46074 800
rect 46386 0 46442 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 51078 0 51134 800
rect 51446 0 51502 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54758 0 54814 800
rect 55126 0 55182 800
rect 55494 0 55550 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61290 0 61346 800
rect 61658 0 61714 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 66074 0 66130 800
rect 66442 0 66498 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 78034 0 78090 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79506 0 79562 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85670 0 85726 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93766 0 93822 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
rect 113454 0 113510 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116306 0 116362 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117410 0 117466 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119618 0 119674 800
rect 119986 0 120042 800
rect 120354 0 120410 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123574 0 123630 800
rect 123942 0 123998 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128726 0 128782 800
rect 129094 0 129150 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130934 0 130990 800
rect 131302 0 131358 800
rect 131670 0 131726 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134522 0 134578 800
rect 134890 0 134946 800
rect 135258 0 135314 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138570 0 138626 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139674 0 139730 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148782 0 148838 800
rect 149150 0 149206 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154946 0 155002 800
rect 155314 0 155370 800
rect 155682 0 155738 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157522 0 157578 800
rect 157890 0 157946 800
rect 158258 0 158314 800
rect 158626 0 158682 800
rect 158994 0 159050 800
rect 159362 0 159418 800
rect 159730 0 159786 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161478 0 161534 800
rect 161846 0 161902 800
rect 162214 0 162270 800
rect 162582 0 162638 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165158 0 165214 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166262 0 166318 800
rect 166630 0 166686 800
rect 166998 0 167054 800
rect 167366 0 167422 800
rect 167734 0 167790 800
rect 168102 0 168158 800
rect 168470 0 168526 800
rect 168838 0 168894 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 170954 0 171010 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173162 0 173218 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 774 119144 1986 119354
rect 2154 119144 3366 119354
rect 3534 119144 4838 119354
rect 5006 119144 6218 119354
rect 6386 119144 7690 119354
rect 7858 119144 9070 119354
rect 9238 119144 10450 119354
rect 10618 119144 11922 119354
rect 12090 119144 13302 119354
rect 13470 119144 14774 119354
rect 14942 119144 16154 119354
rect 16322 119144 17534 119354
rect 17702 119144 19006 119354
rect 19174 119144 20386 119354
rect 20554 119144 21858 119354
rect 22026 119144 23238 119354
rect 23406 119144 24618 119354
rect 24786 119144 26090 119354
rect 26258 119144 27470 119354
rect 27638 119144 28942 119354
rect 29110 119144 30322 119354
rect 30490 119144 31794 119354
rect 31962 119144 33174 119354
rect 33342 119144 34554 119354
rect 34722 119144 36026 119354
rect 36194 119144 37406 119354
rect 37574 119144 38878 119354
rect 39046 119144 40258 119354
rect 40426 119144 41638 119354
rect 41806 119144 43110 119354
rect 43278 119144 44490 119354
rect 44658 119144 45962 119354
rect 46130 119144 47342 119354
rect 47510 119144 48722 119354
rect 48890 119144 50194 119354
rect 50362 119144 51574 119354
rect 51742 119144 53046 119354
rect 53214 119144 54426 119354
rect 54594 119144 55806 119354
rect 55974 119144 57278 119354
rect 57446 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61510 119354
rect 61678 119144 62982 119354
rect 63150 119144 64362 119354
rect 64530 119144 65742 119354
rect 65910 119144 67214 119354
rect 67382 119144 68594 119354
rect 68762 119144 70066 119354
rect 70234 119144 71446 119354
rect 71614 119144 72826 119354
rect 72994 119144 74298 119354
rect 74466 119144 75678 119354
rect 75846 119144 77150 119354
rect 77318 119144 78530 119354
rect 78698 119144 79910 119354
rect 80078 119144 81382 119354
rect 81550 119144 82762 119354
rect 82930 119144 84234 119354
rect 84402 119144 85614 119354
rect 85782 119144 86994 119354
rect 87162 119144 88466 119354
rect 88634 119144 89846 119354
rect 90014 119144 91318 119354
rect 91486 119144 92698 119354
rect 92866 119144 94170 119354
rect 94338 119144 95550 119354
rect 95718 119144 96930 119354
rect 97098 119144 98402 119354
rect 98570 119144 99782 119354
rect 99950 119144 101254 119354
rect 101422 119144 102634 119354
rect 102802 119144 104014 119354
rect 104182 119144 105486 119354
rect 105654 119144 106866 119354
rect 107034 119144 108338 119354
rect 108506 119144 109718 119354
rect 109886 119144 111098 119354
rect 111266 119144 112570 119354
rect 112738 119144 113950 119354
rect 114118 119144 115422 119354
rect 115590 119144 116802 119354
rect 116970 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121034 119354
rect 121202 119144 122506 119354
rect 122674 119144 123886 119354
rect 124054 119144 125358 119354
rect 125526 119144 126738 119354
rect 126906 119144 128118 119354
rect 128286 119144 129590 119354
rect 129758 119144 130970 119354
rect 131138 119144 132442 119354
rect 132610 119144 133822 119354
rect 133990 119144 135202 119354
rect 135370 119144 136674 119354
rect 136842 119144 138054 119354
rect 138222 119144 139526 119354
rect 139694 119144 140906 119354
rect 141074 119144 142286 119354
rect 142454 119144 143758 119354
rect 143926 119144 145138 119354
rect 145306 119144 146610 119354
rect 146778 119144 147990 119354
rect 148158 119144 149370 119354
rect 149538 119144 150842 119354
rect 151010 119144 152222 119354
rect 152390 119144 153694 119354
rect 153862 119144 155074 119354
rect 155242 119144 156546 119354
rect 156714 119144 157926 119354
rect 158094 119144 159306 119354
rect 159474 119144 160778 119354
rect 160946 119144 162158 119354
rect 162326 119144 163630 119354
rect 163798 119144 165010 119354
rect 165178 119144 166390 119354
rect 166558 119144 167862 119354
rect 168030 119144 169242 119354
rect 169410 119144 170714 119354
rect 170882 119144 172094 119354
rect 172262 119144 173474 119354
rect 173642 119144 174946 119354
rect 175114 119144 176326 119354
rect 176494 119144 177798 119354
rect 177966 119144 178186 119354
rect 664 856 178186 119144
rect 664 734 698 856
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7322 856
rect 7490 734 7690 856
rect 7858 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8794 856
rect 8962 734 9162 856
rect 9330 734 9530 856
rect 9698 734 9806 856
rect 9974 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12750 856
rect 12918 734 13118 856
rect 13286 734 13486 856
rect 13654 734 13854 856
rect 14022 734 14222 856
rect 14390 734 14590 856
rect 14758 734 14958 856
rect 15126 734 15326 856
rect 15494 734 15694 856
rect 15862 734 16062 856
rect 16230 734 16430 856
rect 16598 734 16798 856
rect 16966 734 17166 856
rect 17334 734 17534 856
rect 17702 734 17902 856
rect 18070 734 18270 856
rect 18438 734 18638 856
rect 18806 734 19006 856
rect 19174 734 19282 856
rect 19450 734 19650 856
rect 19818 734 20018 856
rect 20186 734 20386 856
rect 20554 734 20754 856
rect 20922 734 21122 856
rect 21290 734 21490 856
rect 21658 734 21858 856
rect 22026 734 22226 856
rect 22394 734 22594 856
rect 22762 734 22962 856
rect 23130 734 23330 856
rect 23498 734 23698 856
rect 23866 734 24066 856
rect 24234 734 24434 856
rect 24602 734 24802 856
rect 24970 734 25170 856
rect 25338 734 25538 856
rect 25706 734 25906 856
rect 26074 734 26274 856
rect 26442 734 26642 856
rect 26810 734 27010 856
rect 27178 734 27378 856
rect 27546 734 27746 856
rect 27914 734 28114 856
rect 28282 734 28482 856
rect 28650 734 28758 856
rect 28926 734 29126 856
rect 29294 734 29494 856
rect 29662 734 29862 856
rect 30030 734 30230 856
rect 30398 734 30598 856
rect 30766 734 30966 856
rect 31134 734 31334 856
rect 31502 734 31702 856
rect 31870 734 32070 856
rect 32238 734 32438 856
rect 32606 734 32806 856
rect 32974 734 33174 856
rect 33342 734 33542 856
rect 33710 734 33910 856
rect 34078 734 34278 856
rect 34446 734 34646 856
rect 34814 734 35014 856
rect 35182 734 35382 856
rect 35550 734 35750 856
rect 35918 734 36118 856
rect 36286 734 36486 856
rect 36654 734 36854 856
rect 37022 734 37222 856
rect 37390 734 37590 856
rect 37758 734 37958 856
rect 38126 734 38234 856
rect 38402 734 38602 856
rect 38770 734 38970 856
rect 39138 734 39338 856
rect 39506 734 39706 856
rect 39874 734 40074 856
rect 40242 734 40442 856
rect 40610 734 40810 856
rect 40978 734 41178 856
rect 41346 734 41546 856
rect 41714 734 41914 856
rect 42082 734 42282 856
rect 42450 734 42650 856
rect 42818 734 43018 856
rect 43186 734 43386 856
rect 43554 734 43754 856
rect 43922 734 44122 856
rect 44290 734 44490 856
rect 44658 734 44858 856
rect 45026 734 45226 856
rect 45394 734 45594 856
rect 45762 734 45962 856
rect 46130 734 46330 856
rect 46498 734 46698 856
rect 46866 734 47066 856
rect 47234 734 47434 856
rect 47602 734 47710 856
rect 47878 734 48078 856
rect 48246 734 48446 856
rect 48614 734 48814 856
rect 48982 734 49182 856
rect 49350 734 49550 856
rect 49718 734 49918 856
rect 50086 734 50286 856
rect 50454 734 50654 856
rect 50822 734 51022 856
rect 51190 734 51390 856
rect 51558 734 51758 856
rect 51926 734 52126 856
rect 52294 734 52494 856
rect 52662 734 52862 856
rect 53030 734 53230 856
rect 53398 734 53598 856
rect 53766 734 53966 856
rect 54134 734 54334 856
rect 54502 734 54702 856
rect 54870 734 55070 856
rect 55238 734 55438 856
rect 55606 734 55806 856
rect 55974 734 56174 856
rect 56342 734 56542 856
rect 56710 734 56910 856
rect 57078 734 57186 856
rect 57354 734 57554 856
rect 57722 734 57922 856
rect 58090 734 58290 856
rect 58458 734 58658 856
rect 58826 734 59026 856
rect 59194 734 59394 856
rect 59562 734 59762 856
rect 59930 734 60130 856
rect 60298 734 60498 856
rect 60666 734 60866 856
rect 61034 734 61234 856
rect 61402 734 61602 856
rect 61770 734 61970 856
rect 62138 734 62338 856
rect 62506 734 62706 856
rect 62874 734 63074 856
rect 63242 734 63442 856
rect 63610 734 63810 856
rect 63978 734 64178 856
rect 64346 734 64546 856
rect 64714 734 64914 856
rect 65082 734 65282 856
rect 65450 734 65650 856
rect 65818 734 66018 856
rect 66186 734 66386 856
rect 66554 734 66662 856
rect 66830 734 67030 856
rect 67198 734 67398 856
rect 67566 734 67766 856
rect 67934 734 68134 856
rect 68302 734 68502 856
rect 68670 734 68870 856
rect 69038 734 69238 856
rect 69406 734 69606 856
rect 69774 734 69974 856
rect 70142 734 70342 856
rect 70510 734 70710 856
rect 70878 734 71078 856
rect 71246 734 71446 856
rect 71614 734 71814 856
rect 71982 734 72182 856
rect 72350 734 72550 856
rect 72718 734 72918 856
rect 73086 734 73286 856
rect 73454 734 73654 856
rect 73822 734 74022 856
rect 74190 734 74390 856
rect 74558 734 74758 856
rect 74926 734 75126 856
rect 75294 734 75494 856
rect 75662 734 75862 856
rect 76030 734 76138 856
rect 76306 734 76506 856
rect 76674 734 76874 856
rect 77042 734 77242 856
rect 77410 734 77610 856
rect 77778 734 77978 856
rect 78146 734 78346 856
rect 78514 734 78714 856
rect 78882 734 79082 856
rect 79250 734 79450 856
rect 79618 734 79818 856
rect 79986 734 80186 856
rect 80354 734 80554 856
rect 80722 734 80922 856
rect 81090 734 81290 856
rect 81458 734 81658 856
rect 81826 734 82026 856
rect 82194 734 82394 856
rect 82562 734 82762 856
rect 82930 734 83130 856
rect 83298 734 83498 856
rect 83666 734 83866 856
rect 84034 734 84234 856
rect 84402 734 84602 856
rect 84770 734 84970 856
rect 85138 734 85338 856
rect 85506 734 85614 856
rect 85782 734 85982 856
rect 86150 734 86350 856
rect 86518 734 86718 856
rect 86886 734 87086 856
rect 87254 734 87454 856
rect 87622 734 87822 856
rect 87990 734 88190 856
rect 88358 734 88558 856
rect 88726 734 88926 856
rect 89094 734 89294 856
rect 89462 734 89662 856
rect 89830 734 90030 856
rect 90198 734 90398 856
rect 90566 734 90766 856
rect 90934 734 91134 856
rect 91302 734 91502 856
rect 91670 734 91870 856
rect 92038 734 92238 856
rect 92406 734 92606 856
rect 92774 734 92974 856
rect 93142 734 93342 856
rect 93510 734 93710 856
rect 93878 734 94078 856
rect 94246 734 94446 856
rect 94614 734 94814 856
rect 94982 734 95090 856
rect 95258 734 95458 856
rect 95626 734 95826 856
rect 95994 734 96194 856
rect 96362 734 96562 856
rect 96730 734 96930 856
rect 97098 734 97298 856
rect 97466 734 97666 856
rect 97834 734 98034 856
rect 98202 734 98402 856
rect 98570 734 98770 856
rect 98938 734 99138 856
rect 99306 734 99506 856
rect 99674 734 99874 856
rect 100042 734 100242 856
rect 100410 734 100610 856
rect 100778 734 100978 856
rect 101146 734 101346 856
rect 101514 734 101714 856
rect 101882 734 102082 856
rect 102250 734 102450 856
rect 102618 734 102818 856
rect 102986 734 103186 856
rect 103354 734 103554 856
rect 103722 734 103922 856
rect 104090 734 104290 856
rect 104458 734 104566 856
rect 104734 734 104934 856
rect 105102 734 105302 856
rect 105470 734 105670 856
rect 105838 734 106038 856
rect 106206 734 106406 856
rect 106574 734 106774 856
rect 106942 734 107142 856
rect 107310 734 107510 856
rect 107678 734 107878 856
rect 108046 734 108246 856
rect 108414 734 108614 856
rect 108782 734 108982 856
rect 109150 734 109350 856
rect 109518 734 109718 856
rect 109886 734 110086 856
rect 110254 734 110454 856
rect 110622 734 110822 856
rect 110990 734 111190 856
rect 111358 734 111558 856
rect 111726 734 111926 856
rect 112094 734 112294 856
rect 112462 734 112662 856
rect 112830 734 113030 856
rect 113198 734 113398 856
rect 113566 734 113766 856
rect 113934 734 114042 856
rect 114210 734 114410 856
rect 114578 734 114778 856
rect 114946 734 115146 856
rect 115314 734 115514 856
rect 115682 734 115882 856
rect 116050 734 116250 856
rect 116418 734 116618 856
rect 116786 734 116986 856
rect 117154 734 117354 856
rect 117522 734 117722 856
rect 117890 734 118090 856
rect 118258 734 118458 856
rect 118626 734 118826 856
rect 118994 734 119194 856
rect 119362 734 119562 856
rect 119730 734 119930 856
rect 120098 734 120298 856
rect 120466 734 120666 856
rect 120834 734 121034 856
rect 121202 734 121402 856
rect 121570 734 121770 856
rect 121938 734 122138 856
rect 122306 734 122506 856
rect 122674 734 122874 856
rect 123042 734 123242 856
rect 123410 734 123518 856
rect 123686 734 123886 856
rect 124054 734 124254 856
rect 124422 734 124622 856
rect 124790 734 124990 856
rect 125158 734 125358 856
rect 125526 734 125726 856
rect 125894 734 126094 856
rect 126262 734 126462 856
rect 126630 734 126830 856
rect 126998 734 127198 856
rect 127366 734 127566 856
rect 127734 734 127934 856
rect 128102 734 128302 856
rect 128470 734 128670 856
rect 128838 734 129038 856
rect 129206 734 129406 856
rect 129574 734 129774 856
rect 129942 734 130142 856
rect 130310 734 130510 856
rect 130678 734 130878 856
rect 131046 734 131246 856
rect 131414 734 131614 856
rect 131782 734 131982 856
rect 132150 734 132350 856
rect 132518 734 132718 856
rect 132886 734 132994 856
rect 133162 734 133362 856
rect 133530 734 133730 856
rect 133898 734 134098 856
rect 134266 734 134466 856
rect 134634 734 134834 856
rect 135002 734 135202 856
rect 135370 734 135570 856
rect 135738 734 135938 856
rect 136106 734 136306 856
rect 136474 734 136674 856
rect 136842 734 137042 856
rect 137210 734 137410 856
rect 137578 734 137778 856
rect 137946 734 138146 856
rect 138314 734 138514 856
rect 138682 734 138882 856
rect 139050 734 139250 856
rect 139418 734 139618 856
rect 139786 734 139986 856
rect 140154 734 140354 856
rect 140522 734 140722 856
rect 140890 734 141090 856
rect 141258 734 141458 856
rect 141626 734 141826 856
rect 141994 734 142194 856
rect 142362 734 142470 856
rect 142638 734 142838 856
rect 143006 734 143206 856
rect 143374 734 143574 856
rect 143742 734 143942 856
rect 144110 734 144310 856
rect 144478 734 144678 856
rect 144846 734 145046 856
rect 145214 734 145414 856
rect 145582 734 145782 856
rect 145950 734 146150 856
rect 146318 734 146518 856
rect 146686 734 146886 856
rect 147054 734 147254 856
rect 147422 734 147622 856
rect 147790 734 147990 856
rect 148158 734 148358 856
rect 148526 734 148726 856
rect 148894 734 149094 856
rect 149262 734 149462 856
rect 149630 734 149830 856
rect 149998 734 150198 856
rect 150366 734 150566 856
rect 150734 734 150934 856
rect 151102 734 151302 856
rect 151470 734 151670 856
rect 151838 734 151946 856
rect 152114 734 152314 856
rect 152482 734 152682 856
rect 152850 734 153050 856
rect 153218 734 153418 856
rect 153586 734 153786 856
rect 153954 734 154154 856
rect 154322 734 154522 856
rect 154690 734 154890 856
rect 155058 734 155258 856
rect 155426 734 155626 856
rect 155794 734 155994 856
rect 156162 734 156362 856
rect 156530 734 156730 856
rect 156898 734 157098 856
rect 157266 734 157466 856
rect 157634 734 157834 856
rect 158002 734 158202 856
rect 158370 734 158570 856
rect 158738 734 158938 856
rect 159106 734 159306 856
rect 159474 734 159674 856
rect 159842 734 160042 856
rect 160210 734 160410 856
rect 160578 734 160778 856
rect 160946 734 161146 856
rect 161314 734 161422 856
rect 161590 734 161790 856
rect 161958 734 162158 856
rect 162326 734 162526 856
rect 162694 734 162894 856
rect 163062 734 163262 856
rect 163430 734 163630 856
rect 163798 734 163998 856
rect 164166 734 164366 856
rect 164534 734 164734 856
rect 164902 734 165102 856
rect 165270 734 165470 856
rect 165638 734 165838 856
rect 166006 734 166206 856
rect 166374 734 166574 856
rect 166742 734 166942 856
rect 167110 734 167310 856
rect 167478 734 167678 856
rect 167846 734 168046 856
rect 168214 734 168414 856
rect 168582 734 168782 856
rect 168950 734 169150 856
rect 169318 734 169518 856
rect 169686 734 169886 856
rect 170054 734 170254 856
rect 170422 734 170622 856
rect 170790 734 170898 856
rect 171066 734 171266 856
rect 171434 734 171634 856
rect 171802 734 172002 856
rect 172170 734 172370 856
rect 172538 734 172738 856
rect 172906 734 173106 856
rect 173274 734 173474 856
rect 173642 734 173842 856
rect 174010 734 174210 856
rect 174378 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175314 856
rect 175482 734 175682 856
rect 175850 734 176050 856
rect 176218 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178186 856
<< metal3 >>
rect 179200 113840 180000 113960
rect 0 111392 800 111512
rect 179200 101872 180000 101992
rect 0 94256 800 94376
rect 179200 89904 180000 90024
rect 179200 77936 180000 78056
rect 0 77120 800 77240
rect 179200 65968 180000 66088
rect 0 59984 800 60104
rect 179200 53864 180000 53984
rect 0 42848 800 42968
rect 179200 41896 180000 42016
rect 179200 29928 180000 30048
rect 0 25712 800 25832
rect 179200 17960 180000 18080
rect 0 8576 800 8696
rect 179200 5992 180000 6112
<< obsm3 >>
rect 800 114040 179200 117741
rect 800 113760 179120 114040
rect 800 111592 179200 113760
rect 880 111312 179200 111592
rect 800 102072 179200 111312
rect 800 101792 179120 102072
rect 800 94456 179200 101792
rect 880 94176 179200 94456
rect 800 90104 179200 94176
rect 800 89824 179120 90104
rect 800 78136 179200 89824
rect 800 77856 179120 78136
rect 800 77320 179200 77856
rect 880 77040 179200 77320
rect 800 66168 179200 77040
rect 800 65888 179120 66168
rect 800 60184 179200 65888
rect 880 59904 179200 60184
rect 800 54064 179200 59904
rect 800 53784 179120 54064
rect 800 43048 179200 53784
rect 880 42768 179200 43048
rect 800 42096 179200 42768
rect 800 41816 179120 42096
rect 800 30128 179200 41816
rect 800 29848 179120 30128
rect 800 25912 179200 29848
rect 880 25632 179200 25912
rect 800 18160 179200 25632
rect 800 17880 179120 18160
rect 800 8776 179200 17880
rect 880 8496 179200 8776
rect 800 6192 179200 8496
rect 800 5912 179120 6192
rect 800 2143 179200 5912
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 63171 110331 65568 117605
rect 66048 110331 80928 117605
rect 81408 110331 96173 117605
<< labels >>
rlabel metal3 s 0 8576 800 8696 6 active
port 1 nsew signal input
rlabel metal3 s 179200 17960 180000 18080 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal2 s 169298 119200 169354 120000 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal2 s 170770 119200 170826 120000 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal3 s 179200 65968 180000 66088 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 0 77120 800 77240 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal3 s 0 94256 800 94376 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal3 s 179200 77936 180000 78056 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal2 s 172150 119200 172206 120000 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal2 s 173530 119200 173586 120000 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal2 s 162214 119200 162270 120000 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 175002 119200 175058 120000 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal3 s 179200 89904 180000 90024 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 0 111392 800 111512 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 176382 119200 176438 120000 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 177854 119200 177910 120000 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 179200 101872 180000 101992 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal3 s 179200 113840 180000 113960 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 179200 41896 180000 42016 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 165066 119200 165122 120000 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 179200 53864 180000 53984 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal2 s 166446 119200 166502 120000 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 0 42848 800 42968 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal2 s 167918 119200 167974 120000 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 43166 119200 43222 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 47398 119200 47454 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 51630 119200 51686 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 55862 119200 55918 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 60186 119200 60242 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 64418 119200 64474 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 68650 119200 68706 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 72882 119200 72938 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 77206 119200 77262 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 81438 119200 81494 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 4894 119200 4950 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 85670 119200 85726 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 94226 119200 94282 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 98458 119200 98514 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 102690 119200 102746 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 111154 119200 111210 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 115478 119200 115534 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 119710 119200 119766 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 123942 119200 123998 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9126 119200 9182 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 128174 119200 128230 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 132498 119200 132554 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 136730 119200 136786 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 140962 119200 141018 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 145194 119200 145250 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 149426 119200 149482 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 153750 119200 153806 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 157982 119200 158038 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 13358 119200 13414 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 17590 119200 17646 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 21914 119200 21970 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 26146 119200 26202 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 30378 119200 30434 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 34610 119200 34666 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 38934 119200 38990 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2042 119200 2098 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 48778 119200 48834 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 53102 119200 53158 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 57334 119200 57390 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 61566 119200 61622 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 65798 119200 65854 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 70122 119200 70178 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 74354 119200 74410 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 82818 119200 82874 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6274 119200 6330 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 91374 119200 91430 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 95606 119200 95662 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 99838 119200 99894 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 104070 119200 104126 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 108394 119200 108450 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 116858 119200 116914 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 121090 119200 121146 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 125414 119200 125470 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 10506 119200 10562 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 129646 119200 129702 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 133878 119200 133934 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 138110 119200 138166 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 142342 119200 142398 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 146666 119200 146722 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 150898 119200 150954 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 155130 119200 155186 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 159362 119200 159418 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 14830 119200 14886 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 19062 119200 19118 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 23294 119200 23350 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 27526 119200 27582 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 31850 119200 31906 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 36082 119200 36138 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 40314 119200 40370 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3422 119200 3478 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 46018 119200 46074 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 50250 119200 50306 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 54482 119200 54538 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 58714 119200 58770 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 63038 119200 63094 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 67270 119200 67326 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 79966 119200 80022 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 84290 119200 84346 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 7746 119200 7802 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 101310 119200 101366 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 105542 119200 105598 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 109774 119200 109830 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 114006 119200 114062 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 122562 119200 122618 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 126794 119200 126850 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 11978 119200 12034 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 131026 119200 131082 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 135258 119200 135314 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 139582 119200 139638 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 143814 119200 143870 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 148046 119200 148102 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 152278 119200 152334 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 156602 119200 156658 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 160834 119200 160890 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 20442 119200 20498 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 24674 119200 24730 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 33230 119200 33286 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 37462 119200 37518 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 41694 119200 41750 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 154946 0 155002 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 157154 0 157210 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 165894 0 165950 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 168102 0 168158 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 129830 0 129886 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 140778 0 140834 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 145102 0 145158 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 123574 0 123630 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 179200 5992 180000 6112 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 user_irq[0]
port 530 nsew signal output
rlabel metal3 s 179200 29928 180000 30048 6 user_irq[1]
port 531 nsew signal output
rlabel metal2 s 163686 119200 163742 120000 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8271392
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_7.magic.gds
string GDS_START 295056
<< end >>

