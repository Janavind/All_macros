magic
tech sky130A
magscale 1 2
timestamp 1653776126
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118380
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9678 119200 9734 120000
rect 11150 119200 11206 120000
rect 12622 119200 12678 120000
rect 14094 119200 14150 120000
rect 15566 119200 15622 120000
rect 17038 119200 17094 120000
rect 18602 119200 18658 120000
rect 20074 119200 20130 120000
rect 21546 119200 21602 120000
rect 23018 119200 23074 120000
rect 24490 119200 24546 120000
rect 25962 119200 26018 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30470 119200 30526 120000
rect 31942 119200 31998 120000
rect 33414 119200 33470 120000
rect 34886 119200 34942 120000
rect 36450 119200 36506 120000
rect 37922 119200 37978 120000
rect 39394 119200 39450 120000
rect 40866 119200 40922 120000
rect 42338 119200 42394 120000
rect 43902 119200 43958 120000
rect 45374 119200 45430 120000
rect 46846 119200 46902 120000
rect 48318 119200 48374 120000
rect 49790 119200 49846 120000
rect 51262 119200 51318 120000
rect 52826 119200 52882 120000
rect 54298 119200 54354 120000
rect 55770 119200 55826 120000
rect 57242 119200 57298 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61750 119200 61806 120000
rect 63222 119200 63278 120000
rect 64694 119200 64750 120000
rect 66166 119200 66222 120000
rect 67638 119200 67694 120000
rect 69110 119200 69166 120000
rect 70674 119200 70730 120000
rect 72146 119200 72202 120000
rect 73618 119200 73674 120000
rect 75090 119200 75146 120000
rect 76562 119200 76618 120000
rect 78126 119200 78182 120000
rect 79598 119200 79654 120000
rect 81070 119200 81126 120000
rect 82542 119200 82598 120000
rect 84014 119200 84070 120000
rect 85486 119200 85542 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89994 119200 90050 120000
rect 91466 119200 91522 120000
rect 92938 119200 92994 120000
rect 94410 119200 94466 120000
rect 95974 119200 96030 120000
rect 97446 119200 97502 120000
rect 98918 119200 98974 120000
rect 100390 119200 100446 120000
rect 101862 119200 101918 120000
rect 103334 119200 103390 120000
rect 104898 119200 104954 120000
rect 106370 119200 106426 120000
rect 107842 119200 107898 120000
rect 109314 119200 109370 120000
rect 110786 119200 110842 120000
rect 112350 119200 112406 120000
rect 113822 119200 113878 120000
rect 115294 119200 115350 120000
rect 116766 119200 116822 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121274 119200 121330 120000
rect 122746 119200 122802 120000
rect 124218 119200 124274 120000
rect 125690 119200 125746 120000
rect 127162 119200 127218 120000
rect 128634 119200 128690 120000
rect 130198 119200 130254 120000
rect 131670 119200 131726 120000
rect 133142 119200 133198 120000
rect 134614 119200 134670 120000
rect 136086 119200 136142 120000
rect 137558 119200 137614 120000
rect 139122 119200 139178 120000
rect 140594 119200 140650 120000
rect 142066 119200 142122 120000
rect 143538 119200 143594 120000
rect 145010 119200 145066 120000
rect 146574 119200 146630 120000
rect 148046 119200 148102 120000
rect 149518 119200 149574 120000
rect 150990 119200 151046 120000
rect 152462 119200 152518 120000
rect 153934 119200 153990 120000
rect 155498 119200 155554 120000
rect 156970 119200 157026 120000
rect 158442 119200 158498 120000
rect 159914 119200 159970 120000
rect 161386 119200 161442 120000
rect 162858 119200 162914 120000
rect 164422 119200 164478 120000
rect 165894 119200 165950 120000
rect 167366 119200 167422 120000
rect 168838 119200 168894 120000
rect 170310 119200 170366 120000
rect 171782 119200 171838 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31298 0 31354 800
rect 31666 0 31722 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35622 0 35678 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37462 0 37518 800
rect 37830 0 37886 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42154 0 42210 800
rect 42522 0 42578 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46202 0 46258 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55954 0 56010 800
rect 56322 0 56378 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57426 0 57482 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62486 0 62542 800
rect 62854 0 62910 800
rect 63222 0 63278 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81346 0 81402 800
rect 81714 0 81770 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 93030 0 93086 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95882 0 95938 800
rect 96250 0 96306 800
rect 96618 0 96674 800
rect 96986 0 97042 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98458 0 98514 800
rect 98826 0 98882 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108946 0 109002 800
rect 109314 0 109370 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116950 0 117006 800
rect 117318 0 117374 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123850 0 123906 800
rect 124218 0 124274 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126426 0 126482 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129278 0 129334 800
rect 129646 0 129702 800
rect 130014 0 130070 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133970 0 134026 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140134 0 140190 800
rect 140502 0 140558 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 141974 0 142030 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146022 0 146078 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147770 0 147826 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151450 0 151506 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153566 0 153622 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155406 0 155462 800
rect 155774 0 155830 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156878 0 156934 800
rect 157246 0 157302 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161938 0 161994 800
rect 162306 0 162362 800
rect 162674 0 162730 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163778 0 163834 800
rect 164146 0 164202 800
rect 164514 0 164570 800
rect 164882 0 164938 800
rect 165250 0 165306 800
rect 165618 0 165674 800
rect 165986 0 166042 800
rect 166354 0 166410 800
rect 166722 0 166778 800
rect 166998 0 167054 800
rect 167366 0 167422 800
rect 167734 0 167790 800
rect 168102 0 168158 800
rect 168470 0 168526 800
rect 168838 0 168894 800
rect 169206 0 169262 800
rect 169574 0 169630 800
rect 169942 0 169998 800
rect 170310 0 170366 800
rect 170678 0 170734 800
rect 171046 0 171102 800
rect 171414 0 171470 800
rect 171782 0 171838 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173254 0 173310 800
rect 173530 0 173586 800
rect 173898 0 173954 800
rect 174266 0 174322 800
rect 174634 0 174690 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176106 0 176162 800
rect 176474 0 176530 800
rect 176842 0 176898 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6586 119354
rect 6754 119144 8058 119354
rect 8226 119144 9622 119354
rect 9790 119144 11094 119354
rect 11262 119144 12566 119354
rect 12734 119144 14038 119354
rect 14206 119144 15510 119354
rect 15678 119144 16982 119354
rect 17150 119144 18546 119354
rect 18714 119144 20018 119354
rect 20186 119144 21490 119354
rect 21658 119144 22962 119354
rect 23130 119144 24434 119354
rect 24602 119144 25906 119354
rect 26074 119144 27470 119354
rect 27638 119144 28942 119354
rect 29110 119144 30414 119354
rect 30582 119144 31886 119354
rect 32054 119144 33358 119354
rect 33526 119144 34830 119354
rect 34998 119144 36394 119354
rect 36562 119144 37866 119354
rect 38034 119144 39338 119354
rect 39506 119144 40810 119354
rect 40978 119144 42282 119354
rect 42450 119144 43846 119354
rect 44014 119144 45318 119354
rect 45486 119144 46790 119354
rect 46958 119144 48262 119354
rect 48430 119144 49734 119354
rect 49902 119144 51206 119354
rect 51374 119144 52770 119354
rect 52938 119144 54242 119354
rect 54410 119144 55714 119354
rect 55882 119144 57186 119354
rect 57354 119144 58658 119354
rect 58826 119144 60130 119354
rect 60298 119144 61694 119354
rect 61862 119144 63166 119354
rect 63334 119144 64638 119354
rect 64806 119144 66110 119354
rect 66278 119144 67582 119354
rect 67750 119144 69054 119354
rect 69222 119144 70618 119354
rect 70786 119144 72090 119354
rect 72258 119144 73562 119354
rect 73730 119144 75034 119354
rect 75202 119144 76506 119354
rect 76674 119144 78070 119354
rect 78238 119144 79542 119354
rect 79710 119144 81014 119354
rect 81182 119144 82486 119354
rect 82654 119144 83958 119354
rect 84126 119144 85430 119354
rect 85598 119144 86994 119354
rect 87162 119144 88466 119354
rect 88634 119144 89938 119354
rect 90106 119144 91410 119354
rect 91578 119144 92882 119354
rect 93050 119144 94354 119354
rect 94522 119144 95918 119354
rect 96086 119144 97390 119354
rect 97558 119144 98862 119354
rect 99030 119144 100334 119354
rect 100502 119144 101806 119354
rect 101974 119144 103278 119354
rect 103446 119144 104842 119354
rect 105010 119144 106314 119354
rect 106482 119144 107786 119354
rect 107954 119144 109258 119354
rect 109426 119144 110730 119354
rect 110898 119144 112294 119354
rect 112462 119144 113766 119354
rect 113934 119144 115238 119354
rect 115406 119144 116710 119354
rect 116878 119144 118182 119354
rect 118350 119144 119654 119354
rect 119822 119144 121218 119354
rect 121386 119144 122690 119354
rect 122858 119144 124162 119354
rect 124330 119144 125634 119354
rect 125802 119144 127106 119354
rect 127274 119144 128578 119354
rect 128746 119144 130142 119354
rect 130310 119144 131614 119354
rect 131782 119144 133086 119354
rect 133254 119144 134558 119354
rect 134726 119144 136030 119354
rect 136198 119144 137502 119354
rect 137670 119144 139066 119354
rect 139234 119144 140538 119354
rect 140706 119144 142010 119354
rect 142178 119144 143482 119354
rect 143650 119144 144954 119354
rect 145122 119144 146518 119354
rect 146686 119144 147990 119354
rect 148158 119144 149462 119354
rect 149630 119144 150934 119354
rect 151102 119144 152406 119354
rect 152574 119144 153878 119354
rect 154046 119144 155442 119354
rect 155610 119144 156914 119354
rect 157082 119144 158386 119354
rect 158554 119144 159858 119354
rect 160026 119144 161330 119354
rect 161498 119144 162802 119354
rect 162970 119144 164366 119354
rect 164534 119144 165838 119354
rect 166006 119144 167310 119354
rect 167478 119144 168782 119354
rect 168950 119144 170254 119354
rect 170422 119144 171726 119354
rect 171894 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178368 119354
rect 756 856 178368 119144
rect 866 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6862 856
rect 7030 734 7230 856
rect 7398 734 7598 856
rect 7766 734 7966 856
rect 8134 734 8334 856
rect 8502 734 8702 856
rect 8870 734 9070 856
rect 9238 734 9438 856
rect 9606 734 9806 856
rect 9974 734 10174 856
rect 10342 734 10542 856
rect 10710 734 10910 856
rect 11078 734 11278 856
rect 11446 734 11646 856
rect 11814 734 12014 856
rect 12182 734 12382 856
rect 12550 734 12750 856
rect 12918 734 13118 856
rect 13286 734 13394 856
rect 13562 734 13762 856
rect 13930 734 14130 856
rect 14298 734 14498 856
rect 14666 734 14866 856
rect 15034 734 15234 856
rect 15402 734 15602 856
rect 15770 734 15970 856
rect 16138 734 16338 856
rect 16506 734 16706 856
rect 16874 734 17074 856
rect 17242 734 17442 856
rect 17610 734 17810 856
rect 17978 734 18178 856
rect 18346 734 18546 856
rect 18714 734 18914 856
rect 19082 734 19282 856
rect 19450 734 19650 856
rect 19818 734 20018 856
rect 20186 734 20294 856
rect 20462 734 20662 856
rect 20830 734 21030 856
rect 21198 734 21398 856
rect 21566 734 21766 856
rect 21934 734 22134 856
rect 22302 734 22502 856
rect 22670 734 22870 856
rect 23038 734 23238 856
rect 23406 734 23606 856
rect 23774 734 23974 856
rect 24142 734 24342 856
rect 24510 734 24710 856
rect 24878 734 25078 856
rect 25246 734 25446 856
rect 25614 734 25814 856
rect 25982 734 26182 856
rect 26350 734 26550 856
rect 26718 734 26826 856
rect 26994 734 27194 856
rect 27362 734 27562 856
rect 27730 734 27930 856
rect 28098 734 28298 856
rect 28466 734 28666 856
rect 28834 734 29034 856
rect 29202 734 29402 856
rect 29570 734 29770 856
rect 29938 734 30138 856
rect 30306 734 30506 856
rect 30674 734 30874 856
rect 31042 734 31242 856
rect 31410 734 31610 856
rect 31778 734 31978 856
rect 32146 734 32346 856
rect 32514 734 32714 856
rect 32882 734 33082 856
rect 33250 734 33358 856
rect 33526 734 33726 856
rect 33894 734 34094 856
rect 34262 734 34462 856
rect 34630 734 34830 856
rect 34998 734 35198 856
rect 35366 734 35566 856
rect 35734 734 35934 856
rect 36102 734 36302 856
rect 36470 734 36670 856
rect 36838 734 37038 856
rect 37206 734 37406 856
rect 37574 734 37774 856
rect 37942 734 38142 856
rect 38310 734 38510 856
rect 38678 734 38878 856
rect 39046 734 39246 856
rect 39414 734 39614 856
rect 39782 734 39982 856
rect 40150 734 40258 856
rect 40426 734 40626 856
rect 40794 734 40994 856
rect 41162 734 41362 856
rect 41530 734 41730 856
rect 41898 734 42098 856
rect 42266 734 42466 856
rect 42634 734 42834 856
rect 43002 734 43202 856
rect 43370 734 43570 856
rect 43738 734 43938 856
rect 44106 734 44306 856
rect 44474 734 44674 856
rect 44842 734 45042 856
rect 45210 734 45410 856
rect 45578 734 45778 856
rect 45946 734 46146 856
rect 46314 734 46514 856
rect 46682 734 46790 856
rect 46958 734 47158 856
rect 47326 734 47526 856
rect 47694 734 47894 856
rect 48062 734 48262 856
rect 48430 734 48630 856
rect 48798 734 48998 856
rect 49166 734 49366 856
rect 49534 734 49734 856
rect 49902 734 50102 856
rect 50270 734 50470 856
rect 50638 734 50838 856
rect 51006 734 51206 856
rect 51374 734 51574 856
rect 51742 734 51942 856
rect 52110 734 52310 856
rect 52478 734 52678 856
rect 52846 734 53046 856
rect 53214 734 53322 856
rect 53490 734 53690 856
rect 53858 734 54058 856
rect 54226 734 54426 856
rect 54594 734 54794 856
rect 54962 734 55162 856
rect 55330 734 55530 856
rect 55698 734 55898 856
rect 56066 734 56266 856
rect 56434 734 56634 856
rect 56802 734 57002 856
rect 57170 734 57370 856
rect 57538 734 57738 856
rect 57906 734 58106 856
rect 58274 734 58474 856
rect 58642 734 58842 856
rect 59010 734 59210 856
rect 59378 734 59578 856
rect 59746 734 59946 856
rect 60114 734 60222 856
rect 60390 734 60590 856
rect 60758 734 60958 856
rect 61126 734 61326 856
rect 61494 734 61694 856
rect 61862 734 62062 856
rect 62230 734 62430 856
rect 62598 734 62798 856
rect 62966 734 63166 856
rect 63334 734 63534 856
rect 63702 734 63902 856
rect 64070 734 64270 856
rect 64438 734 64638 856
rect 64806 734 65006 856
rect 65174 734 65374 856
rect 65542 734 65742 856
rect 65910 734 66110 856
rect 66278 734 66478 856
rect 66646 734 66754 856
rect 66922 734 67122 856
rect 67290 734 67490 856
rect 67658 734 67858 856
rect 68026 734 68226 856
rect 68394 734 68594 856
rect 68762 734 68962 856
rect 69130 734 69330 856
rect 69498 734 69698 856
rect 69866 734 70066 856
rect 70234 734 70434 856
rect 70602 734 70802 856
rect 70970 734 71170 856
rect 71338 734 71538 856
rect 71706 734 71906 856
rect 72074 734 72274 856
rect 72442 734 72642 856
rect 72810 734 73010 856
rect 73178 734 73378 856
rect 73546 734 73654 856
rect 73822 734 74022 856
rect 74190 734 74390 856
rect 74558 734 74758 856
rect 74926 734 75126 856
rect 75294 734 75494 856
rect 75662 734 75862 856
rect 76030 734 76230 856
rect 76398 734 76598 856
rect 76766 734 76966 856
rect 77134 734 77334 856
rect 77502 734 77702 856
rect 77870 734 78070 856
rect 78238 734 78438 856
rect 78606 734 78806 856
rect 78974 734 79174 856
rect 79342 734 79542 856
rect 79710 734 79910 856
rect 80078 734 80186 856
rect 80354 734 80554 856
rect 80722 734 80922 856
rect 81090 734 81290 856
rect 81458 734 81658 856
rect 81826 734 82026 856
rect 82194 734 82394 856
rect 82562 734 82762 856
rect 82930 734 83130 856
rect 83298 734 83498 856
rect 83666 734 83866 856
rect 84034 734 84234 856
rect 84402 734 84602 856
rect 84770 734 84970 856
rect 85138 734 85338 856
rect 85506 734 85706 856
rect 85874 734 86074 856
rect 86242 734 86442 856
rect 86610 734 86718 856
rect 86886 734 87086 856
rect 87254 734 87454 856
rect 87622 734 87822 856
rect 87990 734 88190 856
rect 88358 734 88558 856
rect 88726 734 88926 856
rect 89094 734 89294 856
rect 89462 734 89662 856
rect 89830 734 90030 856
rect 90198 734 90398 856
rect 90566 734 90766 856
rect 90934 734 91134 856
rect 91302 734 91502 856
rect 91670 734 91870 856
rect 92038 734 92238 856
rect 92406 734 92606 856
rect 92774 734 92974 856
rect 93142 734 93342 856
rect 93510 734 93618 856
rect 93786 734 93986 856
rect 94154 734 94354 856
rect 94522 734 94722 856
rect 94890 734 95090 856
rect 95258 734 95458 856
rect 95626 734 95826 856
rect 95994 734 96194 856
rect 96362 734 96562 856
rect 96730 734 96930 856
rect 97098 734 97298 856
rect 97466 734 97666 856
rect 97834 734 98034 856
rect 98202 734 98402 856
rect 98570 734 98770 856
rect 98938 734 99138 856
rect 99306 734 99506 856
rect 99674 734 99874 856
rect 100042 734 100150 856
rect 100318 734 100518 856
rect 100686 734 100886 856
rect 101054 734 101254 856
rect 101422 734 101622 856
rect 101790 734 101990 856
rect 102158 734 102358 856
rect 102526 734 102726 856
rect 102894 734 103094 856
rect 103262 734 103462 856
rect 103630 734 103830 856
rect 103998 734 104198 856
rect 104366 734 104566 856
rect 104734 734 104934 856
rect 105102 734 105302 856
rect 105470 734 105670 856
rect 105838 734 106038 856
rect 106206 734 106406 856
rect 106574 734 106682 856
rect 106850 734 107050 856
rect 107218 734 107418 856
rect 107586 734 107786 856
rect 107954 734 108154 856
rect 108322 734 108522 856
rect 108690 734 108890 856
rect 109058 734 109258 856
rect 109426 734 109626 856
rect 109794 734 109994 856
rect 110162 734 110362 856
rect 110530 734 110730 856
rect 110898 734 111098 856
rect 111266 734 111466 856
rect 111634 734 111834 856
rect 112002 734 112202 856
rect 112370 734 112570 856
rect 112738 734 112938 856
rect 113106 734 113306 856
rect 113474 734 113582 856
rect 113750 734 113950 856
rect 114118 734 114318 856
rect 114486 734 114686 856
rect 114854 734 115054 856
rect 115222 734 115422 856
rect 115590 734 115790 856
rect 115958 734 116158 856
rect 116326 734 116526 856
rect 116694 734 116894 856
rect 117062 734 117262 856
rect 117430 734 117630 856
rect 117798 734 117998 856
rect 118166 734 118366 856
rect 118534 734 118734 856
rect 118902 734 119102 856
rect 119270 734 119470 856
rect 119638 734 119838 856
rect 120006 734 120114 856
rect 120282 734 120482 856
rect 120650 734 120850 856
rect 121018 734 121218 856
rect 121386 734 121586 856
rect 121754 734 121954 856
rect 122122 734 122322 856
rect 122490 734 122690 856
rect 122858 734 123058 856
rect 123226 734 123426 856
rect 123594 734 123794 856
rect 123962 734 124162 856
rect 124330 734 124530 856
rect 124698 734 124898 856
rect 125066 734 125266 856
rect 125434 734 125634 856
rect 125802 734 126002 856
rect 126170 734 126370 856
rect 126538 734 126738 856
rect 126906 734 127014 856
rect 127182 734 127382 856
rect 127550 734 127750 856
rect 127918 734 128118 856
rect 128286 734 128486 856
rect 128654 734 128854 856
rect 129022 734 129222 856
rect 129390 734 129590 856
rect 129758 734 129958 856
rect 130126 734 130326 856
rect 130494 734 130694 856
rect 130862 734 131062 856
rect 131230 734 131430 856
rect 131598 734 131798 856
rect 131966 734 132166 856
rect 132334 734 132534 856
rect 132702 734 132902 856
rect 133070 734 133270 856
rect 133438 734 133546 856
rect 133714 734 133914 856
rect 134082 734 134282 856
rect 134450 734 134650 856
rect 134818 734 135018 856
rect 135186 734 135386 856
rect 135554 734 135754 856
rect 135922 734 136122 856
rect 136290 734 136490 856
rect 136658 734 136858 856
rect 137026 734 137226 856
rect 137394 734 137594 856
rect 137762 734 137962 856
rect 138130 734 138330 856
rect 138498 734 138698 856
rect 138866 734 139066 856
rect 139234 734 139434 856
rect 139602 734 139802 856
rect 139970 734 140078 856
rect 140246 734 140446 856
rect 140614 734 140814 856
rect 140982 734 141182 856
rect 141350 734 141550 856
rect 141718 734 141918 856
rect 142086 734 142286 856
rect 142454 734 142654 856
rect 142822 734 143022 856
rect 143190 734 143390 856
rect 143558 734 143758 856
rect 143926 734 144126 856
rect 144294 734 144494 856
rect 144662 734 144862 856
rect 145030 734 145230 856
rect 145398 734 145598 856
rect 145766 734 145966 856
rect 146134 734 146334 856
rect 146502 734 146702 856
rect 146870 734 146978 856
rect 147146 734 147346 856
rect 147514 734 147714 856
rect 147882 734 148082 856
rect 148250 734 148450 856
rect 148618 734 148818 856
rect 148986 734 149186 856
rect 149354 734 149554 856
rect 149722 734 149922 856
rect 150090 734 150290 856
rect 150458 734 150658 856
rect 150826 734 151026 856
rect 151194 734 151394 856
rect 151562 734 151762 856
rect 151930 734 152130 856
rect 152298 734 152498 856
rect 152666 734 152866 856
rect 153034 734 153234 856
rect 153402 734 153510 856
rect 153678 734 153878 856
rect 154046 734 154246 856
rect 154414 734 154614 856
rect 154782 734 154982 856
rect 155150 734 155350 856
rect 155518 734 155718 856
rect 155886 734 156086 856
rect 156254 734 156454 856
rect 156622 734 156822 856
rect 156990 734 157190 856
rect 157358 734 157558 856
rect 157726 734 157926 856
rect 158094 734 158294 856
rect 158462 734 158662 856
rect 158830 734 159030 856
rect 159198 734 159398 856
rect 159566 734 159766 856
rect 159934 734 160042 856
rect 160210 734 160410 856
rect 160578 734 160778 856
rect 160946 734 161146 856
rect 161314 734 161514 856
rect 161682 734 161882 856
rect 162050 734 162250 856
rect 162418 734 162618 856
rect 162786 734 162986 856
rect 163154 734 163354 856
rect 163522 734 163722 856
rect 163890 734 164090 856
rect 164258 734 164458 856
rect 164626 734 164826 856
rect 164994 734 165194 856
rect 165362 734 165562 856
rect 165730 734 165930 856
rect 166098 734 166298 856
rect 166466 734 166666 856
rect 166834 734 166942 856
rect 167110 734 167310 856
rect 167478 734 167678 856
rect 167846 734 168046 856
rect 168214 734 168414 856
rect 168582 734 168782 856
rect 168950 734 169150 856
rect 169318 734 169518 856
rect 169686 734 169886 856
rect 170054 734 170254 856
rect 170422 734 170622 856
rect 170790 734 170990 856
rect 171158 734 171358 856
rect 171526 734 171726 856
rect 171894 734 172094 856
rect 172262 734 172462 856
rect 172630 734 172830 856
rect 172998 734 173198 856
rect 173366 734 173474 856
rect 173642 734 173842 856
rect 174010 734 174210 856
rect 174378 734 174578 856
rect 174746 734 174946 856
rect 175114 734 175314 856
rect 175482 734 175682 856
rect 175850 734 176050 856
rect 176218 734 176418 856
rect 176586 734 176786 856
rect 176954 734 177154 856
rect 177322 734 177522 856
rect 177690 734 177890 856
rect 178058 734 178258 856
<< metal3 >>
rect 179200 115608 180000 115728
rect 0 111392 800 111512
rect 179200 107040 180000 107160
rect 179200 98472 180000 98592
rect 0 94256 800 94376
rect 179200 89904 180000 90024
rect 179200 81336 180000 81456
rect 0 77120 800 77240
rect 179200 72768 180000 72888
rect 179200 64200 180000 64320
rect 0 59984 800 60104
rect 179200 55632 180000 55752
rect 179200 47064 180000 47184
rect 0 42848 800 42968
rect 179200 38496 180000 38616
rect 179200 29928 180000 30048
rect 0 25712 800 25832
rect 179200 21360 180000 21480
rect 179200 12792 180000 12912
rect 0 8576 800 8696
rect 179200 4224 180000 4344
<< obsm3 >>
rect 1669 115808 179200 118149
rect 1669 115528 179120 115808
rect 1669 107240 179200 115528
rect 1669 106960 179120 107240
rect 1669 98672 179200 106960
rect 1669 98392 179120 98672
rect 1669 90104 179200 98392
rect 1669 89824 179120 90104
rect 1669 81536 179200 89824
rect 1669 81256 179120 81536
rect 1669 72968 179200 81256
rect 1669 72688 179120 72968
rect 1669 64400 179200 72688
rect 1669 64120 179120 64400
rect 1669 55832 179200 64120
rect 1669 55552 179120 55832
rect 1669 47264 179200 55552
rect 1669 46984 179120 47264
rect 1669 38696 179200 46984
rect 1669 38416 179120 38696
rect 1669 30128 179200 38416
rect 1669 29848 179120 30128
rect 1669 21560 179200 29848
rect 1669 21280 179120 21560
rect 1669 12992 179200 21280
rect 1669 12712 179120 12992
rect 1669 4424 179200 12712
rect 1669 4144 179120 4424
rect 1669 2143 179200 4144
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 67587 117632 96909 118013
rect 67587 110331 80928 117632
rect 81408 110331 96288 117632
rect 96768 110331 96909 117632
<< labels >>
rlabel metal2 s 170310 119200 170366 120000 6 active
port 1 nsew signal input
rlabel metal3 s 179200 4224 180000 4344 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 179200 55632 180000 55752 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal3 s 179200 64200 180000 64320 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 179200 72768 180000 72888 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 179200 81336 180000 81456 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal3 s 0 77120 800 77240 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 179200 89904 180000 90024 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 179200 21360 180000 21480 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal3 s 179200 98472 180000 98592 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 179200 107040 180000 107160 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal3 s 0 94256 800 94376 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal3 s 179200 115608 180000 115728 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 0 111392 800 111512 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 179200 29928 180000 30048 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 179200 38496 180000 38616 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 0 8576 800 8696 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 0 25712 800 25832 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 0 42848 800 42968 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 179200 47064 180000 47184 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 45374 119200 45430 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 49790 119200 49846 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 54298 119200 54354 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 58714 119200 58770 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 63222 119200 63278 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 67638 119200 67694 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 76562 119200 76618 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 81070 119200 81126 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 85486 119200 85542 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 89994 119200 90050 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 94410 119200 94466 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 98918 119200 98974 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 103334 119200 103390 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 107842 119200 107898 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 116766 119200 116822 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 121274 119200 121330 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 125690 119200 125746 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 130198 119200 130254 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 148046 119200 148102 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 152462 119200 152518 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 156970 119200 157026 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 161386 119200 161442 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 165894 119200 165950 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 14094 119200 14150 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18602 119200 18658 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 23018 119200 23074 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 27526 119200 27582 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31942 119200 31998 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 36450 119200 36506 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 40866 119200 40922 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 46846 119200 46902 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 60186 119200 60242 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 69110 119200 69166 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 73618 119200 73674 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 95974 119200 96030 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 100390 119200 100446 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 104898 119200 104954 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 109314 119200 109370 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 113822 119200 113878 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 122746 119200 122802 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 127162 119200 127218 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 131670 119200 131726 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 11150 119200 11206 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 136086 119200 136142 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 140594 119200 140650 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 145010 119200 145066 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 149518 119200 149574 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 153934 119200 153990 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 158442 119200 158498 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 162858 119200 162914 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 167366 119200 167422 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15566 119200 15622 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24490 119200 24546 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 33414 119200 33470 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 37922 119200 37978 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 42338 119200 42394 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 48318 119200 48374 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 57242 119200 57298 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 61750 119200 61806 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 66166 119200 66222 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 84014 119200 84070 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 92938 119200 92994 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 97446 119200 97502 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 101862 119200 101918 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 106370 119200 106426 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 110786 119200 110842 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 115294 119200 115350 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 119710 119200 119766 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 128634 119200 128690 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 133142 119200 133198 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12622 119200 12678 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 137558 119200 137614 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 142066 119200 142122 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 146574 119200 146630 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 150990 119200 151046 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 155498 119200 155554 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 159914 119200 159970 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 164422 119200 164478 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 168838 119200 168894 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 17038 119200 17094 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21546 119200 21602 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25962 119200 26018 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 43902 119200 43958 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 171414 0 171470 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 165250 0 165306 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 171782 0 171838 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 176106 0 176162 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 78126 0 78182 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 127070 0 127126 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 166722 0 166778 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 179200 12792 180000 12912 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 user_irq[1]
port 531 nsew signal output
rlabel metal2 s 171782 119200 171838 120000 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8251348
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_7.magic.gds
string GDS_START 282326
<< end >>

