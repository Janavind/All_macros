magic
tech sky130A
magscale 1 2
timestamp 1653073400
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 934 960 179662 117552
<< metal2 >>
rect 294 0 350 800
rect 938 0 994 800
rect 1674 0 1730 800
rect 2318 0 2374 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6550 0 6606 800
rect 7286 0 7342 800
rect 8022 0 8078 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12162 0 12218 800
rect 12898 0 12954 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 15014 0 15070 800
rect 15750 0 15806 800
rect 16394 0 16450 800
rect 17130 0 17186 800
rect 17866 0 17922 800
rect 18510 0 18566 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22006 0 22062 800
rect 22742 0 22798 800
rect 23478 0 23534 800
rect 24122 0 24178 800
rect 24858 0 24914 800
rect 25594 0 25650 800
rect 26238 0 26294 800
rect 26974 0 27030 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29090 0 29146 800
rect 29826 0 29882 800
rect 30470 0 30526 800
rect 31206 0 31262 800
rect 31942 0 31998 800
rect 32586 0 32642 800
rect 33322 0 33378 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38934 0 38990 800
rect 39670 0 39726 800
rect 40314 0 40370 800
rect 41050 0 41106 800
rect 41786 0 41842 800
rect 42430 0 42486 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44546 0 44602 800
rect 45282 0 45338 800
rect 45926 0 45982 800
rect 46662 0 46718 800
rect 47398 0 47454 800
rect 48042 0 48098 800
rect 48778 0 48834 800
rect 49514 0 49570 800
rect 50158 0 50214 800
rect 50894 0 50950 800
rect 51630 0 51686 800
rect 52274 0 52330 800
rect 53010 0 53066 800
rect 53654 0 53710 800
rect 54390 0 54446 800
rect 55126 0 55182 800
rect 55770 0 55826 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57886 0 57942 800
rect 58622 0 58678 800
rect 59358 0 59414 800
rect 60002 0 60058 800
rect 60738 0 60794 800
rect 61474 0 61530 800
rect 62118 0 62174 800
rect 62854 0 62910 800
rect 63590 0 63646 800
rect 64234 0 64290 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66350 0 66406 800
rect 67086 0 67142 800
rect 67730 0 67786 800
rect 68466 0 68522 800
rect 69202 0 69258 800
rect 69846 0 69902 800
rect 70582 0 70638 800
rect 71318 0 71374 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73434 0 73490 800
rect 74078 0 74134 800
rect 74814 0 74870 800
rect 75458 0 75514 800
rect 76194 0 76250 800
rect 76930 0 76986 800
rect 77574 0 77630 800
rect 78310 0 78366 800
rect 79046 0 79102 800
rect 79690 0 79746 800
rect 80426 0 80482 800
rect 81162 0 81218 800
rect 81806 0 81862 800
rect 82542 0 82598 800
rect 83278 0 83334 800
rect 83922 0 83978 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 86038 0 86094 800
rect 86774 0 86830 800
rect 87418 0 87474 800
rect 88154 0 88210 800
rect 88890 0 88946 800
rect 89534 0 89590 800
rect 90270 0 90326 800
rect 91006 0 91062 800
rect 91650 0 91706 800
rect 92386 0 92442 800
rect 93122 0 93178 800
rect 93766 0 93822 800
rect 94502 0 94558 800
rect 95238 0 95294 800
rect 95882 0 95938 800
rect 96618 0 96674 800
rect 97262 0 97318 800
rect 97998 0 98054 800
rect 98734 0 98790 800
rect 99378 0 99434 800
rect 100114 0 100170 800
rect 100850 0 100906 800
rect 101494 0 101550 800
rect 102230 0 102286 800
rect 102966 0 103022 800
rect 103610 0 103666 800
rect 104346 0 104402 800
rect 105082 0 105138 800
rect 105726 0 105782 800
rect 106462 0 106518 800
rect 107106 0 107162 800
rect 107842 0 107898 800
rect 108578 0 108634 800
rect 109222 0 109278 800
rect 109958 0 110014 800
rect 110694 0 110750 800
rect 111338 0 111394 800
rect 112074 0 112130 800
rect 112810 0 112866 800
rect 113454 0 113510 800
rect 114190 0 114246 800
rect 114926 0 114982 800
rect 115570 0 115626 800
rect 116306 0 116362 800
rect 116950 0 117006 800
rect 117686 0 117742 800
rect 118422 0 118478 800
rect 119066 0 119122 800
rect 119802 0 119858 800
rect 120538 0 120594 800
rect 121182 0 121238 800
rect 121918 0 121974 800
rect 122654 0 122710 800
rect 123298 0 123354 800
rect 124034 0 124090 800
rect 124770 0 124826 800
rect 125414 0 125470 800
rect 126150 0 126206 800
rect 126886 0 126942 800
rect 127530 0 127586 800
rect 128266 0 128322 800
rect 128910 0 128966 800
rect 129646 0 129702 800
rect 130382 0 130438 800
rect 131026 0 131082 800
rect 131762 0 131818 800
rect 132498 0 132554 800
rect 133142 0 133198 800
rect 133878 0 133934 800
rect 134614 0 134670 800
rect 135258 0 135314 800
rect 135994 0 136050 800
rect 136730 0 136786 800
rect 137374 0 137430 800
rect 138110 0 138166 800
rect 138754 0 138810 800
rect 139490 0 139546 800
rect 140226 0 140282 800
rect 140870 0 140926 800
rect 141606 0 141662 800
rect 142342 0 142398 800
rect 142986 0 143042 800
rect 143722 0 143778 800
rect 144458 0 144514 800
rect 145102 0 145158 800
rect 145838 0 145894 800
rect 146574 0 146630 800
rect 147218 0 147274 800
rect 147954 0 148010 800
rect 148598 0 148654 800
rect 149334 0 149390 800
rect 150070 0 150126 800
rect 150714 0 150770 800
rect 151450 0 151506 800
rect 152186 0 152242 800
rect 152830 0 152886 800
rect 153566 0 153622 800
rect 154302 0 154358 800
rect 154946 0 155002 800
rect 155682 0 155738 800
rect 156418 0 156474 800
rect 157062 0 157118 800
rect 157798 0 157854 800
rect 158534 0 158590 800
rect 159178 0 159234 800
rect 159914 0 159970 800
rect 160558 0 160614 800
rect 161294 0 161350 800
rect 162030 0 162086 800
rect 162674 0 162730 800
rect 163410 0 163466 800
rect 164146 0 164202 800
rect 164790 0 164846 800
rect 165526 0 165582 800
rect 166262 0 166318 800
rect 166906 0 166962 800
rect 167642 0 167698 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169758 0 169814 800
rect 170402 0 170458 800
rect 171138 0 171194 800
rect 171874 0 171930 800
rect 172518 0 172574 800
rect 173254 0 173310 800
rect 173990 0 174046 800
rect 174634 0 174690 800
rect 175370 0 175426 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177486 0 177542 800
rect 178222 0 178278 800
rect 178866 0 178922 800
rect 179602 0 179658 800
<< obsm2 >>
rect 940 856 179656 117552
rect 1050 734 1618 856
rect 1786 734 2262 856
rect 2430 734 2998 856
rect 3166 734 3734 856
rect 3902 734 4378 856
rect 4546 734 5114 856
rect 5282 734 5850 856
rect 6018 734 6494 856
rect 6662 734 7230 856
rect 7398 734 7966 856
rect 8134 734 8610 856
rect 8778 734 9346 856
rect 9514 734 10082 856
rect 10250 734 10726 856
rect 10894 734 11462 856
rect 11630 734 12106 856
rect 12274 734 12842 856
rect 13010 734 13578 856
rect 13746 734 14222 856
rect 14390 734 14958 856
rect 15126 734 15694 856
rect 15862 734 16338 856
rect 16506 734 17074 856
rect 17242 734 17810 856
rect 17978 734 18454 856
rect 18622 734 19190 856
rect 19358 734 19926 856
rect 20094 734 20570 856
rect 20738 734 21306 856
rect 21474 734 21950 856
rect 22118 734 22686 856
rect 22854 734 23422 856
rect 23590 734 24066 856
rect 24234 734 24802 856
rect 24970 734 25538 856
rect 25706 734 26182 856
rect 26350 734 26918 856
rect 27086 734 27654 856
rect 27822 734 28298 856
rect 28466 734 29034 856
rect 29202 734 29770 856
rect 29938 734 30414 856
rect 30582 734 31150 856
rect 31318 734 31886 856
rect 32054 734 32530 856
rect 32698 734 33266 856
rect 33434 734 33910 856
rect 34078 734 34646 856
rect 34814 734 35382 856
rect 35550 734 36026 856
rect 36194 734 36762 856
rect 36930 734 37498 856
rect 37666 734 38142 856
rect 38310 734 38878 856
rect 39046 734 39614 856
rect 39782 734 40258 856
rect 40426 734 40994 856
rect 41162 734 41730 856
rect 41898 734 42374 856
rect 42542 734 43110 856
rect 43278 734 43754 856
rect 43922 734 44490 856
rect 44658 734 45226 856
rect 45394 734 45870 856
rect 46038 734 46606 856
rect 46774 734 47342 856
rect 47510 734 47986 856
rect 48154 734 48722 856
rect 48890 734 49458 856
rect 49626 734 50102 856
rect 50270 734 50838 856
rect 51006 734 51574 856
rect 51742 734 52218 856
rect 52386 734 52954 856
rect 53122 734 53598 856
rect 53766 734 54334 856
rect 54502 734 55070 856
rect 55238 734 55714 856
rect 55882 734 56450 856
rect 56618 734 57186 856
rect 57354 734 57830 856
rect 57998 734 58566 856
rect 58734 734 59302 856
rect 59470 734 59946 856
rect 60114 734 60682 856
rect 60850 734 61418 856
rect 61586 734 62062 856
rect 62230 734 62798 856
rect 62966 734 63534 856
rect 63702 734 64178 856
rect 64346 734 64914 856
rect 65082 734 65558 856
rect 65726 734 66294 856
rect 66462 734 67030 856
rect 67198 734 67674 856
rect 67842 734 68410 856
rect 68578 734 69146 856
rect 69314 734 69790 856
rect 69958 734 70526 856
rect 70694 734 71262 856
rect 71430 734 71906 856
rect 72074 734 72642 856
rect 72810 734 73378 856
rect 73546 734 74022 856
rect 74190 734 74758 856
rect 74926 734 75402 856
rect 75570 734 76138 856
rect 76306 734 76874 856
rect 77042 734 77518 856
rect 77686 734 78254 856
rect 78422 734 78990 856
rect 79158 734 79634 856
rect 79802 734 80370 856
rect 80538 734 81106 856
rect 81274 734 81750 856
rect 81918 734 82486 856
rect 82654 734 83222 856
rect 83390 734 83866 856
rect 84034 734 84602 856
rect 84770 734 85246 856
rect 85414 734 85982 856
rect 86150 734 86718 856
rect 86886 734 87362 856
rect 87530 734 88098 856
rect 88266 734 88834 856
rect 89002 734 89478 856
rect 89646 734 90214 856
rect 90382 734 90950 856
rect 91118 734 91594 856
rect 91762 734 92330 856
rect 92498 734 93066 856
rect 93234 734 93710 856
rect 93878 734 94446 856
rect 94614 734 95182 856
rect 95350 734 95826 856
rect 95994 734 96562 856
rect 96730 734 97206 856
rect 97374 734 97942 856
rect 98110 734 98678 856
rect 98846 734 99322 856
rect 99490 734 100058 856
rect 100226 734 100794 856
rect 100962 734 101438 856
rect 101606 734 102174 856
rect 102342 734 102910 856
rect 103078 734 103554 856
rect 103722 734 104290 856
rect 104458 734 105026 856
rect 105194 734 105670 856
rect 105838 734 106406 856
rect 106574 734 107050 856
rect 107218 734 107786 856
rect 107954 734 108522 856
rect 108690 734 109166 856
rect 109334 734 109902 856
rect 110070 734 110638 856
rect 110806 734 111282 856
rect 111450 734 112018 856
rect 112186 734 112754 856
rect 112922 734 113398 856
rect 113566 734 114134 856
rect 114302 734 114870 856
rect 115038 734 115514 856
rect 115682 734 116250 856
rect 116418 734 116894 856
rect 117062 734 117630 856
rect 117798 734 118366 856
rect 118534 734 119010 856
rect 119178 734 119746 856
rect 119914 734 120482 856
rect 120650 734 121126 856
rect 121294 734 121862 856
rect 122030 734 122598 856
rect 122766 734 123242 856
rect 123410 734 123978 856
rect 124146 734 124714 856
rect 124882 734 125358 856
rect 125526 734 126094 856
rect 126262 734 126830 856
rect 126998 734 127474 856
rect 127642 734 128210 856
rect 128378 734 128854 856
rect 129022 734 129590 856
rect 129758 734 130326 856
rect 130494 734 130970 856
rect 131138 734 131706 856
rect 131874 734 132442 856
rect 132610 734 133086 856
rect 133254 734 133822 856
rect 133990 734 134558 856
rect 134726 734 135202 856
rect 135370 734 135938 856
rect 136106 734 136674 856
rect 136842 734 137318 856
rect 137486 734 138054 856
rect 138222 734 138698 856
rect 138866 734 139434 856
rect 139602 734 140170 856
rect 140338 734 140814 856
rect 140982 734 141550 856
rect 141718 734 142286 856
rect 142454 734 142930 856
rect 143098 734 143666 856
rect 143834 734 144402 856
rect 144570 734 145046 856
rect 145214 734 145782 856
rect 145950 734 146518 856
rect 146686 734 147162 856
rect 147330 734 147898 856
rect 148066 734 148542 856
rect 148710 734 149278 856
rect 149446 734 150014 856
rect 150182 734 150658 856
rect 150826 734 151394 856
rect 151562 734 152130 856
rect 152298 734 152774 856
rect 152942 734 153510 856
rect 153678 734 154246 856
rect 154414 734 154890 856
rect 155058 734 155626 856
rect 155794 734 156362 856
rect 156530 734 157006 856
rect 157174 734 157742 856
rect 157910 734 158478 856
rect 158646 734 159122 856
rect 159290 734 159858 856
rect 160026 734 160502 856
rect 160670 734 161238 856
rect 161406 734 161974 856
rect 162142 734 162618 856
rect 162786 734 163354 856
rect 163522 734 164090 856
rect 164258 734 164734 856
rect 164902 734 165470 856
rect 165638 734 166206 856
rect 166374 734 166850 856
rect 167018 734 167586 856
rect 167754 734 168322 856
rect 168490 734 168966 856
rect 169134 734 169702 856
rect 169870 734 170346 856
rect 170514 734 171082 856
rect 171250 734 171818 856
rect 171986 734 172462 856
rect 172630 734 173198 856
rect 173366 734 173934 856
rect 174102 734 174578 856
rect 174746 734 175314 856
rect 175482 734 176050 856
rect 176218 734 176694 856
rect 176862 734 177430 856
rect 177598 734 178166 856
rect 178334 734 178810 856
rect 178978 734 179546 856
<< obsm3 >>
rect 4208 1259 173488 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 60595 2048 65568 8941
rect 66048 2048 80928 8941
rect 81408 2048 85501 8941
rect 60595 1259 85501 2048
<< labels >>
rlabel metal2 s 294 0 350 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[100]
port 2 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[101]
port 3 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[102]
port 4 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[103]
port 5 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[104]
port 6 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_data_in[105]
port 7 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[106]
port 8 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[107]
port 9 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[108]
port 10 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[109]
port 11 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_data_in[10]
port 12 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[110]
port 13 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_data_in[111]
port 14 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_data_in[112]
port 15 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_data_in[113]
port 16 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_data_in[114]
port 17 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_data_in[115]
port 18 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[116]
port 19 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_data_in[117]
port 20 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[118]
port 21 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[119]
port 22 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la_data_in[11]
port 23 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[120]
port 24 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[121]
port 25 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[122]
port 26 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[123]
port 27 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_data_in[124]
port 28 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[125]
port 29 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_data_in[126]
port 30 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[127]
port 31 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[12]
port 32 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_data_in[13]
port 33 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_data_in[14]
port 34 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 la_data_in[15]
port 35 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[16]
port 36 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 la_data_in[17]
port 37 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_data_in[18]
port 38 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[19]
port 39 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 la_data_in[1]
port 40 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_data_in[20]
port 41 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_data_in[21]
port 42 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[22]
port 43 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[23]
port 44 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[24]
port 45 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[25]
port 46 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[26]
port 47 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_data_in[27]
port 48 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[28]
port 49 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[29]
port 50 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 la_data_in[2]
port 51 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in[30]
port 52 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_data_in[31]
port 53 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[32]
port 54 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[33]
port 55 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[34]
port 56 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[35]
port 57 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[36]
port 58 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_data_in[37]
port 59 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_data_in[38]
port 60 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_data_in[39]
port 61 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 la_data_in[3]
port 62 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[40]
port 63 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[41]
port 64 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[42]
port 65 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[43]
port 66 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[44]
port 67 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[45]
port 68 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[46]
port 69 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[47]
port 70 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[48]
port 71 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[49]
port 72 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 la_data_in[4]
port 73 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[50]
port 74 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[51]
port 75 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[52]
port 76 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[53]
port 77 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[54]
port 78 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[55]
port 79 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[56]
port 80 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_data_in[57]
port 81 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[58]
port 82 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[59]
port 83 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 la_data_in[5]
port 84 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[60]
port 85 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[61]
port 86 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[62]
port 87 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[63]
port 88 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[64]
port 89 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_data_in[65]
port 90 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[66]
port 91 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[67]
port 92 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[68]
port 93 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[69]
port 94 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 la_data_in[6]
port 95 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[70]
port 96 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[71]
port 97 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[72]
port 98 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[73]
port 99 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[74]
port 100 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_data_in[75]
port 101 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[76]
port 102 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[77]
port 103 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[78]
port 104 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[79]
port 105 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 la_data_in[7]
port 106 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[80]
port 107 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[81]
port 108 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[82]
port 109 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_data_in[83]
port 110 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[84]
port 111 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[85]
port 112 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[86]
port 113 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[87]
port 114 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[88]
port 115 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[89]
port 116 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_data_in[8]
port 117 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[90]
port 118 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[91]
port 119 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_data_in[92]
port 120 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[93]
port 121 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[94]
port 122 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[95]
port 123 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_data_in[96]
port 124 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[97]
port 125 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[98]
port 126 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[99]
port 127 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_data_in[9]
port 128 nsew signal input
rlabel metal2 s 938 0 994 800 6 la_data_out[0]
port 129 nsew signal output
rlabel metal2 s 141606 0 141662 800 6 la_data_out[100]
port 130 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[101]
port 131 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[102]
port 132 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[103]
port 133 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 la_data_out[104]
port 134 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[105]
port 135 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[106]
port 136 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 la_data_out[107]
port 137 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[108]
port 138 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[109]
port 139 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 la_data_out[10]
port 140 nsew signal output
rlabel metal2 s 155682 0 155738 800 6 la_data_out[110]
port 141 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[111]
port 142 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[112]
port 143 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 la_data_out[113]
port 144 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 la_data_out[114]
port 145 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[115]
port 146 nsew signal output
rlabel metal2 s 164146 0 164202 800 6 la_data_out[116]
port 147 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[117]
port 148 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[118]
port 149 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 la_data_out[119]
port 150 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 la_data_out[11]
port 151 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[120]
port 152 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[121]
port 153 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[122]
port 154 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[123]
port 155 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[124]
port 156 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[125]
port 157 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[126]
port 158 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[127]
port 159 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 la_data_out[12]
port 160 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 la_data_out[13]
port 161 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 la_data_out[14]
port 162 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_data_out[15]
port 163 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[16]
port 164 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 la_data_out[17]
port 165 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 la_data_out[18]
port 166 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[19]
port 167 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 la_data_out[1]
port 168 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[20]
port 169 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 la_data_out[21]
port 170 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[22]
port 171 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 la_data_out[23]
port 172 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[24]
port 173 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 la_data_out[25]
port 174 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[26]
port 175 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[27]
port 176 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 la_data_out[28]
port 177 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[29]
port 178 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 la_data_out[2]
port 179 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[30]
port 180 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[31]
port 181 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[32]
port 182 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[33]
port 183 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[34]
port 184 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[35]
port 185 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[36]
port 186 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 la_data_out[37]
port 187 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[38]
port 188 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[39]
port 189 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 la_data_out[3]
port 190 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[40]
port 191 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[41]
port 192 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[42]
port 193 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[43]
port 194 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[44]
port 195 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[45]
port 196 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[46]
port 197 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[47]
port 198 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 la_data_out[48]
port 199 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[49]
port 200 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 la_data_out[4]
port 201 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[50]
port 202 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[51]
port 203 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[52]
port 204 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[53]
port 205 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[54]
port 206 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 la_data_out[55]
port 207 nsew signal output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[56]
port 208 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[57]
port 209 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[58]
port 210 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[59]
port 211 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 la_data_out[5]
port 212 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[60]
port 213 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 la_data_out[61]
port 214 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[62]
port 215 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[63]
port 216 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[64]
port 217 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[65]
port 218 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[66]
port 219 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[67]
port 220 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[68]
port 221 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 la_data_out[69]
port 222 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 la_data_out[6]
port 223 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[70]
port 224 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[71]
port 225 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[72]
port 226 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[73]
port 227 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[74]
port 228 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[75]
port 229 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[76]
port 230 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[77]
port 231 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[78]
port 232 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[79]
port 233 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 la_data_out[7]
port 234 nsew signal output
rlabel metal2 s 113454 0 113510 800 6 la_data_out[80]
port 235 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[81]
port 236 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 la_data_out[82]
port 237 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 la_data_out[83]
port 238 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 la_data_out[84]
port 239 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[85]
port 240 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[86]
port 241 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[87]
port 242 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[88]
port 243 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[89]
port 244 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 la_data_out[8]
port 245 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[90]
port 246 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[91]
port 247 nsew signal output
rlabel metal2 s 130382 0 130438 800 6 la_data_out[92]
port 248 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 la_data_out[93]
port 249 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[94]
port 250 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[95]
port 251 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[96]
port 252 nsew signal output
rlabel metal2 s 137374 0 137430 800 6 la_data_out[97]
port 253 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[98]
port 254 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[99]
port 255 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 la_data_out[9]
port 256 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 257 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 258 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 258 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 258 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 258 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 258 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 258 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6593934
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_13.magic.gds
string GDS_START 267392
<< end >>

