VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.970 1421.780 1042.290 1421.840 ;
        RECT 2898.070 1421.780 2898.390 1421.840 ;
        RECT 1041.970 1421.640 2898.390 1421.780 ;
        RECT 1041.970 1421.580 1042.290 1421.640 ;
        RECT 2898.070 1421.580 2898.390 1421.640 ;
      LAYER via ;
        RECT 1042.000 1421.580 1042.260 1421.840 ;
        RECT 2898.100 1421.580 2898.360 1421.840 ;
      LAYER met2 ;
        RECT 2898.090 1426.795 2898.370 1427.165 ;
        RECT 2898.160 1421.870 2898.300 1426.795 ;
        RECT 1042.000 1421.550 1042.260 1421.870 ;
        RECT 2898.100 1421.550 2898.360 1421.870 ;
        RECT 1042.060 1048.870 1042.200 1421.550 ;
        RECT 1042.060 1048.730 1043.120 1048.870 ;
        RECT 1042.980 999.330 1043.120 1048.730 ;
        RECT 1044.650 999.330 1044.930 1000.000 ;
        RECT 1042.980 999.190 1044.930 999.330 ;
        RECT 1044.650 996.000 1044.930 999.190 ;
      LAYER via2 ;
        RECT 2898.090 1426.840 2898.370 1427.120 ;
      LAYER met3 ;
        RECT 2898.065 1427.130 2898.395 1427.145 ;
        RECT 2917.600 1427.130 2924.800 1427.580 ;
        RECT 2898.065 1426.830 2924.800 1427.130 ;
        RECT 2898.065 1426.815 2898.395 1426.830 ;
        RECT 2917.600 1426.380 2924.800 1426.830 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1006.090 998.140 1006.410 998.200 ;
        RECT 227.630 998.000 289.870 998.140 ;
        RECT 192.350 997.800 192.670 997.860 ;
        RECT 227.630 997.800 227.770 998.000 ;
        RECT 192.350 997.660 227.770 997.800 ;
        RECT 289.730 997.800 289.870 998.000 ;
        RECT 1006.090 998.000 1014.600 998.140 ;
        RECT 1006.090 997.940 1006.410 998.000 ;
        RECT 289.730 997.660 293.780 997.800 ;
        RECT 192.350 997.600 192.670 997.660 ;
        RECT 293.640 997.120 293.780 997.660 ;
        RECT 971.590 997.260 971.910 997.520 ;
        RECT 293.640 996.980 903.970 997.120 ;
        RECT 903.830 996.440 903.970 996.980 ;
        RECT 931.430 996.640 966.070 996.780 ;
        RECT 931.430 996.440 931.570 996.640 ;
        RECT 903.830 996.300 931.570 996.440 ;
        RECT 965.930 996.440 966.070 996.640 ;
        RECT 971.680 996.440 971.820 997.260 ;
        RECT 1014.460 997.120 1014.600 998.000 ;
        RECT 2228.770 997.120 2229.090 997.180 ;
        RECT 1014.460 996.980 2229.090 997.120 ;
        RECT 2228.770 996.920 2229.090 996.980 ;
        RECT 965.930 996.300 971.820 996.440 ;
      LAYER via ;
        RECT 192.380 997.600 192.640 997.860 ;
        RECT 1006.120 997.940 1006.380 998.200 ;
        RECT 971.620 997.260 971.880 997.520 ;
        RECT 2228.800 996.920 2229.060 997.180 ;
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
        RECT 2230.700 3512.170 2230.840 3517.600 ;
        RECT 2228.860 3512.030 2230.840 3512.170 ;
        RECT 1006.120 998.085 1006.380 998.230 ;
        RECT 192.380 997.570 192.640 997.890 ;
        RECT 971.610 997.715 971.890 998.085 ;
        RECT 1006.110 997.715 1006.390 998.085 ;
        RECT 192.440 617.285 192.580 997.570 ;
        RECT 971.680 997.550 971.820 997.715 ;
        RECT 971.620 997.230 971.880 997.550 ;
        RECT 2228.860 997.210 2229.000 3512.030 ;
        RECT 2228.800 996.890 2229.060 997.210 ;
        RECT 192.370 616.915 192.650 617.285 ;
      LAYER via2 ;
        RECT 971.610 997.760 971.890 998.040 ;
        RECT 1006.110 997.760 1006.390 998.040 ;
        RECT 192.370 616.960 192.650 617.240 ;
      LAYER met3 ;
        RECT 971.585 998.050 971.915 998.065 ;
        RECT 1006.085 998.050 1006.415 998.065 ;
        RECT 971.585 997.750 1006.415 998.050 ;
        RECT 971.585 997.735 971.915 997.750 ;
        RECT 1006.085 997.735 1006.415 997.750 ;
        RECT 192.345 617.250 192.675 617.265 ;
        RECT 192.345 616.950 201.170 617.250 ;
        RECT 192.345 616.935 192.675 616.950 ;
        RECT 200.870 614.840 201.170 616.950 ;
        RECT 200.000 614.240 204.000 614.840 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1089.810 395.320 1090.130 395.380 ;
        RECT 1904.470 395.320 1904.790 395.380 ;
        RECT 1089.810 395.180 1904.790 395.320 ;
        RECT 1089.810 395.120 1090.130 395.180 ;
        RECT 1904.470 395.120 1904.790 395.180 ;
      LAYER via ;
        RECT 1089.840 395.120 1090.100 395.380 ;
        RECT 1904.500 395.120 1904.760 395.380 ;
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
        RECT 1905.940 3512.170 1906.080 3517.600 ;
        RECT 1904.560 3512.030 1906.080 3512.170 ;
        RECT 1089.730 400.180 1090.010 404.000 ;
        RECT 1089.730 400.000 1090.040 400.180 ;
        RECT 1089.900 395.410 1090.040 400.000 ;
        RECT 1904.560 395.410 1904.700 3512.030 ;
        RECT 1089.840 395.090 1090.100 395.410 ;
        RECT 1904.500 395.090 1904.760 395.410 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.730 998.680 296.770 998.820 ;
        RECT 191.890 998.140 192.210 998.200 ;
        RECT 220.730 998.140 220.870 998.680 ;
        RECT 191.890 998.000 220.870 998.140 ;
        RECT 191.890 997.940 192.210 998.000 ;
        RECT 296.630 997.460 296.770 998.680 ;
        RECT 1005.720 998.340 1024.720 998.480 ;
        RECT 1005.720 997.800 1005.860 998.340 ;
        RECT 931.430 997.660 1005.860 997.800 ;
        RECT 931.430 997.460 931.570 997.660 ;
        RECT 296.630 997.320 931.570 997.460 ;
        RECT 1024.580 997.460 1024.720 998.340 ;
        RECT 1580.170 997.460 1580.490 997.520 ;
        RECT 1024.580 997.320 1580.490 997.460 ;
        RECT 1580.170 997.260 1580.490 997.320 ;
      LAYER via ;
        RECT 191.920 997.940 192.180 998.200 ;
        RECT 1580.200 997.260 1580.460 997.520 ;
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
        RECT 1581.640 3512.170 1581.780 3517.600 ;
        RECT 1580.260 3512.030 1581.780 3512.170 ;
        RECT 191.920 997.910 192.180 998.230 ;
        RECT 191.980 702.965 192.120 997.910 ;
        RECT 1580.260 997.550 1580.400 3512.030 ;
        RECT 1580.200 997.230 1580.460 997.550 ;
        RECT 191.910 702.595 192.190 702.965 ;
      LAYER via2 ;
        RECT 191.910 702.640 192.190 702.920 ;
      LAYER met3 ;
        RECT 191.885 702.930 192.215 702.945 ;
        RECT 191.885 702.630 201.170 702.930 ;
        RECT 191.885 702.615 192.215 702.630 ;
        RECT 200.870 700.520 201.170 702.630 ;
        RECT 200.000 699.920 204.000 700.520 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1068.650 1012.760 1068.970 1012.820 ;
        RECT 1255.870 1012.760 1256.190 1012.820 ;
        RECT 1068.650 1012.620 1256.190 1012.760 ;
        RECT 1068.650 1012.560 1068.970 1012.620 ;
        RECT 1255.870 1012.560 1256.190 1012.620 ;
      LAYER via ;
        RECT 1068.680 1012.560 1068.940 1012.820 ;
        RECT 1255.900 1012.560 1256.160 1012.820 ;
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
        RECT 1257.340 3512.170 1257.480 3517.600 ;
        RECT 1255.960 3512.030 1257.480 3512.170 ;
        RECT 1255.960 1012.850 1256.100 3512.030 ;
        RECT 1068.680 1012.530 1068.940 1012.850 ;
        RECT 1255.900 1012.530 1256.160 1012.850 ;
        RECT 1066.730 999.330 1067.010 1000.000 ;
        RECT 1068.740 999.330 1068.880 1012.530 ;
        RECT 1066.730 999.190 1068.880 999.330 ;
        RECT 1066.730 996.000 1067.010 999.190 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 1020.240 931.890 1020.300 ;
        RECT 1072.330 1020.240 1072.650 1020.300 ;
        RECT 931.570 1020.100 1072.650 1020.240 ;
        RECT 931.570 1020.040 931.890 1020.100 ;
        RECT 1072.330 1020.040 1072.650 1020.100 ;
      LAYER via ;
        RECT 931.600 1020.040 931.860 1020.300 ;
        RECT 1072.360 1020.040 1072.620 1020.300 ;
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
        RECT 932.580 3415.570 932.720 3517.600 ;
        RECT 931.660 3415.430 932.720 3415.570 ;
        RECT 931.660 1020.330 931.800 3415.430 ;
        RECT 931.600 1020.010 931.860 1020.330 ;
        RECT 1072.360 1020.010 1072.620 1020.330 ;
        RECT 1072.420 999.330 1072.560 1020.010 ;
        RECT 1074.090 999.330 1074.370 1000.000 ;
        RECT 1072.420 999.190 1074.370 999.330 ;
        RECT 1074.090 996.000 1074.370 999.190 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.430 998.680 1048.870 998.820 ;
        RECT 1000.430 998.140 1000.570 998.680 ;
        RECT 903.830 998.000 1000.570 998.140 ;
        RECT 607.270 997.800 607.590 997.860 ;
        RECT 903.830 997.800 903.970 998.000 ;
        RECT 607.270 997.660 903.970 997.800 ;
        RECT 1048.730 997.800 1048.870 998.680 ;
        RECT 1104.070 997.800 1104.390 997.860 ;
        RECT 1048.730 997.660 1104.390 997.800 ;
        RECT 607.270 997.600 607.590 997.660 ;
        RECT 1104.070 997.600 1104.390 997.660 ;
        RECT 1093.030 406.880 1093.350 406.940 ;
        RECT 1104.070 406.880 1104.390 406.940 ;
        RECT 1093.030 406.740 1104.390 406.880 ;
        RECT 1093.030 406.680 1093.350 406.740 ;
        RECT 1104.070 406.680 1104.390 406.740 ;
      LAYER via ;
        RECT 607.300 997.600 607.560 997.860 ;
        RECT 1104.100 997.600 1104.360 997.860 ;
        RECT 1093.060 406.680 1093.320 406.940 ;
        RECT 1104.100 406.680 1104.360 406.940 ;
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
        RECT 608.280 3512.170 608.420 3517.600 ;
        RECT 607.360 3512.030 608.420 3512.170 ;
        RECT 607.360 997.890 607.500 3512.030 ;
        RECT 607.300 997.570 607.560 997.890 ;
        RECT 1104.100 997.570 1104.360 997.890 ;
        RECT 1104.160 406.970 1104.300 997.570 ;
        RECT 1093.060 406.650 1093.320 406.970 ;
        RECT 1104.100 406.650 1104.360 406.970 ;
        RECT 1091.570 403.650 1091.850 404.000 ;
        RECT 1093.120 403.650 1093.260 406.650 ;
        RECT 1091.570 403.510 1093.260 403.650 ;
        RECT 1091.570 400.000 1091.850 403.510 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.970 1019.560 283.290 1019.620 ;
        RECT 1079.690 1019.560 1080.010 1019.620 ;
        RECT 282.970 1019.420 1080.010 1019.560 ;
        RECT 282.970 1019.360 283.290 1019.420 ;
        RECT 1079.690 1019.360 1080.010 1019.420 ;
      LAYER via ;
        RECT 283.000 1019.360 283.260 1019.620 ;
        RECT 1079.720 1019.360 1079.980 1019.620 ;
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
        RECT 283.980 3415.570 284.120 3517.600 ;
        RECT 283.060 3415.430 284.120 3415.570 ;
        RECT 283.060 1019.650 283.200 3415.430 ;
        RECT 283.000 1019.330 283.260 1019.650 ;
        RECT 1079.720 1019.330 1079.980 1019.650 ;
        RECT 1079.780 999.330 1079.920 1019.330 ;
        RECT 1081.450 999.330 1081.730 1000.000 ;
        RECT 1079.780 999.190 1081.730 999.330 ;
        RECT 1081.450 996.000 1081.730 999.190 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.410 400.180 1093.690 404.000 ;
        RECT 1093.410 400.000 1093.720 400.180 ;
        RECT 1093.580 392.885 1093.720 400.000 ;
        RECT 1093.510 392.515 1093.790 392.885 ;
      LAYER via2 ;
        RECT 1093.510 392.560 1093.790 392.840 ;
      LAYER met3 ;
        RECT -4.800 3486.850 2.400 3487.300 ;
        RECT 16.830 3486.850 17.210 3486.860 ;
        RECT -4.800 3486.550 17.210 3486.850 ;
        RECT -4.800 3486.100 2.400 3486.550 ;
        RECT 16.830 3486.540 17.210 3486.550 ;
        RECT 16.830 392.850 17.210 392.860 ;
        RECT 1093.485 392.850 1093.815 392.865 ;
        RECT 16.830 392.550 1093.815 392.850 ;
        RECT 16.830 392.540 17.210 392.550 ;
        RECT 1093.485 392.535 1093.815 392.550 ;
      LAYER via3 ;
        RECT 16.860 3486.540 17.180 3486.860 ;
        RECT 16.860 392.540 17.180 392.860 ;
      LAYER met4 ;
        RECT 16.855 3486.535 17.185 3486.865 ;
        RECT 16.870 392.865 17.170 3486.535 ;
        RECT 16.855 392.535 17.185 392.865 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.870 3225.480 14.190 3225.540 ;
        RECT 23.990 3225.480 24.310 3225.540 ;
        RECT 13.870 3225.340 24.310 3225.480 ;
        RECT 13.870 3225.280 14.190 3225.340 ;
        RECT 23.990 3225.280 24.310 3225.340 ;
        RECT 23.990 786.660 24.310 786.720 ;
        RECT 190.050 786.660 190.370 786.720 ;
        RECT 23.990 786.520 190.370 786.660 ;
        RECT 23.990 786.460 24.310 786.520 ;
        RECT 190.050 786.460 190.370 786.520 ;
      LAYER via ;
        RECT 13.900 3225.280 14.160 3225.540 ;
        RECT 24.020 3225.280 24.280 3225.540 ;
        RECT 24.020 786.460 24.280 786.720 ;
        RECT 190.080 786.460 190.340 786.720 ;
      LAYER met2 ;
        RECT 13.890 3225.395 14.170 3225.765 ;
        RECT 13.900 3225.250 14.160 3225.395 ;
        RECT 24.020 3225.250 24.280 3225.570 ;
        RECT 24.080 786.750 24.220 3225.250 ;
        RECT 24.020 786.430 24.280 786.750 ;
        RECT 190.080 786.430 190.340 786.750 ;
        RECT 190.140 785.245 190.280 786.430 ;
        RECT 190.070 784.875 190.350 785.245 ;
      LAYER via2 ;
        RECT 13.890 3225.440 14.170 3225.720 ;
        RECT 190.070 784.920 190.350 785.200 ;
      LAYER met3 ;
        RECT -4.800 3225.730 2.400 3226.180 ;
        RECT 13.865 3225.730 14.195 3225.745 ;
        RECT -4.800 3225.430 14.195 3225.730 ;
        RECT -4.800 3224.980 2.400 3225.430 ;
        RECT 13.865 3225.415 14.195 3225.430 ;
        RECT 200.000 785.600 204.000 786.200 ;
        RECT 190.045 785.210 190.375 785.225 ;
        RECT 200.870 785.210 201.170 785.600 ;
        RECT 190.045 784.910 201.170 785.210 ;
        RECT 190.045 784.895 190.375 784.910 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2965.290 2.400 2965.740 ;
        RECT 18.670 2965.290 19.050 2965.300 ;
        RECT -4.800 2964.990 19.050 2965.290 ;
        RECT -4.800 2964.540 2.400 2964.990 ;
        RECT 18.670 2964.980 19.050 2964.990 ;
        RECT 200.000 871.280 204.000 871.880 ;
        RECT 18.670 870.210 19.050 870.220 ;
        RECT 200.870 870.210 201.170 871.280 ;
        RECT 18.670 869.910 201.170 870.210 ;
        RECT 18.670 869.900 19.050 869.910 ;
      LAYER via3 ;
        RECT 18.700 2964.980 19.020 2965.300 ;
        RECT 18.700 869.900 19.020 870.220 ;
      LAYER met4 ;
        RECT 18.695 2964.975 19.025 2965.305 ;
        RECT 18.710 870.225 19.010 2964.975 ;
        RECT 18.695 869.895 19.025 870.225 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1077.390 389.540 1077.710 389.600 ;
        RECT 2903.130 389.540 2903.450 389.600 ;
        RECT 1077.390 389.400 2903.450 389.540 ;
        RECT 1077.390 389.340 1077.710 389.400 ;
        RECT 2903.130 389.340 2903.450 389.400 ;
      LAYER via ;
        RECT 1077.420 389.340 1077.680 389.600 ;
        RECT 2903.160 389.340 2903.420 389.600 ;
      LAYER met2 ;
        RECT 2903.150 1692.675 2903.430 1693.045 ;
        RECT 1077.310 400.180 1077.590 404.000 ;
        RECT 1077.310 400.000 1077.620 400.180 ;
        RECT 1077.480 389.630 1077.620 400.000 ;
        RECT 2903.220 389.630 2903.360 1692.675 ;
        RECT 1077.420 389.310 1077.680 389.630 ;
        RECT 2903.160 389.310 2903.420 389.630 ;
      LAYER via2 ;
        RECT 2903.150 1692.720 2903.430 1693.000 ;
      LAYER met3 ;
        RECT 2903.125 1693.010 2903.455 1693.025 ;
        RECT 2917.600 1693.010 2924.800 1693.460 ;
        RECT 2903.125 1692.710 2924.800 1693.010 ;
        RECT 2903.125 1692.695 2903.455 1692.710 ;
        RECT 2917.600 1692.260 2924.800 1692.710 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.250 400.180 1095.530 404.000 ;
        RECT 1095.250 400.000 1095.560 400.180 ;
        RECT 1095.420 392.205 1095.560 400.000 ;
        RECT 1095.350 391.835 1095.630 392.205 ;
      LAYER via2 ;
        RECT 1095.350 391.880 1095.630 392.160 ;
      LAYER met3 ;
        RECT -4.800 2704.170 2.400 2704.620 ;
        RECT 17.750 2704.170 18.130 2704.180 ;
        RECT -4.800 2703.870 18.130 2704.170 ;
        RECT -4.800 2703.420 2.400 2703.870 ;
        RECT 17.750 2703.860 18.130 2703.870 ;
        RECT 17.750 392.170 18.130 392.180 ;
        RECT 1095.325 392.170 1095.655 392.185 ;
        RECT 17.750 391.870 1095.655 392.170 ;
        RECT 17.750 391.860 18.130 391.870 ;
        RECT 1095.325 391.855 1095.655 391.870 ;
      LAYER via3 ;
        RECT 17.780 2703.860 18.100 2704.180 ;
        RECT 17.780 391.860 18.100 392.180 ;
      LAYER met4 ;
        RECT 17.775 2703.855 18.105 2704.185 ;
        RECT 17.790 392.185 18.090 2703.855 ;
        RECT 17.775 391.855 18.105 392.185 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2442.800 17.410 2442.860 ;
        RECT 969.290 2442.800 969.610 2442.860 ;
        RECT 17.090 2442.660 969.610 2442.800 ;
        RECT 17.090 2442.600 17.410 2442.660 ;
        RECT 969.290 2442.600 969.610 2442.660 ;
        RECT 969.290 1013.440 969.610 1013.500 ;
        RECT 1087.510 1013.440 1087.830 1013.500 ;
        RECT 969.290 1013.300 1087.830 1013.440 ;
        RECT 969.290 1013.240 969.610 1013.300 ;
        RECT 1087.510 1013.240 1087.830 1013.300 ;
      LAYER via ;
        RECT 17.120 2442.600 17.380 2442.860 ;
        RECT 969.320 2442.600 969.580 2442.860 ;
        RECT 969.320 1013.240 969.580 1013.500 ;
        RECT 1087.540 1013.240 1087.800 1013.500 ;
      LAYER met2 ;
        RECT 17.110 2443.395 17.390 2443.765 ;
        RECT 17.180 2442.890 17.320 2443.395 ;
        RECT 17.120 2442.570 17.380 2442.890 ;
        RECT 969.320 2442.570 969.580 2442.890 ;
        RECT 969.380 1013.530 969.520 2442.570 ;
        RECT 969.320 1013.210 969.580 1013.530 ;
        RECT 1087.540 1013.210 1087.800 1013.530 ;
        RECT 1087.600 999.330 1087.740 1013.210 ;
        RECT 1088.810 999.330 1089.090 1000.000 ;
        RECT 1087.600 999.190 1089.090 999.330 ;
        RECT 1088.810 996.000 1089.090 999.190 ;
      LAYER via2 ;
        RECT 17.110 2443.440 17.390 2443.720 ;
      LAYER met3 ;
        RECT -4.800 2443.730 2.400 2444.180 ;
        RECT 17.085 2443.730 17.415 2443.745 ;
        RECT -4.800 2443.430 17.415 2443.730 ;
        RECT -4.800 2442.980 2.400 2443.430 ;
        RECT 17.085 2443.415 17.415 2443.430 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2180.660 17.870 2180.720 ;
        RECT 1110.970 2180.660 1111.290 2180.720 ;
        RECT 17.550 2180.520 1111.290 2180.660 ;
        RECT 17.550 2180.460 17.870 2180.520 ;
        RECT 1110.970 2180.460 1111.290 2180.520 ;
      LAYER via ;
        RECT 17.580 2180.460 17.840 2180.720 ;
        RECT 1111.000 2180.460 1111.260 2180.720 ;
      LAYER met2 ;
        RECT 17.570 2182.955 17.850 2183.325 ;
        RECT 17.640 2180.750 17.780 2182.955 ;
        RECT 17.580 2180.430 17.840 2180.750 ;
        RECT 1111.000 2180.430 1111.260 2180.750 ;
        RECT 1111.060 702.285 1111.200 2180.430 ;
        RECT 1110.990 701.915 1111.270 702.285 ;
      LAYER via2 ;
        RECT 17.570 2183.000 17.850 2183.280 ;
        RECT 1110.990 701.960 1111.270 702.240 ;
      LAYER met3 ;
        RECT -4.800 2183.290 2.400 2183.740 ;
        RECT 17.545 2183.290 17.875 2183.305 ;
        RECT -4.800 2182.990 17.875 2183.290 ;
        RECT -4.800 2182.540 2.400 2182.990 ;
        RECT 17.545 2182.975 17.875 2182.990 ;
        RECT 1110.965 702.250 1111.295 702.265 ;
        RECT 1098.790 701.950 1111.295 702.250 ;
        RECT 1098.790 699.840 1099.090 701.950 ;
        RECT 1110.965 701.935 1111.295 701.950 ;
        RECT 1096.000 699.240 1100.000 699.840 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 959.040 17.410 959.100 ;
        RECT 190.050 959.040 190.370 959.100 ;
        RECT 17.090 958.900 190.370 959.040 ;
        RECT 17.090 958.840 17.410 958.900 ;
        RECT 190.050 958.840 190.370 958.900 ;
      LAYER via ;
        RECT 17.120 958.840 17.380 959.100 ;
        RECT 190.080 958.840 190.340 959.100 ;
      LAYER met2 ;
        RECT 17.110 1921.835 17.390 1922.205 ;
        RECT 17.180 959.130 17.320 1921.835 ;
        RECT 17.120 958.810 17.380 959.130 ;
        RECT 190.080 958.810 190.340 959.130 ;
        RECT 190.140 958.645 190.280 958.810 ;
        RECT 190.070 958.275 190.350 958.645 ;
      LAYER via2 ;
        RECT 17.110 1921.880 17.390 1922.160 ;
        RECT 190.070 958.320 190.350 958.600 ;
      LAYER met3 ;
        RECT -4.800 1922.170 2.400 1922.620 ;
        RECT 17.085 1922.170 17.415 1922.185 ;
        RECT -4.800 1921.870 17.415 1922.170 ;
        RECT -4.800 1921.420 2.400 1921.870 ;
        RECT 17.085 1921.855 17.415 1921.870 ;
        RECT 190.045 958.610 190.375 958.625 ;
        RECT 190.045 958.310 201.170 958.610 ;
        RECT 190.045 958.295 190.375 958.310 ;
        RECT 200.870 957.560 201.170 958.310 ;
        RECT 200.000 956.960 204.000 957.560 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1656.380 16.490 1656.440 ;
        RECT 1097.170 1656.380 1097.490 1656.440 ;
        RECT 16.170 1656.240 1097.490 1656.380 ;
        RECT 16.170 1656.180 16.490 1656.240 ;
        RECT 1097.170 1656.180 1097.490 1656.240 ;
      LAYER via ;
        RECT 16.200 1656.180 16.460 1656.440 ;
        RECT 1097.200 1656.180 1097.460 1656.440 ;
      LAYER met2 ;
        RECT 16.190 1661.395 16.470 1661.765 ;
        RECT 16.260 1656.470 16.400 1661.395 ;
        RECT 16.200 1656.150 16.460 1656.470 ;
        RECT 1097.200 1656.150 1097.460 1656.470 ;
        RECT 1097.260 469.270 1097.400 1656.150 ;
        RECT 1097.260 469.130 1097.860 469.270 ;
        RECT 1097.090 403.650 1097.370 404.000 ;
        RECT 1097.720 403.650 1097.860 469.130 ;
        RECT 1097.090 403.510 1097.860 403.650 ;
        RECT 1097.090 400.000 1097.370 403.510 ;
      LAYER via2 ;
        RECT 16.190 1661.440 16.470 1661.720 ;
      LAYER met3 ;
        RECT -4.800 1661.730 2.400 1662.180 ;
        RECT 16.165 1661.730 16.495 1661.745 ;
        RECT -4.800 1661.430 16.495 1661.730 ;
        RECT -4.800 1660.980 2.400 1661.430 ;
        RECT 16.165 1661.415 16.495 1661.430 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1393.900 16.490 1393.960 ;
        RECT 962.390 1393.900 962.710 1393.960 ;
        RECT 16.170 1393.760 962.710 1393.900 ;
        RECT 16.170 1393.700 16.490 1393.760 ;
        RECT 962.390 1393.700 962.710 1393.760 ;
        RECT 962.390 1013.100 962.710 1013.160 ;
        RECT 1094.870 1013.100 1095.190 1013.160 ;
        RECT 962.390 1012.960 1095.190 1013.100 ;
        RECT 962.390 1012.900 962.710 1012.960 ;
        RECT 1094.870 1012.900 1095.190 1012.960 ;
      LAYER via ;
        RECT 16.200 1393.700 16.460 1393.960 ;
        RECT 962.420 1393.700 962.680 1393.960 ;
        RECT 962.420 1012.900 962.680 1013.160 ;
        RECT 1094.900 1012.900 1095.160 1013.160 ;
      LAYER met2 ;
        RECT 16.190 1400.275 16.470 1400.645 ;
        RECT 16.260 1393.990 16.400 1400.275 ;
        RECT 16.200 1393.670 16.460 1393.990 ;
        RECT 962.420 1393.670 962.680 1393.990 ;
        RECT 962.480 1013.190 962.620 1393.670 ;
        RECT 962.420 1012.870 962.680 1013.190 ;
        RECT 1094.900 1012.870 1095.160 1013.190 ;
        RECT 1094.960 999.330 1095.100 1012.870 ;
        RECT 1096.170 999.330 1096.450 1000.000 ;
        RECT 1094.960 999.190 1096.450 999.330 ;
        RECT 1096.170 996.000 1096.450 999.190 ;
      LAYER via2 ;
        RECT 16.190 1400.320 16.470 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.165 1400.610 16.495 1400.625 ;
        RECT -4.800 1400.310 16.495 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.165 1400.295 16.495 1400.310 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1138.900 17.870 1138.960 ;
        RECT 1104.530 1138.900 1104.850 1138.960 ;
        RECT 17.550 1138.760 1104.850 1138.900 ;
        RECT 17.550 1138.700 17.870 1138.760 ;
        RECT 1104.530 1138.700 1104.850 1138.760 ;
      LAYER via ;
        RECT 17.580 1138.700 17.840 1138.960 ;
        RECT 1104.560 1138.700 1104.820 1138.960 ;
      LAYER met2 ;
        RECT 17.570 1139.835 17.850 1140.205 ;
        RECT 17.640 1138.990 17.780 1139.835 ;
        RECT 17.580 1138.670 17.840 1138.990 ;
        RECT 1104.560 1138.670 1104.820 1138.990 ;
        RECT 1104.620 821.285 1104.760 1138.670 ;
        RECT 1104.550 820.915 1104.830 821.285 ;
      LAYER via2 ;
        RECT 17.570 1139.880 17.850 1140.160 ;
        RECT 1104.550 820.960 1104.830 821.240 ;
      LAYER met3 ;
        RECT -4.800 1140.170 2.400 1140.620 ;
        RECT 17.545 1140.170 17.875 1140.185 ;
        RECT -4.800 1139.870 17.875 1140.170 ;
        RECT -4.800 1139.420 2.400 1139.870 ;
        RECT 17.545 1139.855 17.875 1139.870 ;
        RECT 1104.525 821.250 1104.855 821.265 ;
        RECT 1098.790 820.950 1104.855 821.250 ;
        RECT 1098.790 820.200 1099.090 820.950 ;
        RECT 1104.525 820.935 1104.855 820.950 ;
        RECT 1096.000 819.600 1100.000 820.200 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 394.980 17.410 395.040 ;
        RECT 1099.010 394.980 1099.330 395.040 ;
        RECT 17.090 394.840 1099.330 394.980 ;
        RECT 17.090 394.780 17.410 394.840 ;
        RECT 1099.010 394.780 1099.330 394.840 ;
      LAYER via ;
        RECT 17.120 394.780 17.380 395.040 ;
        RECT 1099.040 394.780 1099.300 395.040 ;
      LAYER met2 ;
        RECT 17.110 879.395 17.390 879.765 ;
        RECT 17.180 395.070 17.320 879.395 ;
        RECT 1098.930 400.180 1099.210 404.000 ;
        RECT 1098.930 400.000 1099.240 400.180 ;
        RECT 1099.100 395.070 1099.240 400.000 ;
        RECT 17.120 394.750 17.380 395.070 ;
        RECT 1099.040 394.750 1099.300 395.070 ;
      LAYER via2 ;
        RECT 17.110 879.440 17.390 879.720 ;
      LAYER met3 ;
        RECT -4.800 879.730 2.400 880.180 ;
        RECT 17.085 879.730 17.415 879.745 ;
        RECT -4.800 879.430 17.415 879.730 ;
        RECT -4.800 878.980 2.400 879.430 ;
        RECT 17.085 879.415 17.415 879.430 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 989.555 20.610 989.925 ;
        RECT 1111.450 989.555 1111.730 989.925 ;
        RECT 20.400 618.645 20.540 989.555 ;
        RECT 1111.520 942.325 1111.660 989.555 ;
        RECT 1111.450 941.955 1111.730 942.325 ;
        RECT 20.330 618.275 20.610 618.645 ;
      LAYER via2 ;
        RECT 20.330 989.600 20.610 989.880 ;
        RECT 1111.450 989.600 1111.730 989.880 ;
        RECT 1111.450 942.000 1111.730 942.280 ;
        RECT 20.330 618.320 20.610 618.600 ;
      LAYER met3 ;
        RECT 20.305 989.890 20.635 989.905 ;
        RECT 1111.425 989.890 1111.755 989.905 ;
        RECT 20.305 989.590 1111.755 989.890 ;
        RECT 20.305 989.575 20.635 989.590 ;
        RECT 1111.425 989.575 1111.755 989.590 ;
        RECT 1111.425 942.290 1111.755 942.305 ;
        RECT 1098.790 941.990 1111.755 942.290 ;
        RECT 1098.790 939.880 1099.090 941.990 ;
        RECT 1111.425 941.975 1111.755 941.990 ;
        RECT 1096.000 939.280 1100.000 939.880 ;
        RECT -4.800 618.610 2.400 619.060 ;
        RECT 20.305 618.610 20.635 618.625 ;
        RECT -4.800 618.310 20.635 618.610 ;
        RECT -4.800 617.860 2.400 618.310 ;
        RECT 20.305 618.295 20.635 618.310 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1081.070 393.620 1081.390 393.680 ;
        RECT 2902.670 393.620 2902.990 393.680 ;
        RECT 1081.070 393.480 2902.990 393.620 ;
        RECT 1081.070 393.420 1081.390 393.480 ;
        RECT 2902.670 393.420 2902.990 393.480 ;
      LAYER via ;
        RECT 1081.100 393.420 1081.360 393.680 ;
        RECT 2902.700 393.420 2902.960 393.680 ;
      LAYER met2 ;
        RECT 2902.690 1958.555 2902.970 1958.925 ;
        RECT 1080.990 400.180 1081.270 404.000 ;
        RECT 1080.990 400.000 1081.300 400.180 ;
        RECT 1081.160 393.710 1081.300 400.000 ;
        RECT 2902.760 393.710 2902.900 1958.555 ;
        RECT 1081.100 393.390 1081.360 393.710 ;
        RECT 2902.700 393.390 2902.960 393.710 ;
      LAYER via2 ;
        RECT 2902.690 1958.600 2902.970 1958.880 ;
      LAYER met3 ;
        RECT 2902.665 1958.890 2902.995 1958.905 ;
        RECT 2917.600 1958.890 2924.800 1959.340 ;
        RECT 2902.665 1958.590 2924.800 1958.890 ;
        RECT 2902.665 1958.575 2902.995 1958.590 ;
        RECT 2917.600 1958.140 2924.800 1958.590 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1048.870 2222.140 1049.190 2222.200 ;
        RECT 2900.830 2222.140 2901.150 2222.200 ;
        RECT 1048.870 2222.000 2901.150 2222.140 ;
        RECT 1048.870 2221.940 1049.190 2222.000 ;
        RECT 2900.830 2221.940 2901.150 2222.000 ;
      LAYER via ;
        RECT 1048.900 2221.940 1049.160 2222.200 ;
        RECT 2900.860 2221.940 2901.120 2222.200 ;
      LAYER met2 ;
        RECT 2900.850 2223.755 2901.130 2224.125 ;
        RECT 2900.920 2222.230 2901.060 2223.755 ;
        RECT 1048.900 2221.910 1049.160 2222.230 ;
        RECT 2900.860 2221.910 2901.120 2222.230 ;
        RECT 1048.960 1048.870 1049.100 2221.910 ;
        RECT 1048.960 1048.730 1050.480 1048.870 ;
        RECT 1050.340 999.330 1050.480 1048.730 ;
        RECT 1052.010 999.330 1052.290 1000.000 ;
        RECT 1050.340 999.190 1052.290 999.330 ;
        RECT 1052.010 996.000 1052.290 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2223.800 2901.130 2224.080 ;
      LAYER met3 ;
        RECT 2900.825 2224.090 2901.155 2224.105 ;
        RECT 2917.600 2224.090 2924.800 2224.540 ;
        RECT 2900.825 2223.790 2924.800 2224.090 ;
        RECT 2900.825 2223.775 2901.155 2223.790 ;
        RECT 2917.600 2223.340 2924.800 2223.790 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.770 2484.280 1056.090 2484.340 ;
        RECT 2900.830 2484.280 2901.150 2484.340 ;
        RECT 1055.770 2484.140 2901.150 2484.280 ;
        RECT 1055.770 2484.080 1056.090 2484.140 ;
        RECT 2900.830 2484.080 2901.150 2484.140 ;
      LAYER via ;
        RECT 1055.800 2484.080 1056.060 2484.340 ;
        RECT 2900.860 2484.080 2901.120 2484.340 ;
      LAYER met2 ;
        RECT 2900.850 2489.635 2901.130 2490.005 ;
        RECT 2900.920 2484.370 2901.060 2489.635 ;
        RECT 1055.800 2484.050 1056.060 2484.370 ;
        RECT 2900.860 2484.050 2901.120 2484.370 ;
        RECT 1055.860 1048.870 1056.000 2484.050 ;
        RECT 1055.860 1048.730 1057.840 1048.870 ;
        RECT 1057.700 999.330 1057.840 1048.730 ;
        RECT 1059.370 999.330 1059.650 1000.000 ;
        RECT 1057.700 999.190 1059.650 999.330 ;
        RECT 1059.370 996.000 1059.650 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2489.680 2901.130 2489.960 ;
      LAYER met3 ;
        RECT 2900.825 2489.970 2901.155 2489.985 ;
        RECT 2917.600 2489.970 2924.800 2490.420 ;
        RECT 2900.825 2489.670 2924.800 2489.970 ;
        RECT 2900.825 2489.655 2901.155 2489.670 ;
        RECT 2917.600 2489.220 2924.800 2489.670 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1082.910 393.960 1083.230 394.020 ;
        RECT 2902.210 393.960 2902.530 394.020 ;
        RECT 1082.910 393.820 2902.530 393.960 ;
        RECT 1082.910 393.760 1083.230 393.820 ;
        RECT 2902.210 393.760 2902.530 393.820 ;
      LAYER via ;
        RECT 1082.940 393.760 1083.200 394.020 ;
        RECT 2902.240 393.760 2902.500 394.020 ;
      LAYER met2 ;
        RECT 2902.230 2755.515 2902.510 2755.885 ;
        RECT 1082.830 400.180 1083.110 404.000 ;
        RECT 1082.830 400.000 1083.140 400.180 ;
        RECT 1083.000 394.050 1083.140 400.000 ;
        RECT 2902.300 394.050 2902.440 2755.515 ;
        RECT 1082.940 393.730 1083.200 394.050 ;
        RECT 2902.240 393.730 2902.500 394.050 ;
      LAYER via2 ;
        RECT 2902.230 2755.560 2902.510 2755.840 ;
      LAYER met3 ;
        RECT 2902.205 2755.850 2902.535 2755.865 ;
        RECT 2917.600 2755.850 2924.800 2756.300 ;
        RECT 2902.205 2755.550 2924.800 2755.850 ;
        RECT 2902.205 2755.535 2902.535 2755.550 ;
        RECT 2917.600 2755.100 2924.800 2755.550 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.750 392.940 1085.070 393.000 ;
        RECT 2901.750 392.940 2902.070 393.000 ;
        RECT 1084.750 392.800 2902.070 392.940 ;
        RECT 1084.750 392.740 1085.070 392.800 ;
        RECT 2901.750 392.740 2902.070 392.800 ;
      LAYER via ;
        RECT 1084.780 392.740 1085.040 393.000 ;
        RECT 2901.780 392.740 2902.040 393.000 ;
      LAYER met2 ;
        RECT 2901.770 3020.715 2902.050 3021.085 ;
        RECT 1084.670 400.180 1084.950 404.000 ;
        RECT 1084.670 400.000 1084.980 400.180 ;
        RECT 1084.840 393.030 1084.980 400.000 ;
        RECT 2901.840 393.030 2901.980 3020.715 ;
        RECT 1084.780 392.710 1085.040 393.030 ;
        RECT 2901.780 392.710 2902.040 393.030 ;
      LAYER via2 ;
        RECT 2901.770 3020.760 2902.050 3021.040 ;
      LAYER met3 ;
        RECT 2901.745 3021.050 2902.075 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2901.745 3020.750 2924.800 3021.050 ;
        RECT 2901.745 3020.735 2902.075 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1086.130 394.300 1086.450 394.360 ;
        RECT 2901.290 394.300 2901.610 394.360 ;
        RECT 1086.130 394.160 2901.610 394.300 ;
        RECT 1086.130 394.100 1086.450 394.160 ;
        RECT 2901.290 394.100 2901.610 394.160 ;
      LAYER via ;
        RECT 1086.160 394.100 1086.420 394.360 ;
        RECT 2901.320 394.100 2901.580 394.360 ;
      LAYER met2 ;
        RECT 2901.310 3286.595 2901.590 3286.965 ;
        RECT 1086.050 400.180 1086.330 404.000 ;
        RECT 1086.050 400.000 1086.360 400.180 ;
        RECT 1086.220 394.390 1086.360 400.000 ;
        RECT 2901.380 394.390 2901.520 3286.595 ;
        RECT 1086.160 394.070 1086.420 394.390 ;
        RECT 2901.320 394.070 2901.580 394.390 ;
      LAYER via2 ;
        RECT 2901.310 3286.640 2901.590 3286.920 ;
      LAYER met3 ;
        RECT 2901.285 3286.930 2901.615 3286.945 ;
        RECT 2917.600 3286.930 2924.800 3287.380 ;
        RECT 2901.285 3286.630 2924.800 3286.930 ;
        RECT 2901.285 3286.615 2901.615 3286.630 ;
        RECT 2917.600 3286.180 2924.800 3286.630 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
        RECT 2879.300 3512.170 2879.440 3517.600 ;
        RECT 2877.460 3512.030 2879.440 3512.170 ;
        RECT 2877.460 996.725 2877.600 3512.030 ;
        RECT 192.830 996.355 193.110 996.725 ;
        RECT 2877.390 996.355 2877.670 996.725 ;
        RECT 192.900 530.925 193.040 996.355 ;
        RECT 192.830 530.555 193.110 530.925 ;
      LAYER via2 ;
        RECT 192.830 996.400 193.110 996.680 ;
        RECT 2877.390 996.400 2877.670 996.680 ;
        RECT 192.830 530.600 193.110 530.880 ;
      LAYER met3 ;
        RECT 192.805 996.690 193.135 996.705 ;
        RECT 2877.365 996.690 2877.695 996.705 ;
        RECT 192.805 996.390 2877.695 996.690 ;
        RECT 192.805 996.375 193.135 996.390 ;
        RECT 2877.365 996.375 2877.695 996.390 ;
        RECT 192.805 530.890 193.135 530.905 ;
        RECT 192.805 530.590 201.170 530.890 ;
        RECT 192.805 530.575 193.135 530.590 ;
        RECT 200.870 529.160 201.170 530.590 ;
        RECT 200.000 528.560 204.000 529.160 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1087.970 394.640 1088.290 394.700 ;
        RECT 2553.070 394.640 2553.390 394.700 ;
        RECT 1087.970 394.500 2553.390 394.640 ;
        RECT 1087.970 394.440 1088.290 394.500 ;
        RECT 2553.070 394.440 2553.390 394.500 ;
      LAYER via ;
        RECT 1088.000 394.440 1088.260 394.700 ;
        RECT 2553.100 394.440 2553.360 394.700 ;
      LAYER met2 ;
        RECT 2553.160 3517.910 2554.220 3518.050 ;
        RECT 1087.890 400.180 1088.170 404.000 ;
        RECT 1087.890 400.000 1088.200 400.180 ;
        RECT 1088.060 394.730 1088.200 400.000 ;
        RECT 2553.160 394.730 2553.300 3517.910 ;
        RECT 2554.080 3517.370 2554.220 3517.910 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
        RECT 2555.000 3517.370 2555.140 3517.600 ;
        RECT 2554.080 3517.230 2555.140 3517.370 ;
        RECT 1088.000 394.410 1088.260 394.730 ;
        RECT 2553.100 394.410 2553.360 394.730 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.170 372.880 200.490 372.940 ;
        RECT 201.550 372.880 201.870 372.940 ;
        RECT 200.170 372.740 201.870 372.880 ;
        RECT 200.170 372.680 200.490 372.740 ;
        RECT 201.550 372.680 201.870 372.740 ;
      LAYER via ;
        RECT 200.200 372.680 200.460 372.940 ;
        RECT 201.580 372.680 201.840 372.940 ;
      LAYER met2 ;
        RECT 203.770 996.610 204.050 1000.000 ;
        RECT 201.640 996.470 204.050 996.610 ;
        RECT 201.640 420.970 201.780 996.470 ;
        RECT 203.770 996.000 204.050 996.470 ;
        RECT 200.260 420.830 201.780 420.970 ;
        RECT 200.260 372.970 200.400 420.830 ;
        RECT 200.200 372.650 200.460 372.970 ;
        RECT 201.580 372.650 201.840 372.970 ;
        RECT 201.640 106.605 201.780 372.650 ;
        RECT 201.570 106.235 201.850 106.605 ;
        RECT 2901.310 106.235 2901.590 106.605 ;
        RECT 2901.380 33.165 2901.520 106.235 ;
        RECT 2901.310 32.795 2901.590 33.165 ;
      LAYER via2 ;
        RECT 201.570 106.280 201.850 106.560 ;
        RECT 2901.310 106.280 2901.590 106.560 ;
        RECT 2901.310 32.840 2901.590 33.120 ;
      LAYER met3 ;
        RECT 201.545 106.570 201.875 106.585 ;
        RECT 2901.285 106.570 2901.615 106.585 ;
        RECT 201.545 106.270 2901.615 106.570 ;
        RECT 201.545 106.255 201.875 106.270 ;
        RECT 2901.285 106.255 2901.615 106.270 ;
        RECT 2901.285 33.130 2901.615 33.145 ;
        RECT 2917.600 33.130 2924.800 33.580 ;
        RECT 2901.285 32.830 2924.800 33.130 ;
        RECT 2901.285 32.815 2901.615 32.830 ;
        RECT 2917.600 32.380 2924.800 32.830 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 2284.020 421.290 2284.080 ;
        RECT 2898.070 2284.020 2898.390 2284.080 ;
        RECT 420.970 2283.880 2898.390 2284.020 ;
        RECT 420.970 2283.820 421.290 2283.880 ;
        RECT 2898.070 2283.820 2898.390 2283.880 ;
      LAYER via ;
        RECT 421.000 2283.820 421.260 2284.080 ;
        RECT 2898.100 2283.820 2898.360 2284.080 ;
      LAYER met2 ;
        RECT 2898.090 2290.395 2898.370 2290.765 ;
        RECT 2898.160 2284.110 2898.300 2290.395 ;
        RECT 421.000 2283.790 421.260 2284.110 ;
        RECT 2898.100 2283.790 2898.360 2284.110 ;
        RECT 421.060 1048.870 421.200 2283.790 ;
        RECT 421.060 1048.730 423.040 1048.870 ;
        RECT 422.900 999.330 423.040 1048.730 ;
        RECT 425.030 999.330 425.310 1000.000 ;
        RECT 422.900 999.190 425.310 999.330 ;
        RECT 425.030 996.000 425.310 999.190 ;
      LAYER via2 ;
        RECT 2898.090 2290.440 2898.370 2290.720 ;
      LAYER met3 ;
        RECT 2898.065 2290.730 2898.395 2290.745 ;
        RECT 2917.600 2290.730 2924.800 2291.180 ;
        RECT 2898.065 2290.430 2924.800 2290.730 ;
        RECT 2898.065 2290.415 2898.395 2290.430 ;
        RECT 2917.600 2289.980 2924.800 2290.430 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 2553.300 441.990 2553.360 ;
        RECT 2900.830 2553.300 2901.150 2553.360 ;
        RECT 441.670 2553.160 2901.150 2553.300 ;
        RECT 441.670 2553.100 441.990 2553.160 ;
        RECT 2900.830 2553.100 2901.150 2553.160 ;
      LAYER via ;
        RECT 441.700 2553.100 441.960 2553.360 ;
        RECT 2900.860 2553.100 2901.120 2553.360 ;
      LAYER met2 ;
        RECT 2900.850 2556.275 2901.130 2556.645 ;
        RECT 2900.920 2553.390 2901.060 2556.275 ;
        RECT 441.700 2553.070 441.960 2553.390 ;
        RECT 2900.860 2553.070 2901.120 2553.390 ;
        RECT 441.760 1048.870 441.900 2553.070 ;
        RECT 441.760 1048.730 445.120 1048.870 ;
        RECT 444.980 999.330 445.120 1048.730 ;
        RECT 447.110 999.330 447.390 1000.000 ;
        RECT 444.980 999.190 447.390 999.330 ;
        RECT 447.110 996.000 447.390 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2556.320 2901.130 2556.600 ;
      LAYER met3 ;
        RECT 2900.825 2556.610 2901.155 2556.625 ;
        RECT 2917.600 2556.610 2924.800 2557.060 ;
        RECT 2900.825 2556.310 2924.800 2556.610 ;
        RECT 2900.825 2556.295 2901.155 2556.310 ;
        RECT 2917.600 2555.860 2924.800 2556.310 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 2815.440 469.590 2815.500 ;
        RECT 2899.450 2815.440 2899.770 2815.500 ;
        RECT 469.270 2815.300 2899.770 2815.440 ;
        RECT 469.270 2815.240 469.590 2815.300 ;
        RECT 2899.450 2815.240 2899.770 2815.300 ;
      LAYER via ;
        RECT 469.300 2815.240 469.560 2815.500 ;
        RECT 2899.480 2815.240 2899.740 2815.500 ;
      LAYER met2 ;
        RECT 2899.470 2821.475 2899.750 2821.845 ;
        RECT 2899.540 2815.530 2899.680 2821.475 ;
        RECT 469.300 2815.210 469.560 2815.530 ;
        RECT 2899.480 2815.210 2899.740 2815.530 ;
        RECT 469.360 1048.870 469.500 2815.210 ;
        RECT 469.360 1048.730 469.960 1048.870 ;
        RECT 469.190 999.330 469.470 1000.000 ;
        RECT 469.820 999.330 469.960 1048.730 ;
        RECT 469.190 999.190 469.960 999.330 ;
        RECT 469.190 996.000 469.470 999.190 ;
      LAYER via2 ;
        RECT 2899.470 2821.520 2899.750 2821.800 ;
      LAYER met3 ;
        RECT 2899.445 2821.810 2899.775 2821.825 ;
        RECT 2917.600 2821.810 2924.800 2822.260 ;
        RECT 2899.445 2821.510 2924.800 2821.810 ;
        RECT 2899.445 2821.495 2899.775 2821.510 ;
        RECT 2917.600 2821.060 2924.800 2821.510 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 3084.380 490.290 3084.440 ;
        RECT 2900.830 3084.380 2901.150 3084.440 ;
        RECT 489.970 3084.240 2901.150 3084.380 ;
        RECT 489.970 3084.180 490.290 3084.240 ;
        RECT 2900.830 3084.180 2901.150 3084.240 ;
      LAYER via ;
        RECT 490.000 3084.180 490.260 3084.440 ;
        RECT 2900.860 3084.180 2901.120 3084.440 ;
      LAYER met2 ;
        RECT 2900.850 3087.355 2901.130 3087.725 ;
        RECT 2900.920 3084.470 2901.060 3087.355 ;
        RECT 490.000 3084.150 490.260 3084.470 ;
        RECT 2900.860 3084.150 2901.120 3084.470 ;
        RECT 490.060 999.330 490.200 3084.150 ;
        RECT 491.270 999.330 491.550 1000.000 ;
        RECT 490.060 999.190 491.550 999.330 ;
        RECT 491.270 996.000 491.550 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3087.400 2901.130 3087.680 ;
      LAYER met3 ;
        RECT 2900.825 3087.690 2901.155 3087.705 ;
        RECT 2917.600 3087.690 2924.800 3088.140 ;
        RECT 2900.825 3087.390 2924.800 3087.690 ;
        RECT 2900.825 3087.375 2901.155 3087.390 ;
        RECT 2917.600 3086.940 2924.800 3087.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 3353.660 510.990 3353.720 ;
        RECT 2900.830 3353.660 2901.150 3353.720 ;
        RECT 510.670 3353.520 2901.150 3353.660 ;
        RECT 510.670 3353.460 510.990 3353.520 ;
        RECT 2900.830 3353.460 2901.150 3353.520 ;
      LAYER via ;
        RECT 510.700 3353.460 510.960 3353.720 ;
        RECT 2900.860 3353.460 2901.120 3353.720 ;
      LAYER met2 ;
        RECT 510.700 3353.430 510.960 3353.750 ;
        RECT 2900.860 3353.605 2901.120 3353.750 ;
        RECT 510.760 1048.870 510.900 3353.430 ;
        RECT 2900.850 3353.235 2901.130 3353.605 ;
        RECT 510.760 1048.730 511.360 1048.870 ;
        RECT 511.220 999.330 511.360 1048.730 ;
        RECT 513.350 999.330 513.630 1000.000 ;
        RECT 511.220 999.190 513.630 999.330 ;
        RECT 513.350 996.000 513.630 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3353.280 2901.130 3353.560 ;
      LAYER met3 ;
        RECT 2900.825 3353.570 2901.155 3353.585 ;
        RECT 2917.600 3353.570 2924.800 3354.020 ;
        RECT 2900.825 3353.270 2924.800 3353.570 ;
        RECT 2900.825 3353.255 2901.155 3353.270 ;
        RECT 2917.600 3352.820 2924.800 3353.270 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 533.210 1017.860 533.530 1017.920 ;
        RECT 2794.570 1017.860 2794.890 1017.920 ;
        RECT 533.210 1017.720 2794.890 1017.860 ;
        RECT 533.210 1017.660 533.530 1017.720 ;
        RECT 2794.570 1017.660 2794.890 1017.720 ;
      LAYER via ;
        RECT 533.240 1017.660 533.500 1017.920 ;
        RECT 2794.600 1017.660 2794.860 1017.920 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3512.170 2798.480 3517.600 ;
        RECT 2794.660 3512.030 2798.480 3512.170 ;
        RECT 2794.660 1017.950 2794.800 3512.030 ;
        RECT 533.240 1017.630 533.500 1017.950 ;
        RECT 2794.600 1017.630 2794.860 1017.950 ;
        RECT 533.300 999.330 533.440 1017.630 ;
        RECT 535.430 999.330 535.710 1000.000 ;
        RECT 533.300 999.190 535.710 999.330 ;
        RECT 535.430 996.000 535.710 999.190 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.290 1018.200 555.610 1018.260 ;
        RECT 2470.270 1018.200 2470.590 1018.260 ;
        RECT 555.290 1018.060 2470.590 1018.200 ;
        RECT 555.290 1018.000 555.610 1018.060 ;
        RECT 2470.270 1018.000 2470.590 1018.060 ;
      LAYER via ;
        RECT 555.320 1018.000 555.580 1018.260 ;
        RECT 2470.300 1018.000 2470.560 1018.260 ;
      LAYER met2 ;
        RECT 2470.360 3517.910 2473.260 3518.050 ;
        RECT 2470.360 1018.290 2470.500 3517.910 ;
        RECT 2473.120 3517.370 2473.260 3517.910 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2473.120 3517.230 2474.180 3517.370 ;
        RECT 555.320 1017.970 555.580 1018.290 ;
        RECT 2470.300 1017.970 2470.560 1018.290 ;
        RECT 555.380 999.330 555.520 1017.970 ;
        RECT 557.510 999.330 557.790 1000.000 ;
        RECT 555.380 999.190 557.790 999.330 ;
        RECT 557.510 996.000 557.790 999.190 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.670 1018.540 579.990 1018.600 ;
        RECT 2145.970 1018.540 2146.290 1018.600 ;
        RECT 579.670 1018.400 2146.290 1018.540 ;
        RECT 579.670 1018.340 579.990 1018.400 ;
        RECT 2145.970 1018.340 2146.290 1018.400 ;
      LAYER via ;
        RECT 579.700 1018.340 579.960 1018.600 ;
        RECT 2146.000 1018.340 2146.260 1018.600 ;
      LAYER met2 ;
        RECT 2146.060 3517.910 2148.500 3518.050 ;
        RECT 2146.060 1018.630 2146.200 3517.910 ;
        RECT 2148.360 3517.370 2148.500 3517.910 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2148.360 3517.230 2149.420 3517.370 ;
        RECT 579.700 1018.310 579.960 1018.630 ;
        RECT 2146.000 1018.310 2146.260 1018.630 ;
        RECT 579.760 999.330 579.900 1018.310 ;
        RECT 580.050 999.330 580.330 1000.000 ;
        RECT 579.760 999.190 580.330 999.330 ;
        RECT 580.050 996.000 580.330 999.190 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 1018.880 600.690 1018.940 ;
        RECT 1821.670 1018.880 1821.990 1018.940 ;
        RECT 600.370 1018.740 1821.990 1018.880 ;
        RECT 600.370 1018.680 600.690 1018.740 ;
        RECT 1821.670 1018.680 1821.990 1018.740 ;
      LAYER via ;
        RECT 600.400 1018.680 600.660 1018.940 ;
        RECT 1821.700 1018.680 1821.960 1018.940 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3512.170 1825.120 3517.600 ;
        RECT 1821.760 3512.030 1825.120 3512.170 ;
        RECT 1821.760 1018.970 1821.900 3512.030 ;
        RECT 600.400 1018.650 600.660 1018.970 ;
        RECT 1821.700 1018.650 1821.960 1018.970 ;
        RECT 600.460 999.330 600.600 1018.650 ;
        RECT 602.130 999.330 602.410 1000.000 ;
        RECT 600.460 999.190 602.410 999.330 ;
        RECT 602.130 996.000 602.410 999.190 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 1019.220 622.770 1019.280 ;
        RECT 1497.370 1019.220 1497.690 1019.280 ;
        RECT 622.450 1019.080 1497.690 1019.220 ;
        RECT 622.450 1019.020 622.770 1019.080 ;
        RECT 1497.370 1019.020 1497.690 1019.080 ;
      LAYER via ;
        RECT 622.480 1019.020 622.740 1019.280 ;
        RECT 1497.400 1019.020 1497.660 1019.280 ;
      LAYER met2 ;
        RECT 1497.460 3517.910 1499.900 3518.050 ;
        RECT 1497.460 1019.310 1497.600 3517.910 ;
        RECT 1499.760 3517.370 1499.900 3517.910 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3517.370 1500.820 3517.600 ;
        RECT 1499.760 3517.230 1500.820 3517.370 ;
        RECT 622.480 1018.990 622.740 1019.310 ;
        RECT 1497.400 1018.990 1497.660 1019.310 ;
        RECT 622.540 999.330 622.680 1018.990 ;
        RECT 624.210 999.330 624.490 1000.000 ;
        RECT 622.540 999.190 624.490 999.330 ;
        RECT 624.210 996.000 624.490 999.190 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 1007.915 228.070 1008.285 ;
        RECT 2900.850 1007.915 2901.130 1008.285 ;
        RECT 225.850 999.330 226.130 1000.000 ;
        RECT 227.860 999.330 228.000 1007.915 ;
        RECT 225.850 999.190 228.000 999.330 ;
        RECT 225.850 996.000 226.130 999.190 ;
        RECT 2900.920 231.725 2901.060 1007.915 ;
        RECT 2900.850 231.355 2901.130 231.725 ;
      LAYER via2 ;
        RECT 227.790 1007.960 228.070 1008.240 ;
        RECT 2900.850 1007.960 2901.130 1008.240 ;
        RECT 2900.850 231.400 2901.130 231.680 ;
      LAYER met3 ;
        RECT 227.765 1008.250 228.095 1008.265 ;
        RECT 2900.825 1008.250 2901.155 1008.265 ;
        RECT 227.765 1007.950 2901.155 1008.250 ;
        RECT 227.765 1007.935 228.095 1007.950 ;
        RECT 2900.825 1007.935 2901.155 1007.950 ;
        RECT 2900.825 231.690 2901.155 231.705 ;
        RECT 2917.600 231.690 2924.800 232.140 ;
        RECT 2900.825 231.390 2924.800 231.690 ;
        RECT 2900.825 231.375 2901.155 231.390 ;
        RECT 2917.600 230.940 2924.800 231.390 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 644.530 1019.900 644.850 1019.960 ;
        RECT 1173.070 1019.900 1173.390 1019.960 ;
        RECT 644.530 1019.760 1173.390 1019.900 ;
        RECT 644.530 1019.700 644.850 1019.760 ;
        RECT 1173.070 1019.700 1173.390 1019.760 ;
      LAYER via ;
        RECT 644.560 1019.700 644.820 1019.960 ;
        RECT 1173.100 1019.700 1173.360 1019.960 ;
      LAYER met2 ;
        RECT 1173.160 3517.910 1175.140 3518.050 ;
        RECT 1173.160 1019.990 1173.300 3517.910 ;
        RECT 1175.000 3517.370 1175.140 3517.910 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3517.370 1176.060 3517.600 ;
        RECT 1175.000 3517.230 1176.060 3517.370 ;
        RECT 644.560 1019.670 644.820 1019.990 ;
        RECT 1173.100 1019.670 1173.360 1019.990 ;
        RECT 644.620 999.330 644.760 1019.670 ;
        RECT 646.290 999.330 646.570 1000.000 ;
        RECT 644.620 999.190 646.570 999.330 ;
        RECT 646.290 996.000 646.570 999.190 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 666.610 1020.240 666.930 1020.300 ;
        RECT 848.770 1020.240 849.090 1020.300 ;
        RECT 666.610 1020.100 849.090 1020.240 ;
        RECT 666.610 1020.040 666.930 1020.100 ;
        RECT 848.770 1020.040 849.090 1020.100 ;
      LAYER via ;
        RECT 666.640 1020.040 666.900 1020.300 ;
        RECT 848.800 1020.040 849.060 1020.300 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3512.170 851.760 3517.600 ;
        RECT 848.860 3512.030 851.760 3512.170 ;
        RECT 848.860 1020.330 849.000 3512.030 ;
        RECT 666.640 1020.010 666.900 1020.330 ;
        RECT 848.800 1020.010 849.060 1020.330 ;
        RECT 666.700 999.330 666.840 1020.010 ;
        RECT 668.370 999.330 668.650 1000.000 ;
        RECT 666.700 999.190 668.650 999.330 ;
        RECT 668.370 996.000 668.650 999.190 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3500.200 527.550 3500.260 ;
        RECT 690.070 3500.200 690.390 3500.260 ;
        RECT 527.230 3500.060 690.390 3500.200 ;
        RECT 527.230 3500.000 527.550 3500.060 ;
        RECT 690.070 3500.000 690.390 3500.060 ;
      LAYER via ;
        RECT 527.260 3500.000 527.520 3500.260 ;
        RECT 690.100 3500.000 690.360 3500.260 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3500.290 527.460 3517.600 ;
        RECT 527.260 3499.970 527.520 3500.290 ;
        RECT 690.100 3499.970 690.360 3500.290 ;
        RECT 690.160 999.330 690.300 3499.970 ;
        RECT 690.450 999.330 690.730 1000.000 ;
        RECT 690.160 999.190 690.730 999.330 ;
        RECT 690.450 996.000 690.730 999.190 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3504.620 202.790 3504.680 ;
        RECT 710.770 3504.620 711.090 3504.680 ;
        RECT 202.470 3504.480 711.090 3504.620 ;
        RECT 202.470 3504.420 202.790 3504.480 ;
        RECT 710.770 3504.420 711.090 3504.480 ;
      LAYER via ;
        RECT 202.500 3504.420 202.760 3504.680 ;
        RECT 710.800 3504.420 711.060 3504.680 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3504.710 202.700 3517.600 ;
        RECT 202.500 3504.390 202.760 3504.710 ;
        RECT 710.800 3504.390 711.060 3504.710 ;
        RECT 710.860 999.330 711.000 3504.390 ;
        RECT 712.530 999.330 712.810 1000.000 ;
        RECT 710.860 999.190 712.810 999.330 ;
        RECT 712.530 996.000 712.810 999.190 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3416.220 17.410 3416.280 ;
        RECT 731.470 3416.220 731.790 3416.280 ;
        RECT 17.090 3416.080 731.790 3416.220 ;
        RECT 17.090 3416.020 17.410 3416.080 ;
        RECT 731.470 3416.020 731.790 3416.080 ;
      LAYER via ;
        RECT 17.120 3416.020 17.380 3416.280 ;
        RECT 731.500 3416.020 731.760 3416.280 ;
      LAYER met2 ;
        RECT 17.110 3421.235 17.390 3421.605 ;
        RECT 17.180 3416.310 17.320 3421.235 ;
        RECT 17.120 3415.990 17.380 3416.310 ;
        RECT 731.500 3415.990 731.760 3416.310 ;
        RECT 731.560 1048.870 731.700 3415.990 ;
        RECT 731.560 1048.730 733.080 1048.870 ;
        RECT 732.940 999.330 733.080 1048.730 ;
        RECT 734.610 999.330 734.890 1000.000 ;
        RECT 732.940 999.190 734.890 999.330 ;
        RECT 734.610 996.000 734.890 999.190 ;
      LAYER via2 ;
        RECT 17.110 3421.280 17.390 3421.560 ;
      LAYER met3 ;
        RECT -4.800 3421.570 2.400 3422.020 ;
        RECT 17.085 3421.570 17.415 3421.585 ;
        RECT -4.800 3421.270 17.415 3421.570 ;
        RECT -4.800 3420.820 2.400 3421.270 ;
        RECT 17.085 3421.255 17.415 3421.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3160.540 17.410 3160.600 ;
        RECT 752.170 3160.540 752.490 3160.600 ;
        RECT 17.090 3160.400 752.490 3160.540 ;
        RECT 17.090 3160.340 17.410 3160.400 ;
        RECT 752.170 3160.340 752.490 3160.400 ;
      LAYER via ;
        RECT 17.120 3160.340 17.380 3160.600 ;
        RECT 752.200 3160.340 752.460 3160.600 ;
      LAYER met2 ;
        RECT 17.120 3160.485 17.380 3160.630 ;
        RECT 17.110 3160.115 17.390 3160.485 ;
        RECT 752.200 3160.310 752.460 3160.630 ;
        RECT 752.260 1048.870 752.400 3160.310 ;
        RECT 752.260 1048.730 755.160 1048.870 ;
        RECT 755.020 999.330 755.160 1048.730 ;
        RECT 757.150 999.330 757.430 1000.000 ;
        RECT 755.020 999.190 757.430 999.330 ;
        RECT 757.150 996.000 757.430 999.190 ;
      LAYER via2 ;
        RECT 17.110 3160.160 17.390 3160.440 ;
      LAYER met3 ;
        RECT -4.800 3160.450 2.400 3160.900 ;
        RECT 17.085 3160.450 17.415 3160.465 ;
        RECT -4.800 3160.150 17.415 3160.450 ;
        RECT -4.800 3159.700 2.400 3160.150 ;
        RECT 17.085 3160.135 17.415 3160.150 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2898.400 16.950 2898.460 ;
        RECT 772.870 2898.400 773.190 2898.460 ;
        RECT 16.630 2898.260 773.190 2898.400 ;
        RECT 16.630 2898.200 16.950 2898.260 ;
        RECT 772.870 2898.200 773.190 2898.260 ;
      LAYER via ;
        RECT 16.660 2898.200 16.920 2898.460 ;
        RECT 772.900 2898.200 773.160 2898.460 ;
      LAYER met2 ;
        RECT 16.650 2899.675 16.930 2900.045 ;
        RECT 16.720 2898.490 16.860 2899.675 ;
        RECT 16.660 2898.170 16.920 2898.490 ;
        RECT 772.900 2898.170 773.160 2898.490 ;
        RECT 772.960 1048.870 773.100 2898.170 ;
        RECT 772.960 1048.730 777.240 1048.870 ;
        RECT 777.100 999.330 777.240 1048.730 ;
        RECT 779.230 999.330 779.510 1000.000 ;
        RECT 777.100 999.190 779.510 999.330 ;
        RECT 779.230 996.000 779.510 999.190 ;
      LAYER via2 ;
        RECT 16.650 2899.720 16.930 2900.000 ;
      LAYER met3 ;
        RECT -4.800 2900.010 2.400 2900.460 ;
        RECT 16.625 2900.010 16.955 2900.025 ;
        RECT -4.800 2899.710 16.955 2900.010 ;
        RECT -4.800 2899.260 2.400 2899.710 ;
        RECT 16.625 2899.695 16.955 2899.710 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2635.920 17.410 2635.980 ;
        RECT 800.470 2635.920 800.790 2635.980 ;
        RECT 17.090 2635.780 800.790 2635.920 ;
        RECT 17.090 2635.720 17.410 2635.780 ;
        RECT 800.470 2635.720 800.790 2635.780 ;
      LAYER via ;
        RECT 17.120 2635.720 17.380 2635.980 ;
        RECT 800.500 2635.720 800.760 2635.980 ;
      LAYER met2 ;
        RECT 17.110 2639.235 17.390 2639.605 ;
        RECT 17.180 2636.010 17.320 2639.235 ;
        RECT 17.120 2635.690 17.380 2636.010 ;
        RECT 800.500 2635.690 800.760 2636.010 ;
        RECT 800.560 999.330 800.700 2635.690 ;
        RECT 801.310 999.330 801.590 1000.000 ;
        RECT 800.560 999.190 801.590 999.330 ;
        RECT 801.310 996.000 801.590 999.190 ;
      LAYER via2 ;
        RECT 17.110 2639.280 17.390 2639.560 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 17.085 2639.570 17.415 2639.585 ;
        RECT -4.800 2639.270 17.415 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 17.085 2639.255 17.415 2639.270 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2373.780 17.410 2373.840 ;
        RECT 821.170 2373.780 821.490 2373.840 ;
        RECT 17.090 2373.640 821.490 2373.780 ;
        RECT 17.090 2373.580 17.410 2373.640 ;
        RECT 821.170 2373.580 821.490 2373.640 ;
      LAYER via ;
        RECT 17.120 2373.580 17.380 2373.840 ;
        RECT 821.200 2373.580 821.460 2373.840 ;
      LAYER met2 ;
        RECT 17.110 2378.115 17.390 2378.485 ;
        RECT 17.180 2373.870 17.320 2378.115 ;
        RECT 17.120 2373.550 17.380 2373.870 ;
        RECT 821.200 2373.550 821.460 2373.870 ;
        RECT 821.260 999.330 821.400 2373.550 ;
        RECT 823.390 999.330 823.670 1000.000 ;
        RECT 821.260 999.190 823.670 999.330 ;
        RECT 823.390 996.000 823.670 999.190 ;
      LAYER via2 ;
        RECT 17.110 2378.160 17.390 2378.440 ;
      LAYER met3 ;
        RECT -4.800 2378.450 2.400 2378.900 ;
        RECT 17.085 2378.450 17.415 2378.465 ;
        RECT -4.800 2378.150 17.415 2378.450 ;
        RECT -4.800 2377.700 2.400 2378.150 ;
        RECT 17.085 2378.135 17.415 2378.150 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2111.640 17.410 2111.700 ;
        RECT 841.870 2111.640 842.190 2111.700 ;
        RECT 17.090 2111.500 842.190 2111.640 ;
        RECT 17.090 2111.440 17.410 2111.500 ;
        RECT 841.870 2111.440 842.190 2111.500 ;
      LAYER via ;
        RECT 17.120 2111.440 17.380 2111.700 ;
        RECT 841.900 2111.440 842.160 2111.700 ;
      LAYER met2 ;
        RECT 17.110 2117.675 17.390 2118.045 ;
        RECT 17.180 2111.730 17.320 2117.675 ;
        RECT 17.120 2111.410 17.380 2111.730 ;
        RECT 841.900 2111.410 842.160 2111.730 ;
        RECT 841.960 1048.870 842.100 2111.410 ;
        RECT 841.960 1048.730 843.480 1048.870 ;
        RECT 843.340 999.330 843.480 1048.730 ;
        RECT 845.470 999.330 845.750 1000.000 ;
        RECT 843.340 999.190 845.750 999.330 ;
        RECT 845.470 996.000 845.750 999.190 ;
      LAYER via2 ;
        RECT 17.110 2117.720 17.390 2118.000 ;
      LAYER met3 ;
        RECT -4.800 2118.010 2.400 2118.460 ;
        RECT 17.085 2118.010 17.415 2118.025 ;
        RECT -4.800 2117.710 17.415 2118.010 ;
        RECT -4.800 2117.260 2.400 2117.710 ;
        RECT 17.085 2117.695 17.415 2117.710 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 249.850 1000.860 250.170 1000.920 ;
        RECT 2900.370 1000.860 2900.690 1000.920 ;
        RECT 249.850 1000.720 2900.690 1000.860 ;
        RECT 249.850 1000.660 250.170 1000.720 ;
        RECT 2900.370 1000.660 2900.690 1000.720 ;
      LAYER via ;
        RECT 249.880 1000.660 250.140 1000.920 ;
        RECT 2900.400 1000.660 2900.660 1000.920 ;
      LAYER met2 ;
        RECT 249.880 1000.630 250.140 1000.950 ;
        RECT 2900.400 1000.630 2900.660 1000.950 ;
        RECT 247.930 999.330 248.210 1000.000 ;
        RECT 249.940 999.330 250.080 1000.630 ;
        RECT 247.930 999.190 250.080 999.330 ;
        RECT 247.930 996.000 248.210 999.190 ;
        RECT 2900.460 430.965 2900.600 1000.630 ;
        RECT 2900.390 430.595 2900.670 430.965 ;
      LAYER via2 ;
        RECT 2900.390 430.640 2900.670 430.920 ;
      LAYER met3 ;
        RECT 2900.365 430.930 2900.695 430.945 ;
        RECT 2917.600 430.930 2924.800 431.380 ;
        RECT 2900.365 430.630 2924.800 430.930 ;
        RECT 2900.365 430.615 2900.695 430.630 ;
        RECT 2917.600 430.180 2924.800 430.630 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1856.300 17.870 1856.360 ;
        RECT 862.570 1856.300 862.890 1856.360 ;
        RECT 17.550 1856.160 862.890 1856.300 ;
        RECT 17.550 1856.100 17.870 1856.160 ;
        RECT 862.570 1856.100 862.890 1856.160 ;
      LAYER via ;
        RECT 17.580 1856.100 17.840 1856.360 ;
        RECT 862.600 1856.100 862.860 1856.360 ;
      LAYER met2 ;
        RECT 17.570 1856.555 17.850 1856.925 ;
        RECT 17.640 1856.390 17.780 1856.555 ;
        RECT 17.580 1856.070 17.840 1856.390 ;
        RECT 862.600 1856.070 862.860 1856.390 ;
        RECT 862.660 1048.870 862.800 1856.070 ;
        RECT 862.660 1048.730 865.560 1048.870 ;
        RECT 865.420 999.330 865.560 1048.730 ;
        RECT 867.550 999.330 867.830 1000.000 ;
        RECT 865.420 999.190 867.830 999.330 ;
        RECT 867.550 996.000 867.830 999.190 ;
      LAYER via2 ;
        RECT 17.570 1856.600 17.850 1856.880 ;
      LAYER met3 ;
        RECT -4.800 1856.890 2.400 1857.340 ;
        RECT 17.545 1856.890 17.875 1856.905 ;
        RECT -4.800 1856.590 17.875 1856.890 ;
        RECT -4.800 1856.140 2.400 1856.590 ;
        RECT 17.545 1856.575 17.875 1856.590 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1594.160 16.950 1594.220 ;
        RECT 883.270 1594.160 883.590 1594.220 ;
        RECT 16.630 1594.020 883.590 1594.160 ;
        RECT 16.630 1593.960 16.950 1594.020 ;
        RECT 883.270 1593.960 883.590 1594.020 ;
      LAYER via ;
        RECT 16.660 1593.960 16.920 1594.220 ;
        RECT 883.300 1593.960 883.560 1594.220 ;
      LAYER met2 ;
        RECT 16.650 1596.115 16.930 1596.485 ;
        RECT 16.720 1594.250 16.860 1596.115 ;
        RECT 16.660 1593.930 16.920 1594.250 ;
        RECT 883.300 1593.930 883.560 1594.250 ;
        RECT 883.360 1048.870 883.500 1593.930 ;
        RECT 883.360 1048.730 887.640 1048.870 ;
        RECT 887.500 999.330 887.640 1048.730 ;
        RECT 889.630 999.330 889.910 1000.000 ;
        RECT 887.500 999.190 889.910 999.330 ;
        RECT 889.630 996.000 889.910 999.190 ;
      LAYER via2 ;
        RECT 16.650 1596.160 16.930 1596.440 ;
      LAYER met3 ;
        RECT -4.800 1596.450 2.400 1596.900 ;
        RECT 16.625 1596.450 16.955 1596.465 ;
        RECT -4.800 1596.150 16.955 1596.450 ;
        RECT -4.800 1595.700 2.400 1596.150 ;
        RECT 16.625 1596.135 16.955 1596.150 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1332.020 15.570 1332.080 ;
        RECT 910.870 1332.020 911.190 1332.080 ;
        RECT 15.250 1331.880 911.190 1332.020 ;
        RECT 15.250 1331.820 15.570 1331.880 ;
        RECT 910.870 1331.820 911.190 1331.880 ;
      LAYER via ;
        RECT 15.280 1331.820 15.540 1332.080 ;
        RECT 910.900 1331.820 911.160 1332.080 ;
      LAYER met2 ;
        RECT 15.270 1335.675 15.550 1336.045 ;
        RECT 15.340 1332.110 15.480 1335.675 ;
        RECT 15.280 1331.790 15.540 1332.110 ;
        RECT 910.900 1331.790 911.160 1332.110 ;
        RECT 910.960 999.330 911.100 1331.790 ;
        RECT 911.710 999.330 911.990 1000.000 ;
        RECT 910.960 999.190 911.990 999.330 ;
        RECT 911.710 996.000 911.990 999.190 ;
      LAYER via2 ;
        RECT 15.270 1335.720 15.550 1336.000 ;
      LAYER met3 ;
        RECT -4.800 1336.010 2.400 1336.460 ;
        RECT 15.245 1336.010 15.575 1336.025 ;
        RECT -4.800 1335.710 15.575 1336.010 ;
        RECT -4.800 1335.260 2.400 1335.710 ;
        RECT 15.245 1335.695 15.575 1335.710 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1069.880 16.030 1069.940 ;
        RECT 932.030 1069.880 932.350 1069.940 ;
        RECT 15.710 1069.740 932.350 1069.880 ;
        RECT 15.710 1069.680 16.030 1069.740 ;
        RECT 932.030 1069.680 932.350 1069.740 ;
      LAYER via ;
        RECT 15.740 1069.680 16.000 1069.940 ;
        RECT 932.060 1069.680 932.320 1069.940 ;
      LAYER met2 ;
        RECT 15.730 1074.555 16.010 1074.925 ;
        RECT 15.800 1069.970 15.940 1074.555 ;
        RECT 15.740 1069.650 16.000 1069.970 ;
        RECT 932.060 1069.650 932.320 1069.970 ;
        RECT 932.120 1048.870 932.260 1069.650 ;
        RECT 932.120 1048.730 932.720 1048.870 ;
        RECT 932.580 999.330 932.720 1048.730 ;
        RECT 934.250 999.330 934.530 1000.000 ;
        RECT 932.580 999.190 934.530 999.330 ;
        RECT 934.250 996.000 934.530 999.190 ;
      LAYER via2 ;
        RECT 15.730 1074.600 16.010 1074.880 ;
      LAYER met3 ;
        RECT -4.800 1074.890 2.400 1075.340 ;
        RECT 15.705 1074.890 16.035 1074.905 ;
        RECT -4.800 1074.590 16.035 1074.890 ;
        RECT -4.800 1074.140 2.400 1074.590 ;
        RECT 15.705 1074.575 16.035 1074.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1009.700 16.030 1009.760 ;
        RECT 955.030 1009.700 955.350 1009.760 ;
        RECT 15.710 1009.560 955.350 1009.700 ;
        RECT 15.710 1009.500 16.030 1009.560 ;
        RECT 955.030 1009.500 955.350 1009.560 ;
      LAYER via ;
        RECT 15.740 1009.500 16.000 1009.760 ;
        RECT 955.060 1009.500 955.320 1009.760 ;
      LAYER met2 ;
        RECT 15.740 1009.470 16.000 1009.790 ;
        RECT 955.060 1009.470 955.320 1009.790 ;
        RECT 15.800 814.485 15.940 1009.470 ;
        RECT 955.120 999.330 955.260 1009.470 ;
        RECT 956.330 999.330 956.610 1000.000 ;
        RECT 955.120 999.190 956.610 999.330 ;
        RECT 956.330 996.000 956.610 999.190 ;
        RECT 15.730 814.115 16.010 814.485 ;
      LAYER via2 ;
        RECT 15.730 814.160 16.010 814.440 ;
      LAYER met3 ;
        RECT -4.800 814.450 2.400 814.900 ;
        RECT 15.705 814.450 16.035 814.465 ;
        RECT -4.800 814.150 16.035 814.450 ;
        RECT -4.800 813.700 2.400 814.150 ;
        RECT 15.705 814.135 16.035 814.150 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.950 997.800 243.270 997.860 ;
        RECT 242.950 997.660 262.270 997.800 ;
        RECT 242.950 997.600 243.270 997.660 ;
        RECT 220.870 997.460 221.190 997.520 ;
        RECT 242.030 997.460 242.350 997.520 ;
        RECT 220.870 997.320 242.350 997.460 ;
        RECT 262.130 997.460 262.270 997.660 ;
        RECT 977.110 997.460 977.430 997.520 ;
        RECT 262.130 997.320 289.870 997.460 ;
        RECT 220.870 997.260 221.190 997.320 ;
        RECT 242.030 997.260 242.350 997.320 ;
        RECT 289.730 996.440 289.870 997.320 ;
        RECT 973.520 997.320 977.430 997.460 ;
        RECT 289.730 996.300 296.770 996.440 ;
        RECT 19.850 994.740 20.170 994.800 ;
        RECT 200.630 994.740 200.950 994.800 ;
        RECT 19.850 994.600 200.950 994.740 ;
        RECT 296.630 994.740 296.770 996.300 ;
        RECT 973.520 994.740 973.660 997.320 ;
        RECT 977.110 997.260 977.430 997.320 ;
        RECT 296.630 994.600 973.660 994.740 ;
        RECT 19.850 994.540 20.170 994.600 ;
        RECT 200.630 994.540 200.950 994.600 ;
      LAYER via ;
        RECT 242.980 997.600 243.240 997.860 ;
        RECT 220.900 997.260 221.160 997.520 ;
        RECT 242.060 997.260 242.320 997.520 ;
        RECT 19.880 994.540 20.140 994.800 ;
        RECT 200.660 994.540 200.920 994.800 ;
        RECT 977.140 997.260 977.400 997.520 ;
      LAYER met2 ;
        RECT 200.650 997.715 200.930 998.085 ;
        RECT 220.890 997.715 221.170 998.085 ;
        RECT 200.720 994.830 200.860 997.715 ;
        RECT 220.960 997.550 221.100 997.715 ;
        RECT 242.980 997.570 243.240 997.890 ;
        RECT 220.900 997.230 221.160 997.550 ;
        RECT 242.060 997.290 242.320 997.550 ;
        RECT 243.040 997.290 243.180 997.570 ;
        RECT 242.060 997.230 243.180 997.290 ;
        RECT 977.140 997.290 977.400 997.550 ;
        RECT 978.410 997.290 978.690 1000.000 ;
        RECT 977.140 997.230 978.690 997.290 ;
        RECT 242.120 997.150 243.180 997.230 ;
        RECT 977.200 997.150 978.690 997.230 ;
        RECT 978.410 996.000 978.690 997.150 ;
        RECT 19.880 994.510 20.140 994.830 ;
        RECT 200.660 994.510 200.920 994.830 ;
        RECT 19.940 553.365 20.080 994.510 ;
        RECT 19.870 552.995 20.150 553.365 ;
      LAYER via2 ;
        RECT 200.650 997.760 200.930 998.040 ;
        RECT 220.890 997.760 221.170 998.040 ;
        RECT 19.870 553.040 20.150 553.320 ;
      LAYER met3 ;
        RECT 200.625 998.050 200.955 998.065 ;
        RECT 220.865 998.050 221.195 998.065 ;
        RECT 200.625 997.750 221.195 998.050 ;
        RECT 200.625 997.735 200.955 997.750 ;
        RECT 220.865 997.735 221.195 997.750 ;
        RECT -4.800 553.330 2.400 553.780 ;
        RECT 19.845 553.330 20.175 553.345 ;
        RECT -4.800 553.030 20.175 553.330 ;
        RECT -4.800 552.580 2.400 553.030 ;
        RECT 19.845 553.015 20.175 553.030 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 1008.000 18.790 1008.060 ;
        RECT 1001.030 1008.000 1001.350 1008.060 ;
        RECT 18.470 1007.860 1001.350 1008.000 ;
        RECT 18.470 1007.800 18.790 1007.860 ;
        RECT 1001.030 1007.800 1001.350 1007.860 ;
      LAYER via ;
        RECT 18.500 1007.800 18.760 1008.060 ;
        RECT 1001.060 1007.800 1001.320 1008.060 ;
      LAYER met2 ;
        RECT 18.500 1007.770 18.760 1008.090 ;
        RECT 1001.060 1007.770 1001.320 1008.090 ;
        RECT 18.560 358.205 18.700 1007.770 ;
        RECT 1000.490 999.330 1000.770 1000.000 ;
        RECT 1001.120 999.330 1001.260 1007.770 ;
        RECT 1000.490 999.190 1001.260 999.330 ;
        RECT 1000.490 996.000 1000.770 999.190 ;
        RECT 18.490 357.835 18.770 358.205 ;
      LAYER via2 ;
        RECT 18.490 357.880 18.770 358.160 ;
      LAYER met3 ;
        RECT -4.800 358.170 2.400 358.620 ;
        RECT 18.465 358.170 18.795 358.185 ;
        RECT -4.800 357.870 18.795 358.170 ;
        RECT -4.800 357.420 2.400 357.870 ;
        RECT 18.465 357.855 18.795 357.870 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1007.660 17.870 1007.720 ;
        RECT 1021.270 1007.660 1021.590 1007.720 ;
        RECT 17.550 1007.520 1021.590 1007.660 ;
        RECT 17.550 1007.460 17.870 1007.520 ;
        RECT 1021.270 1007.460 1021.590 1007.520 ;
      LAYER via ;
        RECT 17.580 1007.460 17.840 1007.720 ;
        RECT 1021.300 1007.460 1021.560 1007.720 ;
      LAYER met2 ;
        RECT 17.580 1007.430 17.840 1007.750 ;
        RECT 1021.300 1007.430 1021.560 1007.750 ;
        RECT 17.640 162.365 17.780 1007.430 ;
        RECT 1021.360 999.330 1021.500 1007.430 ;
        RECT 1022.570 999.330 1022.850 1000.000 ;
        RECT 1021.360 999.190 1022.850 999.330 ;
        RECT 1022.570 996.000 1022.850 999.190 ;
        RECT 17.570 161.995 17.850 162.365 ;
      LAYER via2 ;
        RECT 17.570 162.040 17.850 162.320 ;
      LAYER met3 ;
        RECT -4.800 162.330 2.400 162.780 ;
        RECT 17.545 162.330 17.875 162.345 ;
        RECT -4.800 162.030 17.875 162.330 ;
        RECT -4.800 161.580 2.400 162.030 ;
        RECT 17.545 162.015 17.875 162.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 271.930 1011.060 272.250 1011.120 ;
        RECT 1093.490 1011.060 1093.810 1011.120 ;
        RECT 271.930 1010.920 1093.810 1011.060 ;
        RECT 271.930 1010.860 272.250 1010.920 ;
        RECT 1093.490 1010.860 1093.810 1010.920 ;
        RECT 1094.870 634.680 1095.190 634.740 ;
        RECT 2899.450 634.680 2899.770 634.740 ;
        RECT 1094.870 634.540 2899.770 634.680 ;
        RECT 1094.870 634.480 1095.190 634.540 ;
        RECT 2899.450 634.480 2899.770 634.540 ;
      LAYER via ;
        RECT 271.960 1010.860 272.220 1011.120 ;
        RECT 1093.520 1010.860 1093.780 1011.120 ;
        RECT 1094.900 634.480 1095.160 634.740 ;
        RECT 2899.480 634.480 2899.740 634.740 ;
      LAYER met2 ;
        RECT 271.960 1010.830 272.220 1011.150 ;
        RECT 1093.520 1010.830 1093.780 1011.150 ;
        RECT 270.010 999.330 270.290 1000.000 ;
        RECT 272.020 999.330 272.160 1010.830 ;
        RECT 270.010 999.190 272.160 999.330 ;
        RECT 270.010 996.000 270.290 999.190 ;
        RECT 1093.580 759.070 1093.720 1010.830 ;
        RECT 1093.580 758.930 1095.100 759.070 ;
        RECT 1094.960 634.770 1095.100 758.930 ;
        RECT 1094.900 634.450 1095.160 634.770 ;
        RECT 2899.480 634.450 2899.740 634.770 ;
        RECT 2899.540 630.205 2899.680 634.450 ;
        RECT 2899.470 629.835 2899.750 630.205 ;
      LAYER via2 ;
        RECT 2899.470 629.880 2899.750 630.160 ;
      LAYER met3 ;
        RECT 2899.445 630.170 2899.775 630.185 ;
        RECT 2917.600 630.170 2924.800 630.620 ;
        RECT 2899.445 629.870 2924.800 630.170 ;
        RECT 2899.445 629.855 2899.775 629.870 ;
        RECT 2917.600 629.420 2924.800 629.870 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.010 1011.740 294.330 1011.800 ;
        RECT 1102.230 1011.740 1102.550 1011.800 ;
        RECT 294.010 1011.600 1102.550 1011.740 ;
        RECT 294.010 1011.540 294.330 1011.600 ;
        RECT 1102.230 1011.540 1102.550 1011.600 ;
        RECT 1102.230 834.940 1102.550 835.000 ;
        RECT 2899.450 834.940 2899.770 835.000 ;
        RECT 1102.230 834.800 2899.770 834.940 ;
        RECT 1102.230 834.740 1102.550 834.800 ;
        RECT 2899.450 834.740 2899.770 834.800 ;
      LAYER via ;
        RECT 294.040 1011.540 294.300 1011.800 ;
        RECT 1102.260 1011.540 1102.520 1011.800 ;
        RECT 1102.260 834.740 1102.520 835.000 ;
        RECT 2899.480 834.740 2899.740 835.000 ;
      LAYER met2 ;
        RECT 294.040 1011.510 294.300 1011.830 ;
        RECT 1102.260 1011.510 1102.520 1011.830 ;
        RECT 292.090 999.330 292.370 1000.000 ;
        RECT 294.100 999.330 294.240 1011.510 ;
        RECT 292.090 999.190 294.240 999.330 ;
        RECT 292.090 996.000 292.370 999.190 ;
        RECT 1102.320 835.030 1102.460 1011.510 ;
        RECT 1102.260 834.710 1102.520 835.030 ;
        RECT 2899.480 834.710 2899.740 835.030 ;
        RECT 2899.540 829.445 2899.680 834.710 ;
        RECT 2899.470 829.075 2899.750 829.445 ;
      LAYER via2 ;
        RECT 2899.470 829.120 2899.750 829.400 ;
      LAYER met3 ;
        RECT 2899.445 829.410 2899.775 829.425 ;
        RECT 2917.600 829.410 2924.800 829.860 ;
        RECT 2899.445 829.110 2924.800 829.410 ;
        RECT 2899.445 829.095 2899.775 829.110 ;
        RECT 2917.600 828.660 2924.800 829.110 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 315.630 1028.400 315.950 1028.460 ;
        RECT 2900.830 1028.400 2901.150 1028.460 ;
        RECT 315.630 1028.260 2901.150 1028.400 ;
        RECT 315.630 1028.200 315.950 1028.260 ;
        RECT 2900.830 1028.200 2901.150 1028.260 ;
      LAYER via ;
        RECT 315.660 1028.200 315.920 1028.460 ;
        RECT 2900.860 1028.200 2901.120 1028.460 ;
      LAYER met2 ;
        RECT 315.660 1028.170 315.920 1028.490 ;
        RECT 2900.850 1028.315 2901.130 1028.685 ;
        RECT 2900.860 1028.170 2901.120 1028.315 ;
        RECT 314.170 999.330 314.450 1000.000 ;
        RECT 315.720 999.330 315.860 1028.170 ;
        RECT 314.170 999.190 315.860 999.330 ;
        RECT 314.170 996.000 314.450 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1028.360 2901.130 1028.640 ;
      LAYER met3 ;
        RECT 2900.825 1028.650 2901.155 1028.665 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2900.825 1028.350 2924.800 1028.650 ;
        RECT 2900.825 1028.335 2901.155 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 1221.520 331.590 1221.580 ;
        RECT 2900.830 1221.520 2901.150 1221.580 ;
        RECT 331.270 1221.380 2901.150 1221.520 ;
        RECT 331.270 1221.320 331.590 1221.380 ;
        RECT 2900.830 1221.320 2901.150 1221.380 ;
      LAYER via ;
        RECT 331.300 1221.320 331.560 1221.580 ;
        RECT 2900.860 1221.320 2901.120 1221.580 ;
      LAYER met2 ;
        RECT 2900.850 1227.555 2901.130 1227.925 ;
        RECT 2900.920 1221.610 2901.060 1227.555 ;
        RECT 331.300 1221.290 331.560 1221.610 ;
        RECT 2900.860 1221.290 2901.120 1221.610 ;
        RECT 331.360 1048.870 331.500 1221.290 ;
        RECT 331.360 1048.730 334.720 1048.870 ;
        RECT 334.580 999.330 334.720 1048.730 ;
        RECT 336.250 999.330 336.530 1000.000 ;
        RECT 334.580 999.190 336.530 999.330 ;
        RECT 336.250 996.000 336.530 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1227.600 2901.130 1227.880 ;
      LAYER met3 ;
        RECT 2900.825 1227.890 2901.155 1227.905 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2900.825 1227.590 2924.800 1227.890 ;
        RECT 2900.825 1227.575 2901.155 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.970 1490.800 352.290 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 351.970 1490.660 2901.150 1490.800 ;
        RECT 351.970 1490.600 352.290 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 352.000 1490.600 352.260 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1493.435 2901.130 1493.805 ;
        RECT 2900.920 1490.890 2901.060 1493.435 ;
        RECT 352.000 1490.570 352.260 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 352.060 1048.870 352.200 1490.570 ;
        RECT 352.060 1048.730 356.800 1048.870 ;
        RECT 356.660 999.330 356.800 1048.730 ;
        RECT 358.330 999.330 358.610 1000.000 ;
        RECT 356.660 999.190 358.610 999.330 ;
        RECT 358.330 996.000 358.610 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1493.480 2901.130 1493.760 ;
      LAYER met3 ;
        RECT 2900.825 1493.770 2901.155 1493.785 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2900.825 1493.470 2924.800 1493.770 ;
        RECT 2900.825 1493.455 2901.155 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.570 1759.740 379.890 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 379.570 1759.600 2901.150 1759.740 ;
        RECT 379.570 1759.540 379.890 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
      LAYER via ;
        RECT 379.600 1759.540 379.860 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
      LAYER met2 ;
        RECT 379.600 1759.510 379.860 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 379.660 999.330 379.800 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 380.410 999.330 380.690 1000.000 ;
        RECT 379.660 999.190 380.690 999.330 ;
        RECT 380.410 996.000 380.690 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 2021.880 400.590 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 400.270 2021.740 2901.150 2021.880 ;
        RECT 400.270 2021.680 400.590 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 400.300 2021.680 400.560 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2024.515 2901.130 2024.885 ;
        RECT 2900.920 2021.970 2901.060 2024.515 ;
        RECT 400.300 2021.650 400.560 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 400.360 1048.870 400.500 2021.650 ;
        RECT 400.360 1048.730 400.960 1048.870 ;
        RECT 400.820 999.330 400.960 1048.730 ;
        RECT 402.950 999.330 403.230 1000.000 ;
        RECT 400.820 999.190 403.230 999.330 ;
        RECT 402.950 996.000 403.230 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2024.560 2901.130 2024.840 ;
      LAYER met3 ;
        RECT 2900.825 2024.850 2901.155 2024.865 ;
        RECT 2917.600 2024.850 2924.800 2025.300 ;
        RECT 2900.825 2024.550 2924.800 2024.850 ;
        RECT 2900.825 2024.535 2901.155 2024.550 ;
        RECT 2917.600 2024.100 2924.800 2024.550 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 1007.235 213.350 1007.605 ;
        RECT 2904.070 1007.235 2904.350 1007.605 ;
        RECT 211.130 999.330 211.410 1000.000 ;
        RECT 213.140 999.330 213.280 1007.235 ;
        RECT 211.130 999.190 213.280 999.330 ;
        RECT 211.130 996.000 211.410 999.190 ;
        RECT 2904.140 165.765 2904.280 1007.235 ;
        RECT 2904.070 165.395 2904.350 165.765 ;
      LAYER via2 ;
        RECT 213.070 1007.280 213.350 1007.560 ;
        RECT 2904.070 1007.280 2904.350 1007.560 ;
        RECT 2904.070 165.440 2904.350 165.720 ;
      LAYER met3 ;
        RECT 213.045 1007.570 213.375 1007.585 ;
        RECT 2904.045 1007.570 2904.375 1007.585 ;
        RECT 213.045 1007.270 2904.375 1007.570 ;
        RECT 213.045 1007.255 213.375 1007.270 ;
        RECT 2904.045 1007.255 2904.375 1007.270 ;
        RECT 2904.045 165.730 2904.375 165.745 ;
        RECT 2917.600 165.730 2924.800 166.180 ;
        RECT 2904.045 165.430 2924.800 165.730 ;
        RECT 2904.045 165.415 2904.375 165.430 ;
        RECT 2917.600 164.980 2924.800 165.430 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 2422.060 428.190 2422.120 ;
        RECT 2900.830 2422.060 2901.150 2422.120 ;
        RECT 427.870 2421.920 2901.150 2422.060 ;
        RECT 427.870 2421.860 428.190 2421.920 ;
        RECT 2900.830 2421.860 2901.150 2421.920 ;
      LAYER via ;
        RECT 427.900 2421.860 428.160 2422.120 ;
        RECT 2900.860 2421.860 2901.120 2422.120 ;
      LAYER met2 ;
        RECT 2900.850 2422.995 2901.130 2423.365 ;
        RECT 2900.920 2422.150 2901.060 2422.995 ;
        RECT 427.900 2421.830 428.160 2422.150 ;
        RECT 2900.860 2421.830 2901.120 2422.150 ;
        RECT 427.960 1048.870 428.100 2421.830 ;
        RECT 427.960 1048.730 430.400 1048.870 ;
        RECT 430.260 999.330 430.400 1048.730 ;
        RECT 432.390 999.330 432.670 1000.000 ;
        RECT 430.260 999.190 432.670 999.330 ;
        RECT 432.390 996.000 432.670 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2423.040 2901.130 2423.320 ;
      LAYER met3 ;
        RECT 2900.825 2423.330 2901.155 2423.345 ;
        RECT 2917.600 2423.330 2924.800 2423.780 ;
        RECT 2900.825 2423.030 2924.800 2423.330 ;
        RECT 2900.825 2423.015 2901.155 2423.030 ;
        RECT 2917.600 2422.580 2924.800 2423.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 2684.200 448.890 2684.260 ;
        RECT 2900.830 2684.200 2901.150 2684.260 ;
        RECT 448.570 2684.060 2901.150 2684.200 ;
        RECT 448.570 2684.000 448.890 2684.060 ;
        RECT 2900.830 2684.000 2901.150 2684.060 ;
      LAYER via ;
        RECT 448.600 2684.000 448.860 2684.260 ;
        RECT 2900.860 2684.000 2901.120 2684.260 ;
      LAYER met2 ;
        RECT 2900.850 2688.875 2901.130 2689.245 ;
        RECT 2900.920 2684.290 2901.060 2688.875 ;
        RECT 448.600 2683.970 448.860 2684.290 ;
        RECT 2900.860 2683.970 2901.120 2684.290 ;
        RECT 448.660 1048.870 448.800 2683.970 ;
        RECT 448.660 1048.730 452.480 1048.870 ;
        RECT 452.340 999.330 452.480 1048.730 ;
        RECT 454.470 999.330 454.750 1000.000 ;
        RECT 452.340 999.190 454.750 999.330 ;
        RECT 454.470 996.000 454.750 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2688.920 2901.130 2689.200 ;
      LAYER met3 ;
        RECT 2900.825 2689.210 2901.155 2689.225 ;
        RECT 2917.600 2689.210 2924.800 2689.660 ;
        RECT 2900.825 2688.910 2924.800 2689.210 ;
        RECT 2900.825 2688.895 2901.155 2688.910 ;
        RECT 2917.600 2688.460 2924.800 2688.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 2953.480 476.490 2953.540 ;
        RECT 2898.070 2953.480 2898.390 2953.540 ;
        RECT 476.170 2953.340 2898.390 2953.480 ;
        RECT 476.170 2953.280 476.490 2953.340 ;
        RECT 2898.070 2953.280 2898.390 2953.340 ;
      LAYER via ;
        RECT 476.200 2953.280 476.460 2953.540 ;
        RECT 2898.100 2953.280 2898.360 2953.540 ;
      LAYER met2 ;
        RECT 2898.090 2954.755 2898.370 2955.125 ;
        RECT 2898.160 2953.570 2898.300 2954.755 ;
        RECT 476.200 2953.250 476.460 2953.570 ;
        RECT 2898.100 2953.250 2898.360 2953.570 ;
        RECT 476.260 999.330 476.400 2953.250 ;
        RECT 476.550 999.330 476.830 1000.000 ;
        RECT 476.260 999.190 476.830 999.330 ;
        RECT 476.550 996.000 476.830 999.190 ;
      LAYER via2 ;
        RECT 2898.090 2954.800 2898.370 2955.080 ;
      LAYER met3 ;
        RECT 2898.065 2955.090 2898.395 2955.105 ;
        RECT 2917.600 2955.090 2924.800 2955.540 ;
        RECT 2898.065 2954.790 2924.800 2955.090 ;
        RECT 2898.065 2954.775 2898.395 2954.790 ;
        RECT 2917.600 2954.340 2924.800 2954.790 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 3215.620 497.190 3215.680 ;
        RECT 2900.830 3215.620 2901.150 3215.680 ;
        RECT 496.870 3215.480 2901.150 3215.620 ;
        RECT 496.870 3215.420 497.190 3215.480 ;
        RECT 2900.830 3215.420 2901.150 3215.480 ;
      LAYER via ;
        RECT 496.900 3215.420 497.160 3215.680 ;
        RECT 2900.860 3215.420 2901.120 3215.680 ;
      LAYER met2 ;
        RECT 2900.850 3219.955 2901.130 3220.325 ;
        RECT 2900.920 3215.710 2901.060 3219.955 ;
        RECT 496.900 3215.390 497.160 3215.710 ;
        RECT 2900.860 3215.390 2901.120 3215.710 ;
        RECT 496.960 999.330 497.100 3215.390 ;
        RECT 498.630 999.330 498.910 1000.000 ;
        RECT 496.960 999.190 498.910 999.330 ;
        RECT 498.630 996.000 498.910 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3220.000 2901.130 3220.280 ;
      LAYER met3 ;
        RECT 2900.825 3220.290 2901.155 3220.305 ;
        RECT 2917.600 3220.290 2924.800 3220.740 ;
        RECT 2900.825 3219.990 2924.800 3220.290 ;
        RECT 2900.825 3219.975 2901.155 3219.990 ;
        RECT 2917.600 3219.540 2924.800 3219.990 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 3484.900 517.890 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 517.570 3484.760 2901.150 3484.900 ;
        RECT 517.570 3484.700 517.890 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 517.600 3484.700 517.860 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3485.835 2901.130 3486.205 ;
        RECT 2900.920 3484.990 2901.060 3485.835 ;
        RECT 517.600 3484.670 517.860 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 517.660 1048.870 517.800 3484.670 ;
        RECT 517.660 1048.730 518.720 1048.870 ;
        RECT 518.580 999.330 518.720 1048.730 ;
        RECT 520.710 999.330 520.990 1000.000 ;
        RECT 518.580 999.190 520.990 999.330 ;
        RECT 520.710 996.000 520.990 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3485.880 2901.130 3486.160 ;
      LAYER met3 ;
        RECT 2900.825 3486.170 2901.155 3486.185 ;
        RECT 2917.600 3486.170 2924.800 3486.620 ;
        RECT 2900.825 3485.870 2924.800 3486.170 ;
        RECT 2900.825 3485.855 2901.155 3485.870 ;
        RECT 2917.600 3485.420 2924.800 3485.870 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 1011.005 2636.100 3517.600 ;
        RECT 544.270 1010.635 544.550 1011.005 ;
        RECT 2635.890 1010.635 2636.170 1011.005 ;
        RECT 542.790 999.330 543.070 1000.000 ;
        RECT 544.340 999.330 544.480 1010.635 ;
        RECT 542.790 999.190 544.480 999.330 ;
        RECT 542.790 996.000 543.070 999.190 ;
      LAYER via2 ;
        RECT 544.270 1010.680 544.550 1010.960 ;
        RECT 2635.890 1010.680 2636.170 1010.960 ;
      LAYER met3 ;
        RECT 544.245 1010.970 544.575 1010.985 ;
        RECT 2635.865 1010.970 2636.195 1010.985 ;
        RECT 544.245 1010.670 2636.195 1010.970 ;
        RECT 544.245 1010.655 544.575 1010.670 ;
        RECT 2635.865 1010.655 2636.195 1010.670 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 3501.560 559.290 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 558.970 3501.420 2311.890 3501.560 ;
        RECT 558.970 3501.360 559.290 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
      LAYER via ;
        RECT 559.000 3501.360 559.260 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 559.000 3501.330 559.260 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 559.060 1048.870 559.200 3501.330 ;
        RECT 559.060 1048.730 563.800 1048.870 ;
        RECT 563.660 999.330 563.800 1048.730 ;
        RECT 565.330 999.330 565.610 1000.000 ;
        RECT 563.660 999.190 565.610 999.330 ;
        RECT 565.330 996.000 565.610 999.190 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 3502.240 586.890 3502.300 ;
        RECT 1987.270 3502.240 1987.590 3502.300 ;
        RECT 586.570 3502.100 1987.590 3502.240 ;
        RECT 586.570 3502.040 586.890 3502.100 ;
        RECT 1987.270 3502.040 1987.590 3502.100 ;
      LAYER via ;
        RECT 586.600 3502.040 586.860 3502.300 ;
        RECT 1987.300 3502.040 1987.560 3502.300 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3502.330 1987.500 3517.600 ;
        RECT 586.600 3502.010 586.860 3502.330 ;
        RECT 1987.300 3502.010 1987.560 3502.330 ;
        RECT 586.660 999.330 586.800 3502.010 ;
        RECT 587.410 999.330 587.690 1000.000 ;
        RECT 586.660 999.190 587.690 999.330 ;
        RECT 587.410 996.000 587.690 999.190 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 3502.920 608.050 3502.980 ;
        RECT 1662.510 3502.920 1662.830 3502.980 ;
        RECT 607.730 3502.780 1662.830 3502.920 ;
        RECT 607.730 3502.720 608.050 3502.780 ;
        RECT 1662.510 3502.720 1662.830 3502.780 ;
      LAYER via ;
        RECT 607.760 3502.720 608.020 3502.980 ;
        RECT 1662.540 3502.720 1662.800 3502.980 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.010 1662.740 3517.600 ;
        RECT 607.760 3502.690 608.020 3503.010 ;
        RECT 1662.540 3502.690 1662.800 3503.010 ;
        RECT 607.820 999.330 607.960 3502.690 ;
        RECT 609.490 999.330 609.770 1000.000 ;
        RECT 607.820 999.190 609.770 999.330 ;
        RECT 609.490 996.000 609.770 999.190 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.970 3503.600 628.290 3503.660 ;
        RECT 1338.210 3503.600 1338.530 3503.660 ;
        RECT 627.970 3503.460 1338.530 3503.600 ;
        RECT 627.970 3503.400 628.290 3503.460 ;
        RECT 1338.210 3503.400 1338.530 3503.460 ;
      LAYER via ;
        RECT 628.000 3503.400 628.260 3503.660 ;
        RECT 1338.240 3503.400 1338.500 3503.660 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3503.690 1338.440 3517.600 ;
        RECT 628.000 3503.370 628.260 3503.690 ;
        RECT 1338.240 3503.370 1338.500 3503.690 ;
        RECT 628.060 1048.870 628.200 3503.370 ;
        RECT 628.060 1048.730 630.040 1048.870 ;
        RECT 629.900 999.330 630.040 1048.730 ;
        RECT 631.570 999.330 631.850 1000.000 ;
        RECT 629.900 999.190 631.850 999.330 ;
        RECT 631.570 996.000 631.850 999.190 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 1008.595 235.430 1008.965 ;
        RECT 2899.930 1008.595 2900.210 1008.965 ;
        RECT 233.210 999.330 233.490 1000.000 ;
        RECT 235.220 999.330 235.360 1008.595 ;
        RECT 233.210 999.190 235.360 999.330 ;
        RECT 233.210 996.000 233.490 999.190 ;
        RECT 2900.000 365.005 2900.140 1008.595 ;
        RECT 2899.930 364.635 2900.210 365.005 ;
      LAYER via2 ;
        RECT 235.150 1008.640 235.430 1008.920 ;
        RECT 2899.930 1008.640 2900.210 1008.920 ;
        RECT 2899.930 364.680 2900.210 364.960 ;
      LAYER met3 ;
        RECT 235.125 1008.930 235.455 1008.945 ;
        RECT 2899.905 1008.930 2900.235 1008.945 ;
        RECT 235.125 1008.630 2900.235 1008.930 ;
        RECT 235.125 1008.615 235.455 1008.630 ;
        RECT 2899.905 1008.615 2900.235 1008.630 ;
        RECT 2899.905 364.970 2900.235 364.985 ;
        RECT 2917.600 364.970 2924.800 365.420 ;
        RECT 2899.905 364.670 2924.800 364.970 ;
        RECT 2899.905 364.655 2900.235 364.670 ;
        RECT 2917.600 364.220 2924.800 364.670 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 3501.220 648.990 3501.280 ;
        RECT 1013.910 3501.220 1014.230 3501.280 ;
        RECT 648.670 3501.080 1014.230 3501.220 ;
        RECT 648.670 3501.020 648.990 3501.080 ;
        RECT 1013.910 3501.020 1014.230 3501.080 ;
      LAYER via ;
        RECT 648.700 3501.020 648.960 3501.280 ;
        RECT 1013.940 3501.020 1014.200 3501.280 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3501.310 1014.140 3517.600 ;
        RECT 648.700 3500.990 648.960 3501.310 ;
        RECT 1013.940 3500.990 1014.200 3501.310 ;
        RECT 648.760 1048.870 648.900 3500.990 ;
        RECT 648.760 1048.730 652.120 1048.870 ;
        RECT 651.980 999.330 652.120 1048.730 ;
        RECT 653.650 999.330 653.930 1000.000 ;
        RECT 651.980 999.190 653.930 999.330 ;
        RECT 653.650 996.000 653.930 999.190 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 675.350 1013.780 675.670 1013.840 ;
        RECT 683.170 1013.780 683.490 1013.840 ;
        RECT 675.350 1013.640 683.490 1013.780 ;
        RECT 675.350 1013.580 675.670 1013.640 ;
        RECT 683.170 1013.580 683.490 1013.640 ;
      LAYER via ;
        RECT 675.380 1013.580 675.640 1013.840 ;
        RECT 683.200 1013.580 683.460 1013.840 ;
      LAYER met2 ;
        RECT 683.260 3517.910 688.460 3518.050 ;
        RECT 683.260 1013.870 683.400 3517.910 ;
        RECT 688.320 3517.370 688.460 3517.910 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.320 3517.230 689.380 3517.370 ;
        RECT 675.380 1013.550 675.640 1013.870 ;
        RECT 683.200 1013.550 683.460 1013.870 ;
        RECT 675.440 999.330 675.580 1013.550 ;
        RECT 675.730 999.330 676.010 1000.000 ;
        RECT 675.440 999.190 676.010 999.330 ;
        RECT 675.730 996.000 676.010 999.190 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.850 3500.880 365.170 3500.940 ;
        RECT 693.290 3500.880 693.610 3500.940 ;
        RECT 364.850 3500.740 693.610 3500.880 ;
        RECT 364.850 3500.680 365.170 3500.740 ;
        RECT 693.290 3500.680 693.610 3500.740 ;
        RECT 693.290 1014.120 693.610 1014.180 ;
        RECT 696.970 1014.120 697.290 1014.180 ;
        RECT 693.290 1013.980 697.290 1014.120 ;
        RECT 693.290 1013.920 693.610 1013.980 ;
        RECT 696.970 1013.920 697.290 1013.980 ;
      LAYER via ;
        RECT 364.880 3500.680 365.140 3500.940 ;
        RECT 693.320 3500.680 693.580 3500.940 ;
        RECT 693.320 1013.920 693.580 1014.180 ;
        RECT 697.000 1013.920 697.260 1014.180 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3500.970 365.080 3517.600 ;
        RECT 364.880 3500.650 365.140 3500.970 ;
        RECT 693.320 3500.650 693.580 3500.970 ;
        RECT 693.380 1014.210 693.520 3500.650 ;
        RECT 693.320 1013.890 693.580 1014.210 ;
        RECT 697.000 1013.890 697.260 1014.210 ;
        RECT 697.060 999.330 697.200 1013.890 ;
        RECT 697.810 999.330 698.090 1000.000 ;
        RECT 697.060 999.190 698.090 999.330 ;
        RECT 697.810 996.000 698.090 999.190 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.550 3503.940 40.870 3504.000 ;
        RECT 700.190 3503.940 700.510 3504.000 ;
        RECT 40.550 3503.800 700.510 3503.940 ;
        RECT 40.550 3503.740 40.870 3503.800 ;
        RECT 700.190 3503.740 700.510 3503.800 ;
        RECT 700.190 1012.760 700.510 1012.820 ;
        RECT 718.590 1012.760 718.910 1012.820 ;
        RECT 700.190 1012.620 718.910 1012.760 ;
        RECT 700.190 1012.560 700.510 1012.620 ;
        RECT 718.590 1012.560 718.910 1012.620 ;
      LAYER via ;
        RECT 40.580 3503.740 40.840 3504.000 ;
        RECT 700.220 3503.740 700.480 3504.000 ;
        RECT 700.220 1012.560 700.480 1012.820 ;
        RECT 718.620 1012.560 718.880 1012.820 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3504.030 40.780 3517.600 ;
        RECT 40.580 3503.710 40.840 3504.030 ;
        RECT 700.220 3503.710 700.480 3504.030 ;
        RECT 700.280 1012.850 700.420 3503.710 ;
        RECT 700.220 1012.530 700.480 1012.850 ;
        RECT 718.620 1012.530 718.880 1012.850 ;
        RECT 718.680 999.330 718.820 1012.530 ;
        RECT 719.890 999.330 720.170 1000.000 ;
        RECT 718.680 999.190 720.170 999.330 ;
        RECT 719.890 996.000 720.170 999.190 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3284.640 17.410 3284.700 ;
        RECT 738.370 3284.640 738.690 3284.700 ;
        RECT 17.090 3284.500 738.690 3284.640 ;
        RECT 17.090 3284.440 17.410 3284.500 ;
        RECT 738.370 3284.440 738.690 3284.500 ;
      LAYER via ;
        RECT 17.120 3284.440 17.380 3284.700 ;
        RECT 738.400 3284.440 738.660 3284.700 ;
      LAYER met2 ;
        RECT 17.110 3290.675 17.390 3291.045 ;
        RECT 17.180 3284.730 17.320 3290.675 ;
        RECT 17.120 3284.410 17.380 3284.730 ;
        RECT 738.400 3284.410 738.660 3284.730 ;
        RECT 738.460 1048.870 738.600 3284.410 ;
        RECT 738.460 1048.730 740.440 1048.870 ;
        RECT 740.300 999.330 740.440 1048.730 ;
        RECT 741.970 999.330 742.250 1000.000 ;
        RECT 740.300 999.190 742.250 999.330 ;
        RECT 741.970 996.000 742.250 999.190 ;
      LAYER via2 ;
        RECT 17.110 3290.720 17.390 3291.000 ;
      LAYER met3 ;
        RECT -4.800 3291.010 2.400 3291.460 ;
        RECT 17.085 3291.010 17.415 3291.025 ;
        RECT -4.800 3290.710 17.415 3291.010 ;
        RECT -4.800 3290.260 2.400 3290.710 ;
        RECT 17.085 3290.695 17.415 3290.710 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 3029.300 16.490 3029.360 ;
        RECT 759.070 3029.300 759.390 3029.360 ;
        RECT 16.170 3029.160 759.390 3029.300 ;
        RECT 16.170 3029.100 16.490 3029.160 ;
        RECT 759.070 3029.100 759.390 3029.160 ;
      LAYER via ;
        RECT 16.200 3029.100 16.460 3029.360 ;
        RECT 759.100 3029.100 759.360 3029.360 ;
      LAYER met2 ;
        RECT 16.190 3030.235 16.470 3030.605 ;
        RECT 16.260 3029.390 16.400 3030.235 ;
        RECT 16.200 3029.070 16.460 3029.390 ;
        RECT 759.100 3029.070 759.360 3029.390 ;
        RECT 759.160 1048.870 759.300 3029.070 ;
        RECT 759.160 1048.730 762.520 1048.870 ;
        RECT 762.380 999.330 762.520 1048.730 ;
        RECT 764.510 999.330 764.790 1000.000 ;
        RECT 762.380 999.190 764.790 999.330 ;
        RECT 764.510 996.000 764.790 999.190 ;
      LAYER via2 ;
        RECT 16.190 3030.280 16.470 3030.560 ;
      LAYER met3 ;
        RECT -4.800 3030.570 2.400 3031.020 ;
        RECT 16.165 3030.570 16.495 3030.585 ;
        RECT -4.800 3030.270 16.495 3030.570 ;
        RECT -4.800 3029.820 2.400 3030.270 ;
        RECT 16.165 3030.255 16.495 3030.270 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2767.160 17.410 2767.220 ;
        RECT 786.670 2767.160 786.990 2767.220 ;
        RECT 17.090 2767.020 786.990 2767.160 ;
        RECT 17.090 2766.960 17.410 2767.020 ;
        RECT 786.670 2766.960 786.990 2767.020 ;
      LAYER via ;
        RECT 17.120 2766.960 17.380 2767.220 ;
        RECT 786.700 2766.960 786.960 2767.220 ;
      LAYER met2 ;
        RECT 17.110 2769.115 17.390 2769.485 ;
        RECT 17.180 2767.250 17.320 2769.115 ;
        RECT 17.120 2766.930 17.380 2767.250 ;
        RECT 786.700 2766.930 786.960 2767.250 ;
        RECT 786.760 1048.870 786.900 2766.930 ;
        RECT 786.760 1048.730 787.360 1048.870 ;
        RECT 786.590 999.330 786.870 1000.000 ;
        RECT 787.220 999.330 787.360 1048.730 ;
        RECT 786.590 999.190 787.360 999.330 ;
        RECT 786.590 996.000 786.870 999.190 ;
      LAYER via2 ;
        RECT 17.110 2769.160 17.390 2769.440 ;
      LAYER met3 ;
        RECT -4.800 2769.450 2.400 2769.900 ;
        RECT 17.085 2769.450 17.415 2769.465 ;
        RECT -4.800 2769.150 17.415 2769.450 ;
        RECT -4.800 2768.700 2.400 2769.150 ;
        RECT 17.085 2769.135 17.415 2769.150 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2505.020 15.570 2505.080 ;
        RECT 807.370 2505.020 807.690 2505.080 ;
        RECT 15.250 2504.880 807.690 2505.020 ;
        RECT 15.250 2504.820 15.570 2504.880 ;
        RECT 807.370 2504.820 807.690 2504.880 ;
      LAYER via ;
        RECT 15.280 2504.820 15.540 2505.080 ;
        RECT 807.400 2504.820 807.660 2505.080 ;
      LAYER met2 ;
        RECT 15.270 2508.675 15.550 2509.045 ;
        RECT 15.340 2505.110 15.480 2508.675 ;
        RECT 15.280 2504.790 15.540 2505.110 ;
        RECT 807.400 2504.790 807.660 2505.110 ;
        RECT 807.460 999.330 807.600 2504.790 ;
        RECT 808.670 999.330 808.950 1000.000 ;
        RECT 807.460 999.190 808.950 999.330 ;
        RECT 808.670 996.000 808.950 999.190 ;
      LAYER via2 ;
        RECT 15.270 2508.720 15.550 2509.000 ;
      LAYER met3 ;
        RECT -4.800 2509.010 2.400 2509.460 ;
        RECT 15.245 2509.010 15.575 2509.025 ;
        RECT -4.800 2508.710 15.575 2509.010 ;
        RECT -4.800 2508.260 2.400 2508.710 ;
        RECT 15.245 2508.695 15.575 2508.710 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2242.880 16.030 2242.940 ;
        RECT 828.070 2242.880 828.390 2242.940 ;
        RECT 15.710 2242.740 828.390 2242.880 ;
        RECT 15.710 2242.680 16.030 2242.740 ;
        RECT 828.070 2242.680 828.390 2242.740 ;
      LAYER via ;
        RECT 15.740 2242.680 16.000 2242.940 ;
        RECT 828.100 2242.680 828.360 2242.940 ;
      LAYER met2 ;
        RECT 15.730 2247.555 16.010 2247.925 ;
        RECT 15.800 2242.970 15.940 2247.555 ;
        RECT 15.740 2242.650 16.000 2242.970 ;
        RECT 828.100 2242.650 828.360 2242.970 ;
        RECT 828.160 1048.870 828.300 2242.650 ;
        RECT 828.160 1048.730 828.760 1048.870 ;
        RECT 828.620 999.330 828.760 1048.730 ;
        RECT 830.750 999.330 831.030 1000.000 ;
        RECT 828.620 999.190 831.030 999.330 ;
        RECT 830.750 996.000 831.030 999.190 ;
      LAYER via2 ;
        RECT 15.730 2247.600 16.010 2247.880 ;
      LAYER met3 ;
        RECT -4.800 2247.890 2.400 2248.340 ;
        RECT 15.705 2247.890 16.035 2247.905 ;
        RECT -4.800 2247.590 16.035 2247.890 ;
        RECT -4.800 2247.140 2.400 2247.590 ;
        RECT 15.705 2247.575 16.035 2247.590 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 1987.540 17.410 1987.600 ;
        RECT 849.230 1987.540 849.550 1987.600 ;
        RECT 17.090 1987.400 849.550 1987.540 ;
        RECT 17.090 1987.340 17.410 1987.400 ;
        RECT 849.230 1987.340 849.550 1987.400 ;
      LAYER via ;
        RECT 17.120 1987.340 17.380 1987.600 ;
        RECT 849.260 1987.340 849.520 1987.600 ;
      LAYER met2 ;
        RECT 17.120 1987.485 17.380 1987.630 ;
        RECT 17.110 1987.115 17.390 1987.485 ;
        RECT 849.260 1987.310 849.520 1987.630 ;
        RECT 849.320 1048.870 849.460 1987.310 ;
        RECT 849.320 1048.730 850.840 1048.870 ;
        RECT 850.700 999.330 850.840 1048.730 ;
        RECT 852.830 999.330 853.110 1000.000 ;
        RECT 850.700 999.190 853.110 999.330 ;
        RECT 852.830 996.000 853.110 999.190 ;
      LAYER via2 ;
        RECT 17.110 1987.160 17.390 1987.440 ;
      LAYER met3 ;
        RECT -4.800 1987.450 2.400 1987.900 ;
        RECT 17.085 1987.450 17.415 1987.465 ;
        RECT -4.800 1987.150 17.415 1987.450 ;
        RECT -4.800 1986.700 2.400 1987.150 ;
        RECT 17.085 1987.135 17.415 1987.150 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1101.310 565.660 1101.630 565.720 ;
        RECT 2899.450 565.660 2899.770 565.720 ;
        RECT 1101.310 565.520 2899.770 565.660 ;
        RECT 1101.310 565.460 1101.630 565.520 ;
        RECT 2899.450 565.460 2899.770 565.520 ;
      LAYER via ;
        RECT 1101.340 565.460 1101.600 565.720 ;
        RECT 2899.480 565.460 2899.740 565.720 ;
      LAYER met2 ;
        RECT 257.230 1009.955 257.510 1010.325 ;
        RECT 1101.330 1009.955 1101.610 1010.325 ;
        RECT 255.290 999.330 255.570 1000.000 ;
        RECT 257.300 999.330 257.440 1009.955 ;
        RECT 255.290 999.190 257.440 999.330 ;
        RECT 255.290 996.000 255.570 999.190 ;
        RECT 1101.400 565.750 1101.540 1009.955 ;
        RECT 1101.340 565.430 1101.600 565.750 ;
        RECT 2899.480 565.430 2899.740 565.750 ;
        RECT 2899.540 564.245 2899.680 565.430 ;
        RECT 2899.470 563.875 2899.750 564.245 ;
      LAYER via2 ;
        RECT 257.230 1010.000 257.510 1010.280 ;
        RECT 1101.330 1010.000 1101.610 1010.280 ;
        RECT 2899.470 563.920 2899.750 564.200 ;
      LAYER met3 ;
        RECT 257.205 1010.290 257.535 1010.305 ;
        RECT 1101.305 1010.290 1101.635 1010.305 ;
        RECT 257.205 1009.990 1101.635 1010.290 ;
        RECT 257.205 1009.975 257.535 1009.990 ;
        RECT 1101.305 1009.975 1101.635 1009.990 ;
        RECT 2899.445 564.210 2899.775 564.225 ;
        RECT 2917.600 564.210 2924.800 564.660 ;
        RECT 2899.445 563.910 2924.800 564.210 ;
        RECT 2899.445 563.895 2899.775 563.910 ;
        RECT 2917.600 563.460 2924.800 563.910 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1725.400 16.950 1725.460 ;
        RECT 869.470 1725.400 869.790 1725.460 ;
        RECT 16.630 1725.260 869.790 1725.400 ;
        RECT 16.630 1725.200 16.950 1725.260 ;
        RECT 869.470 1725.200 869.790 1725.260 ;
      LAYER via ;
        RECT 16.660 1725.200 16.920 1725.460 ;
        RECT 869.500 1725.200 869.760 1725.460 ;
      LAYER met2 ;
        RECT 16.650 1726.675 16.930 1727.045 ;
        RECT 16.720 1725.490 16.860 1726.675 ;
        RECT 16.660 1725.170 16.920 1725.490 ;
        RECT 869.500 1725.170 869.760 1725.490 ;
        RECT 869.560 1048.870 869.700 1725.170 ;
        RECT 869.560 1048.730 872.920 1048.870 ;
        RECT 872.780 999.330 872.920 1048.730 ;
        RECT 874.910 999.330 875.190 1000.000 ;
        RECT 872.780 999.190 875.190 999.330 ;
        RECT 874.910 996.000 875.190 999.190 ;
      LAYER via2 ;
        RECT 16.650 1726.720 16.930 1727.000 ;
      LAYER met3 ;
        RECT -4.800 1727.010 2.400 1727.460 ;
        RECT 16.625 1727.010 16.955 1727.025 ;
        RECT -4.800 1726.710 16.955 1727.010 ;
        RECT -4.800 1726.260 2.400 1726.710 ;
        RECT 16.625 1726.695 16.955 1726.710 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1462.920 17.870 1462.980 ;
        RECT 897.070 1462.920 897.390 1462.980 ;
        RECT 17.550 1462.780 897.390 1462.920 ;
        RECT 17.550 1462.720 17.870 1462.780 ;
        RECT 897.070 1462.720 897.390 1462.780 ;
      LAYER via ;
        RECT 17.580 1462.720 17.840 1462.980 ;
        RECT 897.100 1462.720 897.360 1462.980 ;
      LAYER met2 ;
        RECT 17.570 1465.555 17.850 1465.925 ;
        RECT 17.640 1463.010 17.780 1465.555 ;
        RECT 17.580 1462.690 17.840 1463.010 ;
        RECT 897.100 1462.690 897.360 1463.010 ;
        RECT 897.160 1048.870 897.300 1462.690 ;
        RECT 897.160 1048.730 897.760 1048.870 ;
        RECT 896.990 999.330 897.270 1000.000 ;
        RECT 897.620 999.330 897.760 1048.730 ;
        RECT 896.990 999.190 897.760 999.330 ;
        RECT 896.990 996.000 897.270 999.190 ;
      LAYER via2 ;
        RECT 17.570 1465.600 17.850 1465.880 ;
      LAYER met3 ;
        RECT -4.800 1465.890 2.400 1466.340 ;
        RECT 17.545 1465.890 17.875 1465.905 ;
        RECT -4.800 1465.590 17.875 1465.890 ;
        RECT -4.800 1465.140 2.400 1465.590 ;
        RECT 17.545 1465.575 17.875 1465.590 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1200.780 15.570 1200.840 ;
        RECT 917.770 1200.780 918.090 1200.840 ;
        RECT 15.250 1200.640 918.090 1200.780 ;
        RECT 15.250 1200.580 15.570 1200.640 ;
        RECT 917.770 1200.580 918.090 1200.640 ;
      LAYER via ;
        RECT 15.280 1200.580 15.540 1200.840 ;
        RECT 917.800 1200.580 918.060 1200.840 ;
      LAYER met2 ;
        RECT 15.270 1205.115 15.550 1205.485 ;
        RECT 15.340 1200.870 15.480 1205.115 ;
        RECT 15.280 1200.550 15.540 1200.870 ;
        RECT 917.800 1200.550 918.060 1200.870 ;
        RECT 917.860 999.330 918.000 1200.550 ;
        RECT 919.070 999.330 919.350 1000.000 ;
        RECT 917.860 999.190 919.350 999.330 ;
        RECT 919.070 996.000 919.350 999.190 ;
      LAYER via2 ;
        RECT 15.270 1205.160 15.550 1205.440 ;
      LAYER met3 ;
        RECT -4.800 1205.450 2.400 1205.900 ;
        RECT 15.245 1205.450 15.575 1205.465 ;
        RECT -4.800 1205.150 15.575 1205.450 ;
        RECT -4.800 1204.700 2.400 1205.150 ;
        RECT 15.245 1205.135 15.575 1205.150 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1010.380 15.570 1010.440 ;
        RECT 940.310 1010.380 940.630 1010.440 ;
        RECT 15.250 1010.240 940.630 1010.380 ;
        RECT 15.250 1010.180 15.570 1010.240 ;
        RECT 940.310 1010.180 940.630 1010.240 ;
      LAYER via ;
        RECT 15.280 1010.180 15.540 1010.440 ;
        RECT 940.340 1010.180 940.600 1010.440 ;
      LAYER met2 ;
        RECT 15.280 1010.150 15.540 1010.470 ;
        RECT 940.340 1010.150 940.600 1010.470 ;
        RECT 15.340 944.365 15.480 1010.150 ;
        RECT 940.400 999.330 940.540 1010.150 ;
        RECT 941.610 999.330 941.890 1000.000 ;
        RECT 940.400 999.190 941.890 999.330 ;
        RECT 941.610 996.000 941.890 999.190 ;
        RECT 15.270 943.995 15.550 944.365 ;
      LAYER via2 ;
        RECT 15.270 944.040 15.550 944.320 ;
      LAYER met3 ;
        RECT -4.800 944.330 2.400 944.780 ;
        RECT 15.245 944.330 15.575 944.345 ;
        RECT -4.800 944.030 15.575 944.330 ;
        RECT -4.800 943.580 2.400 944.030 ;
        RECT 15.245 944.015 15.575 944.030 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1009.360 16.950 1009.420 ;
        RECT 962.390 1009.360 962.710 1009.420 ;
        RECT 16.630 1009.220 962.710 1009.360 ;
        RECT 16.630 1009.160 16.950 1009.220 ;
        RECT 962.390 1009.160 962.710 1009.220 ;
      LAYER via ;
        RECT 16.660 1009.160 16.920 1009.420 ;
        RECT 962.420 1009.160 962.680 1009.420 ;
      LAYER met2 ;
        RECT 16.660 1009.130 16.920 1009.450 ;
        RECT 962.420 1009.130 962.680 1009.450 ;
        RECT 16.720 683.925 16.860 1009.130 ;
        RECT 962.480 999.330 962.620 1009.130 ;
        RECT 963.690 999.330 963.970 1000.000 ;
        RECT 962.480 999.190 963.970 999.330 ;
        RECT 963.690 996.000 963.970 999.190 ;
        RECT 16.650 683.555 16.930 683.925 ;
      LAYER via2 ;
        RECT 16.650 683.600 16.930 683.880 ;
      LAYER met3 ;
        RECT -4.800 683.890 2.400 684.340 ;
        RECT 16.625 683.890 16.955 683.905 ;
        RECT -4.800 683.590 16.955 683.890 ;
        RECT -4.800 683.140 2.400 683.590 ;
        RECT 16.625 683.575 16.955 683.590 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 1008.680 19.250 1008.740 ;
        RECT 984.470 1008.680 984.790 1008.740 ;
        RECT 18.930 1008.540 984.790 1008.680 ;
        RECT 18.930 1008.480 19.250 1008.540 ;
        RECT 984.470 1008.480 984.790 1008.540 ;
      LAYER via ;
        RECT 18.960 1008.480 19.220 1008.740 ;
        RECT 984.500 1008.480 984.760 1008.740 ;
      LAYER met2 ;
        RECT 18.960 1008.450 19.220 1008.770 ;
        RECT 984.500 1008.450 984.760 1008.770 ;
        RECT 19.020 423.485 19.160 1008.450 ;
        RECT 984.560 999.330 984.700 1008.450 ;
        RECT 985.770 999.330 986.050 1000.000 ;
        RECT 984.560 999.190 986.050 999.330 ;
        RECT 985.770 996.000 986.050 999.190 ;
        RECT 18.950 423.115 19.230 423.485 ;
      LAYER via2 ;
        RECT 18.950 423.160 19.230 423.440 ;
      LAYER met3 ;
        RECT -4.800 423.450 2.400 423.900 ;
        RECT 18.925 423.450 19.255 423.465 ;
        RECT -4.800 423.150 19.255 423.450 ;
        RECT -4.800 422.700 2.400 423.150 ;
        RECT 18.925 423.135 19.255 423.150 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 217.650 999.160 217.970 999.220 ;
        RECT 243.410 999.160 243.730 999.220 ;
        RECT 217.650 999.020 243.730 999.160 ;
        RECT 217.650 998.960 217.970 999.020 ;
        RECT 243.410 998.960 243.730 999.020 ;
        RECT 217.650 997.460 217.970 997.520 ;
        RECT 213.830 997.320 217.970 997.460 ;
        RECT 18.010 994.400 18.330 994.460 ;
        RECT 18.010 994.260 131.170 994.400 ;
        RECT 18.010 994.200 18.330 994.260 ;
        RECT 131.030 993.720 131.170 994.260 ;
        RECT 131.030 993.580 200.170 993.720 ;
        RECT 200.030 993.380 200.170 993.580 ;
        RECT 213.830 993.380 213.970 997.320 ;
        RECT 217.650 997.260 217.970 997.320 ;
        RECT 243.410 997.260 243.730 997.520 ;
        RECT 1008.850 997.260 1009.170 997.520 ;
        RECT 243.500 997.120 243.640 997.260 ;
        RECT 243.500 996.980 262.270 997.120 ;
        RECT 262.130 996.100 262.270 996.980 ;
        RECT 262.130 995.960 269.170 996.100 ;
        RECT 269.030 995.420 269.170 995.960 ;
        RECT 275.930 995.960 281.360 996.100 ;
        RECT 275.930 995.420 276.070 995.960 ;
        RECT 281.220 995.760 281.360 995.960 ;
        RECT 281.220 995.620 282.970 995.760 ;
        RECT 269.030 995.280 276.070 995.420 ;
        RECT 282.830 995.080 282.970 995.620 ;
        RECT 282.830 994.940 284.120 995.080 ;
        RECT 283.980 994.740 284.120 994.940 ;
        RECT 283.980 994.600 285.960 994.740 ;
        RECT 285.820 994.400 285.960 994.600 ;
        RECT 1008.940 994.400 1009.080 997.260 ;
        RECT 285.820 994.260 1009.080 994.400 ;
        RECT 200.030 993.240 213.970 993.380 ;
      LAYER via ;
        RECT 217.680 998.960 217.940 999.220 ;
        RECT 243.440 998.960 243.700 999.220 ;
        RECT 18.040 994.200 18.300 994.460 ;
        RECT 217.680 997.260 217.940 997.520 ;
        RECT 243.440 997.260 243.700 997.520 ;
        RECT 1008.880 997.260 1009.140 997.520 ;
      LAYER met2 ;
        RECT 217.680 998.930 217.940 999.250 ;
        RECT 243.440 998.930 243.700 999.250 ;
        RECT 217.740 997.550 217.880 998.930 ;
        RECT 243.500 997.550 243.640 998.930 ;
        RECT 217.680 997.230 217.940 997.550 ;
        RECT 243.440 997.230 243.700 997.550 ;
        RECT 1007.850 997.290 1008.130 1000.000 ;
        RECT 1008.880 997.290 1009.140 997.550 ;
        RECT 1007.850 997.230 1009.140 997.290 ;
        RECT 1007.850 997.150 1009.080 997.230 ;
        RECT 1007.850 996.000 1008.130 997.150 ;
        RECT 18.040 994.170 18.300 994.490 ;
        RECT 18.100 227.645 18.240 994.170 ;
        RECT 18.030 227.275 18.310 227.645 ;
      LAYER via2 ;
        RECT 18.030 227.320 18.310 227.600 ;
      LAYER met3 ;
        RECT -4.800 227.610 2.400 228.060 ;
        RECT 18.005 227.610 18.335 227.625 ;
        RECT -4.800 227.310 18.335 227.610 ;
        RECT -4.800 226.860 2.400 227.310 ;
        RECT 18.005 227.295 18.335 227.310 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 1009.275 1028.930 1009.645 ;
        RECT 1028.720 999.330 1028.860 1009.275 ;
        RECT 1029.930 999.330 1030.210 1000.000 ;
        RECT 1028.720 999.190 1030.210 999.330 ;
        RECT 1029.930 996.000 1030.210 999.190 ;
      LAYER via2 ;
        RECT 1028.650 1009.320 1028.930 1009.600 ;
      LAYER met3 ;
        RECT 1028.625 1009.610 1028.955 1009.625 ;
        RECT 34.350 1009.310 1028.955 1009.610 ;
        RECT 19.590 1008.930 19.970 1008.940 ;
        RECT 34.350 1008.930 34.650 1009.310 ;
        RECT 1028.625 1009.295 1028.955 1009.310 ;
        RECT 19.590 1008.630 34.650 1008.930 ;
        RECT 19.590 1008.620 19.970 1008.630 ;
        RECT -4.800 32.450 2.400 32.900 ;
        RECT 19.590 32.450 19.970 32.460 ;
        RECT -4.800 32.150 19.970 32.450 ;
        RECT -4.800 31.700 2.400 32.150 ;
        RECT 19.590 32.140 19.970 32.150 ;
      LAYER via3 ;
        RECT 19.620 1008.620 19.940 1008.940 ;
        RECT 19.620 32.140 19.940 32.460 ;
      LAYER met4 ;
        RECT 19.615 1008.615 19.945 1008.945 ;
        RECT 19.630 32.465 19.930 1008.615 ;
        RECT 19.615 32.135 19.945 32.465 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 279.290 1010.720 279.610 1010.780 ;
        RECT 1101.770 1010.720 1102.090 1010.780 ;
        RECT 279.290 1010.580 1102.090 1010.720 ;
        RECT 279.290 1010.520 279.610 1010.580 ;
        RECT 1101.770 1010.520 1102.090 1010.580 ;
        RECT 1101.770 765.920 1102.090 765.980 ;
        RECT 2899.450 765.920 2899.770 765.980 ;
        RECT 1101.770 765.780 2899.770 765.920 ;
        RECT 1101.770 765.720 1102.090 765.780 ;
        RECT 2899.450 765.720 2899.770 765.780 ;
      LAYER via ;
        RECT 279.320 1010.520 279.580 1010.780 ;
        RECT 1101.800 1010.520 1102.060 1010.780 ;
        RECT 1101.800 765.720 1102.060 765.980 ;
        RECT 2899.480 765.720 2899.740 765.980 ;
      LAYER met2 ;
        RECT 279.320 1010.490 279.580 1010.810 ;
        RECT 1101.800 1010.490 1102.060 1010.810 ;
        RECT 277.370 999.330 277.650 1000.000 ;
        RECT 279.380 999.330 279.520 1010.490 ;
        RECT 277.370 999.190 279.520 999.330 ;
        RECT 277.370 996.000 277.650 999.190 ;
        RECT 1101.860 766.010 1102.000 1010.490 ;
        RECT 1101.800 765.690 1102.060 766.010 ;
        RECT 2899.480 765.690 2899.740 766.010 ;
        RECT 2899.540 763.485 2899.680 765.690 ;
        RECT 2899.470 763.115 2899.750 763.485 ;
      LAYER via2 ;
        RECT 2899.470 763.160 2899.750 763.440 ;
      LAYER met3 ;
        RECT 2899.445 763.450 2899.775 763.465 ;
        RECT 2917.600 763.450 2924.800 763.900 ;
        RECT 2899.445 763.150 2924.800 763.450 ;
        RECT 2899.445 763.135 2899.775 763.150 ;
        RECT 2917.600 762.700 2924.800 763.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.370 1012.080 301.690 1012.140 ;
        RECT 1103.150 1012.080 1103.470 1012.140 ;
        RECT 301.370 1011.940 1103.470 1012.080 ;
        RECT 301.370 1011.880 301.690 1011.940 ;
        RECT 1103.150 1011.880 1103.470 1011.940 ;
        RECT 1103.150 965.840 1103.470 965.900 ;
        RECT 2899.450 965.840 2899.770 965.900 ;
        RECT 1103.150 965.700 2899.770 965.840 ;
        RECT 1103.150 965.640 1103.470 965.700 ;
        RECT 2899.450 965.640 2899.770 965.700 ;
      LAYER via ;
        RECT 301.400 1011.880 301.660 1012.140 ;
        RECT 1103.180 1011.880 1103.440 1012.140 ;
        RECT 1103.180 965.640 1103.440 965.900 ;
        RECT 2899.480 965.640 2899.740 965.900 ;
      LAYER met2 ;
        RECT 301.400 1011.850 301.660 1012.170 ;
        RECT 1103.180 1011.850 1103.440 1012.170 ;
        RECT 299.450 999.330 299.730 1000.000 ;
        RECT 301.460 999.330 301.600 1011.850 ;
        RECT 299.450 999.190 301.600 999.330 ;
        RECT 299.450 996.000 299.730 999.190 ;
        RECT 1103.240 965.930 1103.380 1011.850 ;
        RECT 1103.180 965.610 1103.440 965.930 ;
        RECT 2899.480 965.610 2899.740 965.930 ;
        RECT 2899.540 962.725 2899.680 965.610 ;
        RECT 2899.470 962.355 2899.750 962.725 ;
      LAYER via2 ;
        RECT 2899.470 962.400 2899.750 962.680 ;
      LAYER met3 ;
        RECT 2899.445 962.690 2899.775 962.705 ;
        RECT 2917.600 962.690 2924.800 963.140 ;
        RECT 2899.445 962.390 2924.800 962.690 ;
        RECT 2899.445 962.375 2899.775 962.390 ;
        RECT 2917.600 961.940 2924.800 962.390 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.470 1159.300 317.790 1159.360 ;
        RECT 2898.990 1159.300 2899.310 1159.360 ;
        RECT 317.470 1159.160 2899.310 1159.300 ;
        RECT 317.470 1159.100 317.790 1159.160 ;
        RECT 2898.990 1159.100 2899.310 1159.160 ;
      LAYER via ;
        RECT 317.500 1159.100 317.760 1159.360 ;
        RECT 2899.020 1159.100 2899.280 1159.360 ;
      LAYER met2 ;
        RECT 2899.010 1161.595 2899.290 1161.965 ;
        RECT 2899.080 1159.390 2899.220 1161.595 ;
        RECT 317.500 1159.070 317.760 1159.390 ;
        RECT 2899.020 1159.070 2899.280 1159.390 ;
        RECT 317.560 1048.870 317.700 1159.070 ;
        RECT 317.560 1048.730 320.000 1048.870 ;
        RECT 319.860 999.330 320.000 1048.730 ;
        RECT 321.530 999.330 321.810 1000.000 ;
        RECT 319.860 999.190 321.810 999.330 ;
        RECT 321.530 996.000 321.810 999.190 ;
      LAYER via2 ;
        RECT 2899.010 1161.640 2899.290 1161.920 ;
      LAYER met3 ;
        RECT 2898.985 1161.930 2899.315 1161.945 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2898.985 1161.630 2924.800 1161.930 ;
        RECT 2898.985 1161.615 2899.315 1161.630 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 338.170 1359.560 338.490 1359.620 ;
        RECT 2900.830 1359.560 2901.150 1359.620 ;
        RECT 338.170 1359.420 2901.150 1359.560 ;
        RECT 338.170 1359.360 338.490 1359.420 ;
        RECT 2900.830 1359.360 2901.150 1359.420 ;
      LAYER via ;
        RECT 338.200 1359.360 338.460 1359.620 ;
        RECT 2900.860 1359.360 2901.120 1359.620 ;
      LAYER met2 ;
        RECT 2900.850 1360.835 2901.130 1361.205 ;
        RECT 2900.920 1359.650 2901.060 1360.835 ;
        RECT 338.200 1359.330 338.460 1359.650 ;
        RECT 2900.860 1359.330 2901.120 1359.650 ;
        RECT 338.260 1048.870 338.400 1359.330 ;
        RECT 338.260 1048.730 342.080 1048.870 ;
        RECT 341.940 999.330 342.080 1048.730 ;
        RECT 343.610 999.330 343.890 1000.000 ;
        RECT 341.940 999.190 343.890 999.330 ;
        RECT 343.610 996.000 343.890 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1360.880 2901.130 1361.160 ;
      LAYER met3 ;
        RECT 2900.825 1361.170 2901.155 1361.185 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2900.825 1360.870 2924.800 1361.170 ;
        RECT 2900.825 1360.855 2901.155 1360.870 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 1621.700 366.090 1621.760 ;
        RECT 2899.910 1621.700 2900.230 1621.760 ;
        RECT 365.770 1621.560 2900.230 1621.700 ;
        RECT 365.770 1621.500 366.090 1621.560 ;
        RECT 2899.910 1621.500 2900.230 1621.560 ;
      LAYER via ;
        RECT 365.800 1621.500 366.060 1621.760 ;
        RECT 2899.940 1621.500 2900.200 1621.760 ;
      LAYER met2 ;
        RECT 2899.930 1626.035 2900.210 1626.405 ;
        RECT 2900.000 1621.790 2900.140 1626.035 ;
        RECT 365.800 1621.470 366.060 1621.790 ;
        RECT 2899.940 1621.470 2900.200 1621.790 ;
        RECT 365.860 1048.870 366.000 1621.470 ;
        RECT 365.860 1048.730 366.460 1048.870 ;
        RECT 365.690 999.330 365.970 1000.000 ;
        RECT 366.320 999.330 366.460 1048.730 ;
        RECT 365.690 999.190 366.460 999.330 ;
        RECT 365.690 996.000 365.970 999.190 ;
      LAYER via2 ;
        RECT 2899.930 1626.080 2900.210 1626.360 ;
      LAYER met3 ;
        RECT 2899.905 1626.370 2900.235 1626.385 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2899.905 1626.070 2924.800 1626.370 ;
        RECT 2899.905 1626.055 2900.235 1626.070 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.470 1890.980 386.790 1891.040 ;
        RECT 2900.830 1890.980 2901.150 1891.040 ;
        RECT 386.470 1890.840 2901.150 1890.980 ;
        RECT 386.470 1890.780 386.790 1890.840 ;
        RECT 2900.830 1890.780 2901.150 1890.840 ;
      LAYER via ;
        RECT 386.500 1890.780 386.760 1891.040 ;
        RECT 2900.860 1890.780 2901.120 1891.040 ;
      LAYER met2 ;
        RECT 2900.850 1891.915 2901.130 1892.285 ;
        RECT 2900.920 1891.070 2901.060 1891.915 ;
        RECT 386.500 1890.750 386.760 1891.070 ;
        RECT 2900.860 1890.750 2901.120 1891.070 ;
        RECT 386.560 999.330 386.700 1890.750 ;
        RECT 388.230 999.330 388.510 1000.000 ;
        RECT 386.560 999.190 388.510 999.330 ;
        RECT 388.230 996.000 388.510 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1891.960 2901.130 1892.240 ;
      LAYER met3 ;
        RECT 2900.825 1892.250 2901.155 1892.265 ;
        RECT 2917.600 1892.250 2924.800 1892.700 ;
        RECT 2900.825 1891.950 2924.800 1892.250 ;
        RECT 2900.825 1891.935 2901.155 1891.950 ;
        RECT 2917.600 1891.500 2924.800 1891.950 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 2153.120 407.490 2153.180 ;
        RECT 2900.830 2153.120 2901.150 2153.180 ;
        RECT 407.170 2152.980 2901.150 2153.120 ;
        RECT 407.170 2152.920 407.490 2152.980 ;
        RECT 2900.830 2152.920 2901.150 2152.980 ;
      LAYER via ;
        RECT 407.200 2152.920 407.460 2153.180 ;
        RECT 2900.860 2152.920 2901.120 2153.180 ;
      LAYER met2 ;
        RECT 2900.850 2157.795 2901.130 2158.165 ;
        RECT 2900.920 2153.210 2901.060 2157.795 ;
        RECT 407.200 2152.890 407.460 2153.210 ;
        RECT 2900.860 2152.890 2901.120 2153.210 ;
        RECT 407.260 1048.870 407.400 2152.890 ;
        RECT 407.260 1048.730 408.320 1048.870 ;
        RECT 408.180 999.330 408.320 1048.730 ;
        RECT 410.310 999.330 410.590 1000.000 ;
        RECT 408.180 999.190 410.590 999.330 ;
        RECT 410.310 996.000 410.590 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2157.840 2901.130 2158.120 ;
      LAYER met3 ;
        RECT 2900.825 2158.130 2901.155 2158.145 ;
        RECT 2917.600 2158.130 2924.800 2158.580 ;
        RECT 2900.825 2157.830 2924.800 2158.130 ;
        RECT 2900.825 2157.815 2901.155 2157.830 ;
        RECT 2917.600 2157.380 2924.800 2157.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.410 997.260 220.730 997.520 ;
        RECT 220.500 993.040 220.640 997.260 ;
        RECT 2903.590 993.720 2903.910 993.780 ;
        RECT 358.730 993.580 2903.910 993.720 ;
        RECT 220.500 992.900 262.270 993.040 ;
        RECT 262.130 992.360 262.270 992.900 ;
        RECT 282.830 992.900 289.870 993.040 ;
        RECT 282.830 992.700 282.970 992.900 ;
        RECT 275.930 992.560 282.970 992.700 ;
        RECT 275.930 992.360 276.070 992.560 ;
        RECT 262.130 992.220 276.070 992.360 ;
        RECT 289.730 992.360 289.870 992.900 ;
        RECT 358.730 992.360 358.870 993.580 ;
        RECT 2903.590 993.520 2903.910 993.580 ;
        RECT 289.730 992.220 296.770 992.360 ;
        RECT 296.630 992.020 296.770 992.220 ;
        RECT 337.800 992.220 358.870 992.360 ;
        RECT 337.800 992.020 337.940 992.220 ;
        RECT 296.630 991.880 337.940 992.020 ;
      LAYER via ;
        RECT 220.440 997.260 220.700 997.520 ;
        RECT 2903.620 993.520 2903.880 993.780 ;
      LAYER met2 ;
        RECT 218.490 997.290 218.770 1000.000 ;
        RECT 220.440 997.290 220.700 997.550 ;
        RECT 218.490 997.230 220.700 997.290 ;
        RECT 218.490 997.150 220.640 997.230 ;
        RECT 218.490 996.000 218.770 997.150 ;
        RECT 2903.620 993.490 2903.880 993.810 ;
        RECT 2903.680 99.125 2903.820 993.490 ;
        RECT 2903.610 98.755 2903.890 99.125 ;
      LAYER via2 ;
        RECT 2903.610 98.800 2903.890 99.080 ;
      LAYER met3 ;
        RECT 2903.585 99.090 2903.915 99.105 ;
        RECT 2917.600 99.090 2924.800 99.540 ;
        RECT 2903.585 98.790 2924.800 99.090 ;
        RECT 2903.585 98.775 2903.915 98.790 ;
        RECT 2917.600 98.340 2924.800 98.790 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 2353.040 435.090 2353.100 ;
        RECT 2898.070 2353.040 2898.390 2353.100 ;
        RECT 434.770 2352.900 2898.390 2353.040 ;
        RECT 434.770 2352.840 435.090 2352.900 ;
        RECT 2898.070 2352.840 2898.390 2352.900 ;
      LAYER via ;
        RECT 434.800 2352.840 435.060 2353.100 ;
        RECT 2898.100 2352.840 2898.360 2353.100 ;
      LAYER met2 ;
        RECT 2898.090 2357.035 2898.370 2357.405 ;
        RECT 2898.160 2353.130 2898.300 2357.035 ;
        RECT 434.800 2352.810 435.060 2353.130 ;
        RECT 2898.100 2352.810 2898.360 2353.130 ;
        RECT 434.860 1048.870 435.000 2352.810 ;
        RECT 434.860 1048.730 437.760 1048.870 ;
        RECT 437.620 999.330 437.760 1048.730 ;
        RECT 439.750 999.330 440.030 1000.000 ;
        RECT 437.620 999.190 440.030 999.330 ;
        RECT 439.750 996.000 440.030 999.190 ;
      LAYER via2 ;
        RECT 2898.090 2357.080 2898.370 2357.360 ;
      LAYER met3 ;
        RECT 2898.065 2357.370 2898.395 2357.385 ;
        RECT 2917.600 2357.370 2924.800 2357.820 ;
        RECT 2898.065 2357.070 2924.800 2357.370 ;
        RECT 2898.065 2357.055 2898.395 2357.070 ;
        RECT 2917.600 2356.620 2924.800 2357.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 2622.320 455.790 2622.380 ;
        RECT 2900.830 2622.320 2901.150 2622.380 ;
        RECT 455.470 2622.180 2901.150 2622.320 ;
        RECT 455.470 2622.120 455.790 2622.180 ;
        RECT 2900.830 2622.120 2901.150 2622.180 ;
      LAYER via ;
        RECT 455.500 2622.120 455.760 2622.380 ;
        RECT 2900.860 2622.120 2901.120 2622.380 ;
      LAYER met2 ;
        RECT 455.500 2622.090 455.760 2622.410 ;
        RECT 2900.850 2622.235 2901.130 2622.605 ;
        RECT 2900.860 2622.090 2901.120 2622.235 ;
        RECT 455.560 1048.870 455.700 2622.090 ;
        RECT 455.560 1048.730 459.840 1048.870 ;
        RECT 459.700 999.330 459.840 1048.730 ;
        RECT 461.830 999.330 462.110 1000.000 ;
        RECT 459.700 999.190 462.110 999.330 ;
        RECT 461.830 996.000 462.110 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2622.280 2901.130 2622.560 ;
      LAYER met3 ;
        RECT 2900.825 2622.570 2901.155 2622.585 ;
        RECT 2917.600 2622.570 2924.800 2623.020 ;
        RECT 2900.825 2622.270 2924.800 2622.570 ;
        RECT 2900.825 2622.255 2901.155 2622.270 ;
        RECT 2917.600 2621.820 2924.800 2622.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 2884.460 483.390 2884.520 ;
        RECT 2898.070 2884.460 2898.390 2884.520 ;
        RECT 483.070 2884.320 2898.390 2884.460 ;
        RECT 483.070 2884.260 483.390 2884.320 ;
        RECT 2898.070 2884.260 2898.390 2884.320 ;
      LAYER via ;
        RECT 483.100 2884.260 483.360 2884.520 ;
        RECT 2898.100 2884.260 2898.360 2884.520 ;
      LAYER met2 ;
        RECT 2898.090 2888.115 2898.370 2888.485 ;
        RECT 2898.160 2884.550 2898.300 2888.115 ;
        RECT 483.100 2884.230 483.360 2884.550 ;
        RECT 2898.100 2884.230 2898.360 2884.550 ;
        RECT 483.160 999.330 483.300 2884.230 ;
        RECT 483.910 999.330 484.190 1000.000 ;
        RECT 483.160 999.190 484.190 999.330 ;
        RECT 483.910 996.000 484.190 999.190 ;
      LAYER via2 ;
        RECT 2898.090 2888.160 2898.370 2888.440 ;
      LAYER met3 ;
        RECT 2898.065 2888.450 2898.395 2888.465 ;
        RECT 2917.600 2888.450 2924.800 2888.900 ;
        RECT 2898.065 2888.150 2924.800 2888.450 ;
        RECT 2898.065 2888.135 2898.395 2888.150 ;
        RECT 2917.600 2887.700 2924.800 2888.150 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 3153.400 504.090 3153.460 ;
        RECT 2899.910 3153.400 2900.230 3153.460 ;
        RECT 503.770 3153.260 2900.230 3153.400 ;
        RECT 503.770 3153.200 504.090 3153.260 ;
        RECT 2899.910 3153.200 2900.230 3153.260 ;
      LAYER via ;
        RECT 503.800 3153.200 504.060 3153.460 ;
        RECT 2899.940 3153.200 2900.200 3153.460 ;
      LAYER met2 ;
        RECT 2899.930 3153.995 2900.210 3154.365 ;
        RECT 2900.000 3153.490 2900.140 3153.995 ;
        RECT 503.800 3153.170 504.060 3153.490 ;
        RECT 2899.940 3153.170 2900.200 3153.490 ;
        RECT 503.860 999.330 504.000 3153.170 ;
        RECT 505.990 999.330 506.270 1000.000 ;
        RECT 503.860 999.190 506.270 999.330 ;
        RECT 505.990 996.000 506.270 999.190 ;
      LAYER via2 ;
        RECT 2899.930 3154.040 2900.210 3154.320 ;
      LAYER met3 ;
        RECT 2899.905 3154.330 2900.235 3154.345 ;
        RECT 2917.600 3154.330 2924.800 3154.780 ;
        RECT 2899.905 3154.030 2924.800 3154.330 ;
        RECT 2899.905 3154.015 2900.235 3154.030 ;
        RECT 2917.600 3153.580 2924.800 3154.030 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 3415.880 524.790 3415.940 ;
        RECT 2900.830 3415.880 2901.150 3415.940 ;
        RECT 524.470 3415.740 2901.150 3415.880 ;
        RECT 524.470 3415.680 524.790 3415.740 ;
        RECT 2900.830 3415.680 2901.150 3415.740 ;
      LAYER via ;
        RECT 524.500 3415.680 524.760 3415.940 ;
        RECT 2900.860 3415.680 2901.120 3415.940 ;
      LAYER met2 ;
        RECT 2900.850 3419.195 2901.130 3419.565 ;
        RECT 2900.920 3415.970 2901.060 3419.195 ;
        RECT 524.500 3415.650 524.760 3415.970 ;
        RECT 2900.860 3415.650 2901.120 3415.970 ;
        RECT 524.560 1048.870 524.700 3415.650 ;
        RECT 524.560 1048.730 526.080 1048.870 ;
        RECT 525.940 999.330 526.080 1048.730 ;
        RECT 528.070 999.330 528.350 1000.000 ;
        RECT 525.940 999.190 528.350 999.330 ;
        RECT 528.070 996.000 528.350 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3419.240 2901.130 3419.520 ;
      LAYER met3 ;
        RECT 2900.825 3419.530 2901.155 3419.545 ;
        RECT 2917.600 3419.530 2924.800 3419.980 ;
        RECT 2900.825 3419.230 2924.800 3419.530 ;
        RECT 2900.825 3419.215 2901.155 3419.230 ;
        RECT 2917.600 3418.780 2924.800 3419.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.845 2717.520 3517.600 ;
        RECT 545.190 3501.475 545.470 3501.845 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
        RECT 545.260 1048.870 545.400 3501.475 ;
        RECT 545.260 1048.730 548.160 1048.870 ;
        RECT 548.020 999.330 548.160 1048.730 ;
        RECT 550.150 999.330 550.430 1000.000 ;
        RECT 548.020 999.190 550.430 999.330 ;
        RECT 550.150 996.000 550.430 999.190 ;
      LAYER via2 ;
        RECT 545.190 3501.520 545.470 3501.800 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 545.165 3501.810 545.495 3501.825 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 545.165 3501.510 2717.615 3501.810 ;
        RECT 545.165 3501.495 545.495 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.525 2392.760 3517.600 ;
        RECT 572.790 3502.155 573.070 3502.525 ;
        RECT 2392.550 3502.155 2392.830 3502.525 ;
        RECT 572.860 1048.870 573.000 3502.155 ;
        RECT 572.860 1048.730 573.460 1048.870 ;
        RECT 572.690 999.330 572.970 1000.000 ;
        RECT 573.320 999.330 573.460 1048.730 ;
        RECT 572.690 999.190 573.460 999.330 ;
        RECT 572.690 996.000 572.970 999.190 ;
      LAYER via2 ;
        RECT 572.790 3502.200 573.070 3502.480 ;
        RECT 2392.550 3502.200 2392.830 3502.480 ;
      LAYER met3 ;
        RECT 572.765 3502.490 573.095 3502.505 ;
        RECT 2392.525 3502.490 2392.855 3502.505 ;
        RECT 572.765 3502.190 2392.855 3502.490 ;
        RECT 572.765 3502.175 573.095 3502.190 ;
        RECT 2392.525 3502.175 2392.855 3502.190 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 3501.900 593.790 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 593.470 3501.760 2068.550 3501.900 ;
        RECT 593.470 3501.700 593.790 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 593.500 3501.700 593.760 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 593.500 3501.670 593.760 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 593.560 999.330 593.700 3501.670 ;
        RECT 594.770 999.330 595.050 1000.000 ;
        RECT 593.560 999.190 595.050 999.330 ;
        RECT 594.770 996.000 595.050 999.190 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 3502.580 614.490 3502.640 ;
        RECT 1743.930 3502.580 1744.250 3502.640 ;
        RECT 614.170 3502.440 1744.250 3502.580 ;
        RECT 614.170 3502.380 614.490 3502.440 ;
        RECT 1743.930 3502.380 1744.250 3502.440 ;
      LAYER via ;
        RECT 614.200 3502.380 614.460 3502.640 ;
        RECT 1743.960 3502.380 1744.220 3502.640 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.670 1744.160 3517.600 ;
        RECT 614.200 3502.350 614.460 3502.670 ;
        RECT 1743.960 3502.350 1744.220 3502.670 ;
        RECT 614.260 1048.870 614.400 3502.350 ;
        RECT 614.260 1048.730 615.320 1048.870 ;
        RECT 615.180 999.330 615.320 1048.730 ;
        RECT 616.850 999.330 617.130 1000.000 ;
        RECT 615.180 999.190 617.130 999.330 ;
        RECT 616.850 996.000 617.130 999.190 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.870 3503.260 635.190 3503.320 ;
        RECT 1419.170 3503.260 1419.490 3503.320 ;
        RECT 634.870 3503.120 1419.490 3503.260 ;
        RECT 634.870 3503.060 635.190 3503.120 ;
        RECT 1419.170 3503.060 1419.490 3503.120 ;
      LAYER via ;
        RECT 634.900 3503.060 635.160 3503.320 ;
        RECT 1419.200 3503.060 1419.460 3503.320 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3503.350 1419.400 3517.600 ;
        RECT 634.900 3503.030 635.160 3503.350 ;
        RECT 1419.200 3503.030 1419.460 3503.350 ;
        RECT 634.960 1048.870 635.100 3503.030 ;
        RECT 634.960 1048.730 637.400 1048.870 ;
        RECT 637.260 999.330 637.400 1048.730 ;
        RECT 638.930 999.330 639.210 1000.000 ;
        RECT 637.260 999.190 639.210 999.330 ;
        RECT 638.930 996.000 639.210 999.190 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.490 997.600 242.810 997.860 ;
        RECT 242.580 995.080 242.720 997.600 ;
        RECT 242.580 994.940 274.920 995.080 ;
        RECT 274.780 994.740 274.920 994.940 ;
        RECT 274.780 994.600 276.070 994.740 ;
        RECT 275.930 994.400 276.070 994.600 ;
        RECT 275.930 994.260 283.660 994.400 ;
        RECT 283.520 993.380 283.660 994.260 ;
        RECT 2904.510 994.060 2904.830 994.120 ;
        RECT 351.830 993.920 2904.830 994.060 ;
        RECT 351.830 993.720 351.970 993.920 ;
        RECT 2904.510 993.860 2904.830 993.920 ;
        RECT 331.130 993.580 338.170 993.720 ;
        RECT 283.520 993.240 308.040 993.380 ;
        RECT 307.900 993.040 308.040 993.240 ;
        RECT 331.130 993.040 331.270 993.580 ;
        RECT 338.030 993.380 338.170 993.580 ;
        RECT 344.930 993.580 351.970 993.720 ;
        RECT 344.930 993.380 345.070 993.580 ;
        RECT 338.030 993.240 345.070 993.380 ;
        RECT 307.900 992.900 331.270 993.040 ;
      LAYER via ;
        RECT 242.520 997.600 242.780 997.860 ;
        RECT 2904.540 993.860 2904.800 994.120 ;
      LAYER met2 ;
        RECT 240.570 997.970 240.850 1000.000 ;
        RECT 240.570 997.890 242.720 997.970 ;
        RECT 240.570 997.830 242.780 997.890 ;
        RECT 240.570 996.000 240.850 997.830 ;
        RECT 242.520 997.570 242.780 997.830 ;
        RECT 2904.540 993.830 2904.800 994.150 ;
        RECT 2904.600 298.365 2904.740 993.830 ;
        RECT 2904.530 297.995 2904.810 298.365 ;
      LAYER via2 ;
        RECT 2904.530 298.040 2904.810 298.320 ;
      LAYER met3 ;
        RECT 2904.505 298.330 2904.835 298.345 ;
        RECT 2917.600 298.330 2924.800 298.780 ;
        RECT 2904.505 298.030 2924.800 298.330 ;
        RECT 2904.505 298.015 2904.835 298.030 ;
        RECT 2917.600 297.580 2924.800 298.030 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 655.570 3504.960 655.890 3505.020 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 655.570 3504.820 1095.190 3504.960 ;
        RECT 655.570 3504.760 655.890 3504.820 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
      LAYER via ;
        RECT 655.600 3504.760 655.860 3505.020 ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 655.600 3504.730 655.860 3505.050 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 655.660 1048.870 655.800 3504.730 ;
        RECT 655.660 1048.730 659.480 1048.870 ;
        RECT 659.340 999.330 659.480 1048.730 ;
        RECT 661.010 999.330 661.290 1000.000 ;
        RECT 659.340 999.190 661.290 999.330 ;
        RECT 661.010 996.000 661.290 999.190 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 3499.860 683.950 3499.920 ;
        RECT 770.570 3499.860 770.890 3499.920 ;
        RECT 683.630 3499.720 770.890 3499.860 ;
        RECT 683.630 3499.660 683.950 3499.720 ;
        RECT 770.570 3499.660 770.890 3499.720 ;
      LAYER via ;
        RECT 683.660 3499.660 683.920 3499.920 ;
        RECT 770.600 3499.660 770.860 3499.920 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3499.950 770.800 3517.600 ;
        RECT 683.660 3499.630 683.920 3499.950 ;
        RECT 770.600 3499.630 770.860 3499.950 ;
        RECT 683.090 999.330 683.370 1000.000 ;
        RECT 683.720 999.330 683.860 3499.630 ;
        RECT 683.090 999.190 683.860 999.330 ;
        RECT 683.090 996.000 683.370 999.190 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3500.540 446.130 3500.600 ;
        RECT 703.870 3500.540 704.190 3500.600 ;
        RECT 445.810 3500.400 704.190 3500.540 ;
        RECT 445.810 3500.340 446.130 3500.400 ;
        RECT 703.870 3500.340 704.190 3500.400 ;
      LAYER via ;
        RECT 445.840 3500.340 446.100 3500.600 ;
        RECT 703.900 3500.340 704.160 3500.600 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3500.630 446.040 3517.600 ;
        RECT 445.840 3500.310 446.100 3500.630 ;
        RECT 703.900 3500.310 704.160 3500.630 ;
        RECT 703.960 999.330 704.100 3500.310 ;
        RECT 705.170 999.330 705.450 1000.000 ;
        RECT 703.960 999.190 705.450 999.330 ;
        RECT 705.170 996.000 705.450 999.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3504.280 121.830 3504.340 ;
        RECT 724.570 3504.280 724.890 3504.340 ;
        RECT 121.510 3504.140 724.890 3504.280 ;
        RECT 121.510 3504.080 121.830 3504.140 ;
        RECT 724.570 3504.080 724.890 3504.140 ;
      LAYER via ;
        RECT 121.540 3504.080 121.800 3504.340 ;
        RECT 724.600 3504.080 724.860 3504.340 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3504.370 121.740 3517.600 ;
        RECT 121.540 3504.050 121.800 3504.370 ;
        RECT 724.600 3504.050 724.860 3504.370 ;
        RECT 724.660 1048.870 724.800 3504.050 ;
        RECT 724.660 1048.730 725.720 1048.870 ;
        RECT 725.580 999.330 725.720 1048.730 ;
        RECT 727.250 999.330 727.530 1000.000 ;
        RECT 725.580 999.190 727.530 999.330 ;
        RECT 727.250 996.000 727.530 999.190 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 3354.000 17.410 3354.060 ;
        RECT 745.270 3354.000 745.590 3354.060 ;
        RECT 17.090 3353.860 745.590 3354.000 ;
        RECT 17.090 3353.800 17.410 3353.860 ;
        RECT 745.270 3353.800 745.590 3353.860 ;
      LAYER via ;
        RECT 17.120 3353.800 17.380 3354.060 ;
        RECT 745.300 3353.800 745.560 3354.060 ;
      LAYER met2 ;
        RECT 17.110 3355.955 17.390 3356.325 ;
        RECT 17.180 3354.090 17.320 3355.955 ;
        RECT 17.120 3353.770 17.380 3354.090 ;
        RECT 745.300 3353.770 745.560 3354.090 ;
        RECT 745.360 1048.870 745.500 3353.770 ;
        RECT 745.360 1048.730 747.800 1048.870 ;
        RECT 747.660 999.330 747.800 1048.730 ;
        RECT 749.790 999.330 750.070 1000.000 ;
        RECT 747.660 999.190 750.070 999.330 ;
        RECT 749.790 996.000 750.070 999.190 ;
      LAYER via2 ;
        RECT 17.110 3356.000 17.390 3356.280 ;
      LAYER met3 ;
        RECT -4.800 3356.290 2.400 3356.740 ;
        RECT 17.085 3356.290 17.415 3356.305 ;
        RECT -4.800 3355.990 17.415 3356.290 ;
        RECT -4.800 3355.540 2.400 3355.990 ;
        RECT 17.085 3355.975 17.415 3355.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 3091.520 16.030 3091.580 ;
        RECT 765.970 3091.520 766.290 3091.580 ;
        RECT 15.710 3091.380 766.290 3091.520 ;
        RECT 15.710 3091.320 16.030 3091.380 ;
        RECT 765.970 3091.320 766.290 3091.380 ;
      LAYER via ;
        RECT 15.740 3091.320 16.000 3091.580 ;
        RECT 766.000 3091.320 766.260 3091.580 ;
      LAYER met2 ;
        RECT 15.730 3095.515 16.010 3095.885 ;
        RECT 15.800 3091.610 15.940 3095.515 ;
        RECT 15.740 3091.290 16.000 3091.610 ;
        RECT 766.000 3091.290 766.260 3091.610 ;
        RECT 766.060 1048.870 766.200 3091.290 ;
        RECT 766.060 1048.730 769.880 1048.870 ;
        RECT 769.740 999.330 769.880 1048.730 ;
        RECT 771.870 999.330 772.150 1000.000 ;
        RECT 769.740 999.190 772.150 999.330 ;
        RECT 771.870 996.000 772.150 999.190 ;
      LAYER via2 ;
        RECT 15.730 3095.560 16.010 3095.840 ;
      LAYER met3 ;
        RECT -4.800 3095.850 2.400 3096.300 ;
        RECT 15.705 3095.850 16.035 3095.865 ;
        RECT -4.800 3095.550 16.035 3095.850 ;
        RECT -4.800 3095.100 2.400 3095.550 ;
        RECT 15.705 3095.535 16.035 3095.550 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2829.380 17.410 2829.440 ;
        RECT 793.570 2829.380 793.890 2829.440 ;
        RECT 17.090 2829.240 793.890 2829.380 ;
        RECT 17.090 2829.180 17.410 2829.240 ;
        RECT 793.570 2829.180 793.890 2829.240 ;
      LAYER via ;
        RECT 17.120 2829.180 17.380 2829.440 ;
        RECT 793.600 2829.180 793.860 2829.440 ;
      LAYER met2 ;
        RECT 17.110 2834.395 17.390 2834.765 ;
        RECT 17.180 2829.470 17.320 2834.395 ;
        RECT 17.120 2829.150 17.380 2829.470 ;
        RECT 793.600 2829.150 793.860 2829.470 ;
        RECT 793.660 999.330 793.800 2829.150 ;
        RECT 793.950 999.330 794.230 1000.000 ;
        RECT 793.660 999.190 794.230 999.330 ;
        RECT 793.950 996.000 794.230 999.190 ;
      LAYER via2 ;
        RECT 17.110 2834.440 17.390 2834.720 ;
      LAYER met3 ;
        RECT -4.800 2834.730 2.400 2835.180 ;
        RECT 17.085 2834.730 17.415 2834.745 ;
        RECT -4.800 2834.430 17.415 2834.730 ;
        RECT -4.800 2833.980 2.400 2834.430 ;
        RECT 17.085 2834.415 17.415 2834.430 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 2574.040 17.410 2574.100 ;
        RECT 814.270 2574.040 814.590 2574.100 ;
        RECT 17.090 2573.900 814.590 2574.040 ;
        RECT 17.090 2573.840 17.410 2573.900 ;
        RECT 814.270 2573.840 814.590 2573.900 ;
      LAYER via ;
        RECT 17.120 2573.840 17.380 2574.100 ;
        RECT 814.300 2573.840 814.560 2574.100 ;
      LAYER met2 ;
        RECT 17.110 2573.955 17.390 2574.325 ;
        RECT 17.120 2573.810 17.380 2573.955 ;
        RECT 814.300 2573.810 814.560 2574.130 ;
        RECT 814.360 999.330 814.500 2573.810 ;
        RECT 816.030 999.330 816.310 1000.000 ;
        RECT 814.360 999.190 816.310 999.330 ;
        RECT 816.030 996.000 816.310 999.190 ;
      LAYER via2 ;
        RECT 17.110 2574.000 17.390 2574.280 ;
      LAYER met3 ;
        RECT -4.800 2574.290 2.400 2574.740 ;
        RECT 17.085 2574.290 17.415 2574.305 ;
        RECT -4.800 2573.990 17.415 2574.290 ;
        RECT -4.800 2573.540 2.400 2573.990 ;
        RECT 17.085 2573.975 17.415 2573.990 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2311.900 16.490 2311.960 ;
        RECT 834.970 2311.900 835.290 2311.960 ;
        RECT 16.170 2311.760 835.290 2311.900 ;
        RECT 16.170 2311.700 16.490 2311.760 ;
        RECT 834.970 2311.700 835.290 2311.760 ;
      LAYER via ;
        RECT 16.200 2311.700 16.460 2311.960 ;
        RECT 835.000 2311.700 835.260 2311.960 ;
      LAYER met2 ;
        RECT 16.190 2312.835 16.470 2313.205 ;
        RECT 16.260 2311.990 16.400 2312.835 ;
        RECT 16.200 2311.670 16.460 2311.990 ;
        RECT 835.000 2311.670 835.260 2311.990 ;
        RECT 835.060 1048.870 835.200 2311.670 ;
        RECT 835.060 1048.730 836.120 1048.870 ;
        RECT 835.980 999.330 836.120 1048.730 ;
        RECT 838.110 999.330 838.390 1000.000 ;
        RECT 835.980 999.190 838.390 999.330 ;
        RECT 838.110 996.000 838.390 999.190 ;
      LAYER via2 ;
        RECT 16.190 2312.880 16.470 2313.160 ;
      LAYER met3 ;
        RECT -4.800 2313.170 2.400 2313.620 ;
        RECT 16.165 2313.170 16.495 2313.185 ;
        RECT -4.800 2312.870 16.495 2313.170 ;
        RECT -4.800 2312.420 2.400 2312.870 ;
        RECT 16.165 2312.855 16.495 2312.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2049.420 16.030 2049.480 ;
        RECT 855.670 2049.420 855.990 2049.480 ;
        RECT 15.710 2049.280 855.990 2049.420 ;
        RECT 15.710 2049.220 16.030 2049.280 ;
        RECT 855.670 2049.220 855.990 2049.280 ;
      LAYER via ;
        RECT 15.740 2049.220 16.000 2049.480 ;
        RECT 855.700 2049.220 855.960 2049.480 ;
      LAYER met2 ;
        RECT 15.730 2052.395 16.010 2052.765 ;
        RECT 15.800 2049.510 15.940 2052.395 ;
        RECT 15.740 2049.190 16.000 2049.510 ;
        RECT 855.700 2049.190 855.960 2049.510 ;
        RECT 855.760 1048.870 855.900 2049.190 ;
        RECT 855.760 1048.730 858.200 1048.870 ;
        RECT 858.060 999.330 858.200 1048.730 ;
        RECT 860.190 999.330 860.470 1000.000 ;
        RECT 858.060 999.190 860.470 999.330 ;
        RECT 860.190 996.000 860.470 999.190 ;
      LAYER via2 ;
        RECT 15.730 2052.440 16.010 2052.720 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 15.705 2052.730 16.035 2052.745 ;
        RECT -4.800 2052.430 16.035 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 15.705 2052.415 16.035 2052.430 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1100.390 503.440 1100.710 503.500 ;
        RECT 2899.450 503.440 2899.770 503.500 ;
        RECT 1100.390 503.300 2899.770 503.440 ;
        RECT 1100.390 503.240 1100.710 503.300 ;
        RECT 2899.450 503.240 2899.770 503.300 ;
      LAYER via ;
        RECT 1100.420 503.240 1100.680 503.500 ;
        RECT 2899.480 503.240 2899.740 503.500 ;
      LAYER met2 ;
        RECT 264.590 1011.315 264.870 1011.685 ;
        RECT 1100.410 1011.315 1100.690 1011.685 ;
        RECT 262.650 999.330 262.930 1000.000 ;
        RECT 264.660 999.330 264.800 1011.315 ;
        RECT 262.650 999.190 264.800 999.330 ;
        RECT 262.650 996.000 262.930 999.190 ;
        RECT 1100.480 503.530 1100.620 1011.315 ;
        RECT 1100.420 503.210 1100.680 503.530 ;
        RECT 2899.480 503.210 2899.740 503.530 ;
        RECT 2899.540 497.605 2899.680 503.210 ;
        RECT 2899.470 497.235 2899.750 497.605 ;
      LAYER via2 ;
        RECT 264.590 1011.360 264.870 1011.640 ;
        RECT 1100.410 1011.360 1100.690 1011.640 ;
        RECT 2899.470 497.280 2899.750 497.560 ;
      LAYER met3 ;
        RECT 264.565 1011.650 264.895 1011.665 ;
        RECT 1100.385 1011.650 1100.715 1011.665 ;
        RECT 264.565 1011.350 1100.715 1011.650 ;
        RECT 264.565 1011.335 264.895 1011.350 ;
        RECT 1100.385 1011.335 1100.715 1011.350 ;
        RECT 2899.445 497.570 2899.775 497.585 ;
        RECT 2917.600 497.570 2924.800 498.020 ;
        RECT 2899.445 497.270 2924.800 497.570 ;
        RECT 2899.445 497.255 2899.775 497.270 ;
        RECT 2917.600 496.820 2924.800 497.270 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1787.280 16.030 1787.340 ;
        RECT 876.370 1787.280 876.690 1787.340 ;
        RECT 15.710 1787.140 876.690 1787.280 ;
        RECT 15.710 1787.080 16.030 1787.140 ;
        RECT 876.370 1787.080 876.690 1787.140 ;
      LAYER via ;
        RECT 15.740 1787.080 16.000 1787.340 ;
        RECT 876.400 1787.080 876.660 1787.340 ;
      LAYER met2 ;
        RECT 15.730 1791.955 16.010 1792.325 ;
        RECT 15.800 1787.370 15.940 1791.955 ;
        RECT 15.740 1787.050 16.000 1787.370 ;
        RECT 876.400 1787.050 876.660 1787.370 ;
        RECT 876.460 1048.870 876.600 1787.050 ;
        RECT 876.460 1048.730 880.280 1048.870 ;
        RECT 880.140 999.330 880.280 1048.730 ;
        RECT 882.270 999.330 882.550 1000.000 ;
        RECT 880.140 999.190 882.550 999.330 ;
        RECT 882.270 996.000 882.550 999.190 ;
      LAYER via2 ;
        RECT 15.730 1792.000 16.010 1792.280 ;
      LAYER met3 ;
        RECT -4.800 1792.290 2.400 1792.740 ;
        RECT 15.705 1792.290 16.035 1792.305 ;
        RECT -4.800 1791.990 16.035 1792.290 ;
        RECT -4.800 1791.540 2.400 1791.990 ;
        RECT 15.705 1791.975 16.035 1791.990 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1525.140 17.870 1525.200 ;
        RECT 903.970 1525.140 904.290 1525.200 ;
        RECT 17.550 1525.000 904.290 1525.140 ;
        RECT 17.550 1524.940 17.870 1525.000 ;
        RECT 903.970 1524.940 904.290 1525.000 ;
      LAYER via ;
        RECT 17.580 1524.940 17.840 1525.200 ;
        RECT 904.000 1524.940 904.260 1525.200 ;
      LAYER met2 ;
        RECT 17.570 1530.835 17.850 1531.205 ;
        RECT 17.640 1525.230 17.780 1530.835 ;
        RECT 17.580 1524.910 17.840 1525.230 ;
        RECT 904.000 1524.910 904.260 1525.230 ;
        RECT 904.060 999.330 904.200 1524.910 ;
        RECT 904.350 999.330 904.630 1000.000 ;
        RECT 904.060 999.190 904.630 999.330 ;
        RECT 904.350 996.000 904.630 999.190 ;
      LAYER via2 ;
        RECT 17.570 1530.880 17.850 1531.160 ;
      LAYER met3 ;
        RECT -4.800 1531.170 2.400 1531.620 ;
        RECT 17.545 1531.170 17.875 1531.185 ;
        RECT -4.800 1530.870 17.875 1531.170 ;
        RECT -4.800 1530.420 2.400 1530.870 ;
        RECT 17.545 1530.855 17.875 1530.870 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1269.800 17.870 1269.860 ;
        RECT 924.670 1269.800 924.990 1269.860 ;
        RECT 17.550 1269.660 924.990 1269.800 ;
        RECT 17.550 1269.600 17.870 1269.660 ;
        RECT 924.670 1269.600 924.990 1269.660 ;
      LAYER via ;
        RECT 17.580 1269.600 17.840 1269.860 ;
        RECT 924.700 1269.600 924.960 1269.860 ;
      LAYER met2 ;
        RECT 17.570 1270.395 17.850 1270.765 ;
        RECT 17.640 1269.890 17.780 1270.395 ;
        RECT 17.580 1269.570 17.840 1269.890 ;
        RECT 924.700 1269.570 924.960 1269.890 ;
        RECT 924.760 1048.870 924.900 1269.570 ;
        RECT 924.760 1048.730 925.360 1048.870 ;
        RECT 925.220 999.330 925.360 1048.730 ;
        RECT 926.890 999.330 927.170 1000.000 ;
        RECT 925.220 999.190 927.170 999.330 ;
        RECT 926.890 996.000 927.170 999.190 ;
      LAYER via2 ;
        RECT 17.570 1270.440 17.850 1270.720 ;
      LAYER met3 ;
        RECT -4.800 1270.730 2.400 1271.180 ;
        RECT 17.545 1270.730 17.875 1270.745 ;
        RECT -4.800 1270.430 17.875 1270.730 ;
        RECT -4.800 1269.980 2.400 1270.430 ;
        RECT 17.545 1270.415 17.875 1270.430 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1010.040 17.870 1010.100 ;
        RECT 947.670 1010.040 947.990 1010.100 ;
        RECT 17.550 1009.900 947.990 1010.040 ;
        RECT 17.550 1009.840 17.870 1009.900 ;
        RECT 947.670 1009.840 947.990 1009.900 ;
      LAYER via ;
        RECT 17.580 1009.840 17.840 1010.100 ;
        RECT 947.700 1009.840 947.960 1010.100 ;
      LAYER met2 ;
        RECT 17.580 1009.810 17.840 1010.130 ;
        RECT 947.700 1009.810 947.960 1010.130 ;
        RECT 17.640 1009.645 17.780 1009.810 ;
        RECT 17.570 1009.275 17.850 1009.645 ;
        RECT 947.760 999.330 947.900 1009.810 ;
        RECT 948.970 999.330 949.250 1000.000 ;
        RECT 947.760 999.190 949.250 999.330 ;
        RECT 948.970 996.000 949.250 999.190 ;
      LAYER via2 ;
        RECT 17.570 1009.320 17.850 1009.600 ;
      LAYER met3 ;
        RECT -4.800 1009.610 2.400 1010.060 ;
        RECT 17.545 1009.610 17.875 1009.625 ;
        RECT -4.800 1009.310 17.875 1009.610 ;
        RECT -4.800 1008.860 2.400 1009.310 ;
        RECT 17.545 1009.295 17.875 1009.310 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1009.020 16.490 1009.080 ;
        RECT 969.750 1009.020 970.070 1009.080 ;
        RECT 16.170 1008.880 970.070 1009.020 ;
        RECT 16.170 1008.820 16.490 1008.880 ;
        RECT 969.750 1008.820 970.070 1008.880 ;
      LAYER via ;
        RECT 16.200 1008.820 16.460 1009.080 ;
        RECT 969.780 1008.820 970.040 1009.080 ;
      LAYER met2 ;
        RECT 16.200 1008.790 16.460 1009.110 ;
        RECT 969.780 1008.790 970.040 1009.110 ;
        RECT 16.260 749.205 16.400 1008.790 ;
        RECT 969.840 999.330 969.980 1008.790 ;
        RECT 971.050 999.330 971.330 1000.000 ;
        RECT 969.840 999.190 971.330 999.330 ;
        RECT 971.050 996.000 971.330 999.190 ;
        RECT 16.190 748.835 16.470 749.205 ;
      LAYER via2 ;
        RECT 16.190 748.880 16.470 749.160 ;
      LAYER met3 ;
        RECT -4.800 749.170 2.400 749.620 ;
        RECT 16.165 749.170 16.495 749.185 ;
        RECT -4.800 748.870 16.495 749.170 ;
        RECT -4.800 748.420 2.400 748.870 ;
        RECT 16.165 748.855 16.495 748.870 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.390 1008.340 19.710 1008.400 ;
        RECT 991.830 1008.340 992.150 1008.400 ;
        RECT 19.390 1008.200 992.150 1008.340 ;
        RECT 19.390 1008.140 19.710 1008.200 ;
        RECT 991.830 1008.140 992.150 1008.200 ;
      LAYER via ;
        RECT 19.420 1008.140 19.680 1008.400 ;
        RECT 991.860 1008.140 992.120 1008.400 ;
      LAYER met2 ;
        RECT 19.420 1008.110 19.680 1008.430 ;
        RECT 991.860 1008.110 992.120 1008.430 ;
        RECT 19.480 488.085 19.620 1008.110 ;
        RECT 991.920 999.330 992.060 1008.110 ;
        RECT 993.130 999.330 993.410 1000.000 ;
        RECT 991.920 999.190 993.410 999.330 ;
        RECT 993.130 996.000 993.410 999.190 ;
        RECT 19.410 487.715 19.690 488.085 ;
      LAYER via2 ;
        RECT 19.410 487.760 19.690 488.040 ;
      LAYER met3 ;
        RECT -4.800 488.050 2.400 488.500 ;
        RECT 19.385 488.050 19.715 488.065 ;
        RECT -4.800 487.750 19.715 488.050 ;
        RECT -4.800 487.300 2.400 487.750 ;
        RECT 19.385 487.735 19.715 487.750 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 293.090 997.260 293.410 997.520 ;
        RECT 972.510 997.260 972.830 997.520 ;
        RECT 293.180 996.780 293.320 997.260 ;
        RECT 293.180 996.640 331.270 996.780 ;
        RECT 196.490 995.420 196.810 995.480 ;
        RECT 201.090 995.420 201.410 995.480 ;
        RECT 196.490 995.280 201.410 995.420 ;
        RECT 196.490 995.220 196.810 995.280 ;
        RECT 201.090 995.220 201.410 995.280 ;
        RECT 331.130 995.080 331.270 996.640 ;
        RECT 972.600 995.760 972.740 997.260 ;
        RECT 903.830 995.620 931.570 995.760 ;
        RECT 903.830 995.080 903.970 995.620 ;
        RECT 931.430 995.420 931.570 995.620 ;
        RECT 971.680 995.620 972.740 995.760 ;
        RECT 931.430 995.280 966.070 995.420 ;
        RECT 331.130 994.940 903.970 995.080 ;
        RECT 965.930 995.080 966.070 995.280 ;
        RECT 971.680 995.080 971.820 995.620 ;
        RECT 965.930 994.940 971.820 995.080 ;
        RECT 17.090 296.720 17.410 296.780 ;
        RECT 196.490 296.720 196.810 296.780 ;
        RECT 17.090 296.580 196.810 296.720 ;
        RECT 17.090 296.520 17.410 296.580 ;
        RECT 196.490 296.520 196.810 296.580 ;
      LAYER via ;
        RECT 293.120 997.260 293.380 997.520 ;
        RECT 972.540 997.260 972.800 997.520 ;
        RECT 196.520 995.220 196.780 995.480 ;
        RECT 201.120 995.220 201.380 995.480 ;
        RECT 17.120 296.520 17.380 296.780 ;
        RECT 196.520 296.520 196.780 296.780 ;
      LAYER met2 ;
        RECT 1015.210 997.970 1015.490 1000.000 ;
        RECT 1014.000 997.830 1015.490 997.970 ;
        RECT 293.120 997.405 293.380 997.550 ;
        RECT 972.540 997.405 972.800 997.550 ;
        RECT 1014.000 997.405 1014.140 997.830 ;
        RECT 201.110 997.035 201.390 997.405 ;
        RECT 293.110 997.035 293.390 997.405 ;
        RECT 972.530 997.035 972.810 997.405 ;
        RECT 1013.930 997.035 1014.210 997.405 ;
        RECT 201.180 995.510 201.320 997.035 ;
        RECT 1015.210 996.000 1015.490 997.830 ;
        RECT 196.520 995.190 196.780 995.510 ;
        RECT 201.120 995.190 201.380 995.510 ;
        RECT 196.580 296.810 196.720 995.190 ;
        RECT 17.120 296.490 17.380 296.810 ;
        RECT 196.520 296.490 196.780 296.810 ;
        RECT 17.180 292.925 17.320 296.490 ;
        RECT 17.110 292.555 17.390 292.925 ;
      LAYER via2 ;
        RECT 201.110 997.080 201.390 997.360 ;
        RECT 293.110 997.080 293.390 997.360 ;
        RECT 972.530 997.080 972.810 997.360 ;
        RECT 1013.930 997.080 1014.210 997.360 ;
        RECT 17.110 292.600 17.390 292.880 ;
      LAYER met3 ;
        RECT 201.085 997.370 201.415 997.385 ;
        RECT 293.085 997.370 293.415 997.385 ;
        RECT 201.085 997.070 293.415 997.370 ;
        RECT 201.085 997.055 201.415 997.070 ;
        RECT 293.085 997.055 293.415 997.070 ;
        RECT 972.505 997.370 972.835 997.385 ;
        RECT 1013.905 997.370 1014.235 997.385 ;
        RECT 972.505 997.070 1014.235 997.370 ;
        RECT 972.505 997.055 972.835 997.070 ;
        RECT 1013.905 997.055 1014.235 997.070 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 17.085 292.890 17.415 292.905 ;
        RECT -4.800 292.590 17.415 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 17.085 292.575 17.415 292.590 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 997.290 1036.290 997.405 ;
        RECT 1037.290 997.290 1037.570 1000.000 ;
        RECT 1036.010 997.150 1037.570 997.290 ;
        RECT 1036.010 997.035 1036.290 997.150 ;
        RECT 1037.290 996.000 1037.570 997.150 ;
      LAYER via2 ;
        RECT 1036.010 997.080 1036.290 997.360 ;
      LAYER met3 ;
        RECT 1018.710 997.370 1019.090 997.380 ;
        RECT 1035.985 997.370 1036.315 997.385 ;
        RECT 1018.710 997.070 1036.315 997.370 ;
        RECT 1018.710 997.060 1019.090 997.070 ;
        RECT 1035.985 997.055 1036.315 997.070 ;
        RECT 15.910 993.970 16.290 993.980 ;
        RECT 1018.710 993.970 1019.090 993.980 ;
        RECT 15.910 993.670 1019.090 993.970 ;
        RECT 15.910 993.660 16.290 993.670 ;
        RECT 1018.710 993.660 1019.090 993.670 ;
        RECT -4.800 97.050 2.400 97.500 ;
        RECT 15.910 97.050 16.290 97.060 ;
        RECT -4.800 96.750 16.290 97.050 ;
        RECT -4.800 96.300 2.400 96.750 ;
        RECT 15.910 96.740 16.290 96.750 ;
      LAYER via3 ;
        RECT 1018.740 997.060 1019.060 997.380 ;
        RECT 15.940 993.660 16.260 993.980 ;
        RECT 1018.740 993.660 1019.060 993.980 ;
        RECT 15.940 96.740 16.260 97.060 ;
      LAYER met4 ;
        RECT 1018.735 997.055 1019.065 997.385 ;
        RECT 1018.750 993.985 1019.050 997.055 ;
        RECT 15.935 993.655 16.265 993.985 ;
        RECT 1018.735 993.655 1019.065 993.985 ;
        RECT 15.950 97.065 16.250 993.655 ;
        RECT 15.935 96.735 16.265 97.065 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.650 1011.400 286.970 1011.460 ;
        RECT 1100.850 1011.400 1101.170 1011.460 ;
        RECT 286.650 1011.260 1101.170 1011.400 ;
        RECT 286.650 1011.200 286.970 1011.260 ;
        RECT 1100.850 1011.200 1101.170 1011.260 ;
        RECT 1100.850 696.900 1101.170 696.960 ;
        RECT 2899.450 696.900 2899.770 696.960 ;
        RECT 1100.850 696.760 2899.770 696.900 ;
        RECT 1100.850 696.700 1101.170 696.760 ;
        RECT 2899.450 696.700 2899.770 696.760 ;
      LAYER via ;
        RECT 286.680 1011.200 286.940 1011.460 ;
        RECT 1100.880 1011.200 1101.140 1011.460 ;
        RECT 1100.880 696.700 1101.140 696.960 ;
        RECT 2899.480 696.700 2899.740 696.960 ;
      LAYER met2 ;
        RECT 286.680 1011.170 286.940 1011.490 ;
        RECT 1100.880 1011.170 1101.140 1011.490 ;
        RECT 284.730 999.330 285.010 1000.000 ;
        RECT 286.740 999.330 286.880 1011.170 ;
        RECT 284.730 999.190 286.880 999.330 ;
        RECT 284.730 996.000 285.010 999.190 ;
        RECT 1100.940 696.990 1101.080 1011.170 ;
        RECT 1100.880 696.670 1101.140 696.990 ;
        RECT 2899.480 696.845 2899.740 696.990 ;
        RECT 2899.470 696.475 2899.750 696.845 ;
      LAYER via2 ;
        RECT 2899.470 696.520 2899.750 696.800 ;
      LAYER met3 ;
        RECT 2899.445 696.810 2899.775 696.825 ;
        RECT 2917.600 696.810 2924.800 697.260 ;
        RECT 2899.445 696.510 2924.800 696.810 ;
        RECT 2899.445 696.495 2899.775 696.510 ;
        RECT 2917.600 696.060 2924.800 696.510 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 308.730 1012.420 309.050 1012.480 ;
        RECT 1102.690 1012.420 1103.010 1012.480 ;
        RECT 308.730 1012.280 1103.010 1012.420 ;
        RECT 308.730 1012.220 309.050 1012.280 ;
        RECT 1102.690 1012.220 1103.010 1012.280 ;
        RECT 1102.690 896.820 1103.010 896.880 ;
        RECT 2899.450 896.820 2899.770 896.880 ;
        RECT 1102.690 896.680 2899.770 896.820 ;
        RECT 1102.690 896.620 1103.010 896.680 ;
        RECT 2899.450 896.620 2899.770 896.680 ;
      LAYER via ;
        RECT 308.760 1012.220 309.020 1012.480 ;
        RECT 1102.720 1012.220 1102.980 1012.480 ;
        RECT 1102.720 896.620 1102.980 896.880 ;
        RECT 2899.480 896.620 2899.740 896.880 ;
      LAYER met2 ;
        RECT 308.760 1012.190 309.020 1012.510 ;
        RECT 1102.720 1012.190 1102.980 1012.510 ;
        RECT 306.810 999.330 307.090 1000.000 ;
        RECT 308.820 999.330 308.960 1012.190 ;
        RECT 306.810 999.190 308.960 999.330 ;
        RECT 306.810 996.000 307.090 999.190 ;
        RECT 1102.780 896.910 1102.920 1012.190 ;
        RECT 1102.720 896.590 1102.980 896.910 ;
        RECT 2899.480 896.590 2899.740 896.910 ;
        RECT 2899.540 896.085 2899.680 896.590 ;
        RECT 2899.470 895.715 2899.750 896.085 ;
      LAYER via2 ;
        RECT 2899.470 895.760 2899.750 896.040 ;
      LAYER met3 ;
        RECT 2899.445 896.050 2899.775 896.065 ;
        RECT 2917.600 896.050 2924.800 896.500 ;
        RECT 2899.445 895.750 2924.800 896.050 ;
        RECT 2899.445 895.735 2899.775 895.750 ;
        RECT 2917.600 895.300 2924.800 895.750 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 1090.280 324.690 1090.340 ;
        RECT 2900.830 1090.280 2901.150 1090.340 ;
        RECT 324.370 1090.140 2901.150 1090.280 ;
        RECT 324.370 1090.080 324.690 1090.140 ;
        RECT 2900.830 1090.080 2901.150 1090.140 ;
      LAYER via ;
        RECT 324.400 1090.080 324.660 1090.340 ;
        RECT 2900.860 1090.080 2901.120 1090.340 ;
      LAYER met2 ;
        RECT 2900.850 1094.955 2901.130 1095.325 ;
        RECT 2900.920 1090.370 2901.060 1094.955 ;
        RECT 324.400 1090.050 324.660 1090.370 ;
        RECT 2900.860 1090.050 2901.120 1090.370 ;
        RECT 324.460 1048.870 324.600 1090.050 ;
        RECT 324.460 1048.730 327.360 1048.870 ;
        RECT 327.220 999.330 327.360 1048.730 ;
        RECT 328.890 999.330 329.170 1000.000 ;
        RECT 327.220 999.190 329.170 999.330 ;
        RECT 328.890 996.000 329.170 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1095.000 2901.130 1095.280 ;
      LAYER met3 ;
        RECT 2900.825 1095.290 2901.155 1095.305 ;
        RECT 2917.600 1095.290 2924.800 1095.740 ;
        RECT 2900.825 1094.990 2924.800 1095.290 ;
        RECT 2900.825 1094.975 2901.155 1094.990 ;
        RECT 2917.600 1094.540 2924.800 1094.990 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 1290.540 345.390 1290.600 ;
        RECT 2898.070 1290.540 2898.390 1290.600 ;
        RECT 345.070 1290.400 2898.390 1290.540 ;
        RECT 345.070 1290.340 345.390 1290.400 ;
        RECT 2898.070 1290.340 2898.390 1290.400 ;
      LAYER via ;
        RECT 345.100 1290.340 345.360 1290.600 ;
        RECT 2898.100 1290.340 2898.360 1290.600 ;
      LAYER met2 ;
        RECT 2898.090 1294.195 2898.370 1294.565 ;
        RECT 2898.160 1290.630 2898.300 1294.195 ;
        RECT 345.100 1290.310 345.360 1290.630 ;
        RECT 2898.100 1290.310 2898.360 1290.630 ;
        RECT 345.160 1048.870 345.300 1290.310 ;
        RECT 345.160 1048.730 349.440 1048.870 ;
        RECT 349.300 999.330 349.440 1048.730 ;
        RECT 350.970 999.330 351.250 1000.000 ;
        RECT 349.300 999.190 351.250 999.330 ;
        RECT 350.970 996.000 351.250 999.190 ;
      LAYER via2 ;
        RECT 2898.090 1294.240 2898.370 1294.520 ;
      LAYER met3 ;
        RECT 2898.065 1294.530 2898.395 1294.545 ;
        RECT 2917.600 1294.530 2924.800 1294.980 ;
        RECT 2898.065 1294.230 2924.800 1294.530 ;
        RECT 2898.065 1294.215 2898.395 1294.230 ;
        RECT 2917.600 1293.780 2924.800 1294.230 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 1559.480 372.990 1559.540 ;
        RECT 2900.830 1559.480 2901.150 1559.540 ;
        RECT 372.670 1559.340 2901.150 1559.480 ;
        RECT 372.670 1559.280 372.990 1559.340 ;
        RECT 2900.830 1559.280 2901.150 1559.340 ;
      LAYER via ;
        RECT 372.700 1559.280 372.960 1559.540 ;
        RECT 2900.860 1559.280 2901.120 1559.540 ;
      LAYER met2 ;
        RECT 2900.850 1560.075 2901.130 1560.445 ;
        RECT 2900.920 1559.570 2901.060 1560.075 ;
        RECT 372.700 1559.250 372.960 1559.570 ;
        RECT 2900.860 1559.250 2901.120 1559.570 ;
        RECT 372.760 999.330 372.900 1559.250 ;
        RECT 373.050 999.330 373.330 1000.000 ;
        RECT 372.760 999.190 373.330 999.330 ;
        RECT 373.050 996.000 373.330 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1560.120 2901.130 1560.400 ;
      LAYER met3 ;
        RECT 2900.825 1560.410 2901.155 1560.425 ;
        RECT 2917.600 1560.410 2924.800 1560.860 ;
        RECT 2900.825 1560.110 2924.800 1560.410 ;
        RECT 2900.825 1560.095 2901.155 1560.110 ;
        RECT 2917.600 1559.660 2924.800 1560.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.370 1821.960 393.690 1822.020 ;
        RECT 2900.830 1821.960 2901.150 1822.020 ;
        RECT 393.370 1821.820 2901.150 1821.960 ;
        RECT 393.370 1821.760 393.690 1821.820 ;
        RECT 2900.830 1821.760 2901.150 1821.820 ;
      LAYER via ;
        RECT 393.400 1821.760 393.660 1822.020 ;
        RECT 2900.860 1821.760 2901.120 1822.020 ;
      LAYER met2 ;
        RECT 2900.850 1825.275 2901.130 1825.645 ;
        RECT 2900.920 1822.050 2901.060 1825.275 ;
        RECT 393.400 1821.730 393.660 1822.050 ;
        RECT 2900.860 1821.730 2901.120 1822.050 ;
        RECT 393.460 999.330 393.600 1821.730 ;
        RECT 395.590 999.330 395.870 1000.000 ;
        RECT 393.460 999.190 395.870 999.330 ;
        RECT 395.590 996.000 395.870 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1825.320 2901.130 1825.600 ;
      LAYER met3 ;
        RECT 2900.825 1825.610 2901.155 1825.625 ;
        RECT 2917.600 1825.610 2924.800 1826.060 ;
        RECT 2900.825 1825.310 2924.800 1825.610 ;
        RECT 2900.825 1825.295 2901.155 1825.310 ;
        RECT 2917.600 1824.860 2924.800 1825.310 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 2090.900 414.390 2090.960 ;
        RECT 2900.830 2090.900 2901.150 2090.960 ;
        RECT 414.070 2090.760 2901.150 2090.900 ;
        RECT 414.070 2090.700 414.390 2090.760 ;
        RECT 2900.830 2090.700 2901.150 2090.760 ;
      LAYER via ;
        RECT 414.100 2090.700 414.360 2090.960 ;
        RECT 2900.860 2090.700 2901.120 2090.960 ;
      LAYER met2 ;
        RECT 2900.850 2091.155 2901.130 2091.525 ;
        RECT 2900.920 2090.990 2901.060 2091.155 ;
        RECT 414.100 2090.670 414.360 2090.990 ;
        RECT 2900.860 2090.670 2901.120 2090.990 ;
        RECT 414.160 1048.870 414.300 2090.670 ;
        RECT 414.160 1048.730 415.680 1048.870 ;
        RECT 415.540 999.330 415.680 1048.730 ;
        RECT 417.670 999.330 417.950 1000.000 ;
        RECT 415.540 999.190 417.950 999.330 ;
        RECT 417.670 996.000 417.950 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2091.200 2901.130 2091.480 ;
      LAYER met3 ;
        RECT 2900.825 2091.490 2901.155 2091.505 ;
        RECT 2917.600 2091.490 2924.800 2091.940 ;
        RECT 2900.825 2091.190 2924.800 2091.490 ;
        RECT 2900.825 2091.175 2901.155 2091.190 ;
        RECT 2917.600 2090.740 2924.800 2091.190 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.470 32.200 386.790 32.260 ;
        RECT 576.910 32.200 577.230 32.260 ;
        RECT 386.470 32.060 577.230 32.200 ;
        RECT 386.470 32.000 386.790 32.060 ;
        RECT 576.910 32.000 577.230 32.060 ;
        RECT 576.910 15.200 577.230 15.260 ;
        RECT 629.350 15.200 629.670 15.260 ;
        RECT 576.910 15.060 629.670 15.200 ;
        RECT 576.910 15.000 577.230 15.060 ;
        RECT 629.350 15.000 629.670 15.060 ;
      LAYER via ;
        RECT 386.500 32.000 386.760 32.260 ;
        RECT 576.940 32.000 577.200 32.260 ;
        RECT 576.940 15.000 577.200 15.260 ;
        RECT 629.380 15.000 629.640 15.260 ;
      LAYER met2 ;
        RECT 389.610 400.250 389.890 404.000 ;
        RECT 388.400 400.110 389.890 400.250 ;
        RECT 388.400 387.330 388.540 400.110 ;
        RECT 389.610 400.000 389.890 400.110 ;
        RECT 386.560 387.190 388.540 387.330 ;
        RECT 386.560 32.290 386.700 387.190 ;
        RECT 386.500 31.970 386.760 32.290 ;
        RECT 576.940 31.970 577.200 32.290 ;
        RECT 577.000 15.290 577.140 31.970 ;
        RECT 576.940 14.970 577.200 15.290 ;
        RECT 629.380 14.970 629.640 15.290 ;
        RECT 629.440 2.400 629.580 14.970 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 926.050 109.040 926.370 109.100 ;
        RECT 2401.270 109.040 2401.590 109.100 ;
        RECT 926.050 108.900 2401.590 109.040 ;
        RECT 926.050 108.840 926.370 108.900 ;
        RECT 2401.270 108.840 2401.590 108.900 ;
      LAYER via ;
        RECT 926.080 108.840 926.340 109.100 ;
        RECT 2401.300 108.840 2401.560 109.100 ;
      LAYER met2 ;
        RECT 925.510 400.250 925.790 404.000 ;
        RECT 925.220 400.110 925.790 400.250 ;
        RECT 925.220 398.890 925.360 400.110 ;
        RECT 925.510 400.000 925.790 400.110 ;
        RECT 925.220 398.750 925.820 398.890 ;
        RECT 925.680 376.450 925.820 398.750 ;
        RECT 925.680 376.310 926.280 376.450 ;
        RECT 926.140 109.130 926.280 376.310 ;
        RECT 926.080 108.810 926.340 109.130 ;
        RECT 2401.300 108.810 2401.560 109.130 ;
        RECT 2401.360 82.870 2401.500 108.810 ;
        RECT 2401.360 82.730 2402.880 82.870 ;
        RECT 2402.740 2.400 2402.880 82.730 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.590 375.940 925.910 376.000 ;
        RECT 929.730 375.940 930.050 376.000 ;
        RECT 925.590 375.800 930.050 375.940 ;
        RECT 925.590 375.740 925.910 375.800 ;
        RECT 929.730 375.740 930.050 375.800 ;
        RECT 925.590 108.700 925.910 108.760 ;
        RECT 2415.070 108.700 2415.390 108.760 ;
        RECT 925.590 108.560 2415.390 108.700 ;
        RECT 925.590 108.500 925.910 108.560 ;
        RECT 2415.070 108.500 2415.390 108.560 ;
      LAYER via ;
        RECT 925.620 375.740 925.880 376.000 ;
        RECT 929.760 375.740 930.020 376.000 ;
        RECT 925.620 108.500 925.880 108.760 ;
        RECT 2415.100 108.500 2415.360 108.760 ;
      LAYER met2 ;
        RECT 931.030 400.250 931.310 404.000 ;
        RECT 929.820 400.110 931.310 400.250 ;
        RECT 929.820 376.030 929.960 400.110 ;
        RECT 931.030 400.000 931.310 400.110 ;
        RECT 925.620 375.710 925.880 376.030 ;
        RECT 929.760 375.710 930.020 376.030 ;
        RECT 925.680 108.790 925.820 375.710 ;
        RECT 925.620 108.470 925.880 108.790 ;
        RECT 2415.100 108.470 2415.360 108.790 ;
        RECT 2415.160 82.870 2415.300 108.470 ;
        RECT 2415.160 82.730 2420.360 82.870 ;
        RECT 2420.220 2.400 2420.360 82.730 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.950 108.360 933.270 108.420 ;
        RECT 2435.770 108.360 2436.090 108.420 ;
        RECT 932.950 108.220 2436.090 108.360 ;
        RECT 932.950 108.160 933.270 108.220 ;
        RECT 2435.770 108.160 2436.090 108.220 ;
      LAYER via ;
        RECT 932.980 108.160 933.240 108.420 ;
        RECT 2435.800 108.160 2436.060 108.420 ;
      LAYER met2 ;
        RECT 936.090 400.250 936.370 404.000 ;
        RECT 934.880 400.110 936.370 400.250 ;
        RECT 934.880 324.370 935.020 400.110 ;
        RECT 936.090 400.000 936.370 400.110 ;
        RECT 933.040 324.230 935.020 324.370 ;
        RECT 933.040 108.450 933.180 324.230 ;
        RECT 932.980 108.130 933.240 108.450 ;
        RECT 2435.800 108.130 2436.060 108.450 ;
        RECT 2435.860 1.770 2436.000 108.130 ;
        RECT 2437.950 1.770 2438.510 2.400 ;
        RECT 2435.860 1.630 2438.510 1.770 ;
        RECT 2437.950 -4.800 2438.510 1.630 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 939.390 108.020 939.710 108.080 ;
        RECT 2449.570 108.020 2449.890 108.080 ;
        RECT 939.390 107.880 2449.890 108.020 ;
        RECT 939.390 107.820 939.710 107.880 ;
        RECT 2449.570 107.820 2449.890 107.880 ;
        RECT 2449.570 17.580 2449.890 17.640 ;
        RECT 2453.710 17.580 2454.030 17.640 ;
        RECT 2449.570 17.440 2454.030 17.580 ;
        RECT 2449.570 17.380 2449.890 17.440 ;
        RECT 2453.710 17.380 2454.030 17.440 ;
      LAYER via ;
        RECT 939.420 107.820 939.680 108.080 ;
        RECT 2449.600 107.820 2449.860 108.080 ;
        RECT 2449.600 17.380 2449.860 17.640 ;
        RECT 2453.740 17.380 2454.000 17.640 ;
      LAYER met2 ;
        RECT 941.610 400.250 941.890 404.000 ;
        RECT 940.400 400.110 941.890 400.250 ;
        RECT 940.400 324.370 940.540 400.110 ;
        RECT 941.610 400.000 941.890 400.110 ;
        RECT 939.480 324.230 940.540 324.370 ;
        RECT 939.480 108.110 939.620 324.230 ;
        RECT 939.420 107.790 939.680 108.110 ;
        RECT 2449.600 107.790 2449.860 108.110 ;
        RECT 2449.660 17.670 2449.800 107.790 ;
        RECT 2449.600 17.350 2449.860 17.670 ;
        RECT 2453.740 17.350 2454.000 17.670 ;
        RECT 2453.800 1.770 2453.940 17.350 ;
        RECT 2455.430 1.770 2455.990 2.400 ;
        RECT 2453.800 1.630 2455.990 1.770 ;
        RECT 2455.430 -4.800 2455.990 1.630 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.750 107.680 947.070 107.740 ;
        RECT 2470.270 107.680 2470.590 107.740 ;
        RECT 946.750 107.540 2470.590 107.680 ;
        RECT 946.750 107.480 947.070 107.540 ;
        RECT 2470.270 107.480 2470.590 107.540 ;
      LAYER via ;
        RECT 946.780 107.480 947.040 107.740 ;
        RECT 2470.300 107.480 2470.560 107.740 ;
      LAYER met2 ;
        RECT 947.130 400.250 947.410 404.000 ;
        RECT 946.840 400.110 947.410 400.250 ;
        RECT 946.840 107.770 946.980 400.110 ;
        RECT 947.130 400.000 947.410 400.110 ;
        RECT 946.780 107.450 947.040 107.770 ;
        RECT 2470.300 107.450 2470.560 107.770 ;
        RECT 2470.360 82.870 2470.500 107.450 ;
        RECT 2470.360 82.730 2473.720 82.870 ;
        RECT 2473.580 2.400 2473.720 82.730 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.270 22.340 952.590 22.400 ;
        RECT 2490.970 22.340 2491.290 22.400 ;
        RECT 952.270 22.200 2491.290 22.340 ;
        RECT 952.270 22.140 952.590 22.200 ;
        RECT 2490.970 22.140 2491.290 22.200 ;
      LAYER via ;
        RECT 952.300 22.140 952.560 22.400 ;
        RECT 2491.000 22.140 2491.260 22.400 ;
      LAYER met2 ;
        RECT 952.190 400.180 952.470 404.000 ;
        RECT 952.190 400.000 952.500 400.180 ;
        RECT 952.360 22.430 952.500 400.000 ;
        RECT 952.300 22.110 952.560 22.430 ;
        RECT 2491.000 22.110 2491.260 22.430 ;
        RECT 2491.060 2.400 2491.200 22.110 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.730 376.280 953.050 376.340 ;
        RECT 956.410 376.280 956.730 376.340 ;
        RECT 952.730 376.140 956.730 376.280 ;
        RECT 952.730 376.080 953.050 376.140 ;
        RECT 956.410 376.080 956.730 376.140 ;
        RECT 952.730 22.680 953.050 22.740 ;
        RECT 2508.910 22.680 2509.230 22.740 ;
        RECT 952.730 22.540 2509.230 22.680 ;
        RECT 952.730 22.480 953.050 22.540 ;
        RECT 2508.910 22.480 2509.230 22.540 ;
      LAYER via ;
        RECT 952.760 376.080 953.020 376.340 ;
        RECT 956.440 376.080 956.700 376.340 ;
        RECT 952.760 22.480 953.020 22.740 ;
        RECT 2508.940 22.480 2509.200 22.740 ;
      LAYER met2 ;
        RECT 957.710 400.250 957.990 404.000 ;
        RECT 956.500 400.110 957.990 400.250 ;
        RECT 956.500 376.370 956.640 400.110 ;
        RECT 957.710 400.000 957.990 400.110 ;
        RECT 952.760 376.050 953.020 376.370 ;
        RECT 956.440 376.050 956.700 376.370 ;
        RECT 952.820 22.770 952.960 376.050 ;
        RECT 952.760 22.450 953.020 22.770 ;
        RECT 2508.940 22.450 2509.200 22.770 ;
        RECT 2509.000 2.400 2509.140 22.450 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.170 376.280 959.490 376.340 ;
        RECT 961.930 376.280 962.250 376.340 ;
        RECT 959.170 376.140 962.250 376.280 ;
        RECT 959.170 376.080 959.490 376.140 ;
        RECT 961.930 376.080 962.250 376.140 ;
        RECT 959.170 23.020 959.490 23.080 ;
        RECT 2526.850 23.020 2527.170 23.080 ;
        RECT 959.170 22.880 2527.170 23.020 ;
        RECT 959.170 22.820 959.490 22.880 ;
        RECT 2526.850 22.820 2527.170 22.880 ;
      LAYER via ;
        RECT 959.200 376.080 959.460 376.340 ;
        RECT 961.960 376.080 962.220 376.340 ;
        RECT 959.200 22.820 959.460 23.080 ;
        RECT 2526.880 22.820 2527.140 23.080 ;
      LAYER met2 ;
        RECT 963.230 400.250 963.510 404.000 ;
        RECT 962.020 400.110 963.510 400.250 ;
        RECT 962.020 376.370 962.160 400.110 ;
        RECT 963.230 400.000 963.510 400.110 ;
        RECT 959.200 376.050 959.460 376.370 ;
        RECT 961.960 376.050 962.220 376.370 ;
        RECT 959.260 23.110 959.400 376.050 ;
        RECT 959.200 22.790 959.460 23.110 ;
        RECT 2526.880 22.790 2527.140 23.110 ;
        RECT 2526.940 2.400 2527.080 22.790 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.070 376.280 966.390 376.340 ;
        RECT 967.450 376.280 967.770 376.340 ;
        RECT 966.070 376.140 967.770 376.280 ;
        RECT 966.070 376.080 966.390 376.140 ;
        RECT 967.450 376.080 967.770 376.140 ;
        RECT 966.530 23.360 966.850 23.420 ;
        RECT 2544.330 23.360 2544.650 23.420 ;
        RECT 966.530 23.220 2544.650 23.360 ;
        RECT 966.530 23.160 966.850 23.220 ;
        RECT 2544.330 23.160 2544.650 23.220 ;
      LAYER via ;
        RECT 966.100 376.080 966.360 376.340 ;
        RECT 967.480 376.080 967.740 376.340 ;
        RECT 966.560 23.160 966.820 23.420 ;
        RECT 2544.360 23.160 2544.620 23.420 ;
      LAYER met2 ;
        RECT 968.290 400.250 968.570 404.000 ;
        RECT 967.540 400.110 968.570 400.250 ;
        RECT 967.540 376.370 967.680 400.110 ;
        RECT 968.290 400.000 968.570 400.110 ;
        RECT 966.100 376.050 966.360 376.370 ;
        RECT 967.480 376.050 967.740 376.370 ;
        RECT 966.160 82.870 966.300 376.050 ;
        RECT 966.160 82.730 966.760 82.870 ;
        RECT 966.620 23.450 966.760 82.730 ;
        RECT 966.560 23.130 966.820 23.450 ;
        RECT 2544.360 23.130 2544.620 23.450 ;
        RECT 2544.420 2.400 2544.560 23.130 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.970 23.700 973.290 23.760 ;
        RECT 2562.270 23.700 2562.590 23.760 ;
        RECT 972.970 23.560 2562.590 23.700 ;
        RECT 972.970 23.500 973.290 23.560 ;
        RECT 2562.270 23.500 2562.590 23.560 ;
      LAYER via ;
        RECT 973.000 23.500 973.260 23.760 ;
        RECT 2562.300 23.500 2562.560 23.760 ;
      LAYER met2 ;
        RECT 973.810 400.250 974.090 404.000 ;
        RECT 973.060 400.110 974.090 400.250 ;
        RECT 973.060 23.790 973.200 400.110 ;
        RECT 973.810 400.000 974.090 400.110 ;
        RECT 973.000 23.470 973.260 23.790 ;
        RECT 2562.300 23.470 2562.560 23.790 ;
        RECT 2562.360 2.400 2562.500 23.470 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.590 40.700 442.910 40.760 ;
        RECT 583.350 40.700 583.670 40.760 ;
        RECT 442.590 40.560 583.670 40.700 ;
        RECT 442.590 40.500 442.910 40.560 ;
        RECT 583.350 40.500 583.670 40.560 ;
        RECT 583.350 19.960 583.670 20.020 ;
        RECT 806.450 19.960 806.770 20.020 ;
        RECT 583.350 19.820 806.770 19.960 ;
        RECT 583.350 19.760 583.670 19.820 ;
        RECT 806.450 19.760 806.770 19.820 ;
      LAYER via ;
        RECT 442.620 40.500 442.880 40.760 ;
        RECT 583.380 40.500 583.640 40.760 ;
        RECT 583.380 19.760 583.640 20.020 ;
        RECT 806.480 19.760 806.740 20.020 ;
      LAYER met2 ;
        RECT 443.430 400.250 443.710 404.000 ;
        RECT 442.680 400.110 443.710 400.250 ;
        RECT 442.680 40.790 442.820 400.110 ;
        RECT 443.430 400.000 443.710 400.110 ;
        RECT 442.620 40.470 442.880 40.790 ;
        RECT 583.380 40.470 583.640 40.790 ;
        RECT 583.440 20.050 583.580 40.470 ;
        RECT 583.380 19.730 583.640 20.050 ;
        RECT 806.480 19.730 806.740 20.050 ;
        RECT 806.540 2.400 806.680 19.730 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.430 375.940 973.750 376.000 ;
        RECT 978.030 375.940 978.350 376.000 ;
        RECT 973.430 375.800 978.350 375.940 ;
        RECT 973.430 375.740 973.750 375.800 ;
        RECT 978.030 375.740 978.350 375.800 ;
        RECT 973.430 27.440 973.750 27.500 ;
        RECT 2579.750 27.440 2580.070 27.500 ;
        RECT 973.430 27.300 2580.070 27.440 ;
        RECT 973.430 27.240 973.750 27.300 ;
        RECT 2579.750 27.240 2580.070 27.300 ;
      LAYER via ;
        RECT 973.460 375.740 973.720 376.000 ;
        RECT 978.060 375.740 978.320 376.000 ;
        RECT 973.460 27.240 973.720 27.500 ;
        RECT 2579.780 27.240 2580.040 27.500 ;
      LAYER met2 ;
        RECT 978.870 400.250 979.150 404.000 ;
        RECT 978.120 400.110 979.150 400.250 ;
        RECT 978.120 376.030 978.260 400.110 ;
        RECT 978.870 400.000 979.150 400.110 ;
        RECT 973.460 375.710 973.720 376.030 ;
        RECT 978.060 375.710 978.320 376.030 ;
        RECT 973.520 27.530 973.660 375.710 ;
        RECT 973.460 27.210 973.720 27.530 ;
        RECT 2579.780 27.210 2580.040 27.530 ;
        RECT 2579.840 2.400 2579.980 27.210 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 979.870 380.020 980.190 380.080 ;
        RECT 983.090 380.020 983.410 380.080 ;
        RECT 979.870 379.880 983.410 380.020 ;
        RECT 979.870 379.820 980.190 379.880 ;
        RECT 983.090 379.820 983.410 379.880 ;
        RECT 979.870 27.100 980.190 27.160 ;
        RECT 2597.690 27.100 2598.010 27.160 ;
        RECT 979.870 26.960 2598.010 27.100 ;
        RECT 979.870 26.900 980.190 26.960 ;
        RECT 2597.690 26.900 2598.010 26.960 ;
      LAYER via ;
        RECT 979.900 379.820 980.160 380.080 ;
        RECT 983.120 379.820 983.380 380.080 ;
        RECT 979.900 26.900 980.160 27.160 ;
        RECT 2597.720 26.900 2597.980 27.160 ;
      LAYER met2 ;
        RECT 984.390 400.250 984.670 404.000 ;
        RECT 983.180 400.110 984.670 400.250 ;
        RECT 983.180 380.110 983.320 400.110 ;
        RECT 984.390 400.000 984.670 400.110 ;
        RECT 979.900 379.790 980.160 380.110 ;
        RECT 983.120 379.790 983.380 380.110 ;
        RECT 979.960 27.190 980.100 379.790 ;
        RECT 979.900 26.870 980.160 27.190 ;
        RECT 2597.720 26.870 2597.980 27.190 ;
        RECT 2597.780 2.400 2597.920 26.870 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 986.770 386.480 987.090 386.540 ;
        RECT 988.610 386.480 988.930 386.540 ;
        RECT 986.770 386.340 988.930 386.480 ;
        RECT 986.770 386.280 987.090 386.340 ;
        RECT 988.610 386.280 988.930 386.340 ;
        RECT 986.770 26.760 987.090 26.820 ;
        RECT 2615.170 26.760 2615.490 26.820 ;
        RECT 986.770 26.620 2615.490 26.760 ;
        RECT 986.770 26.560 987.090 26.620 ;
        RECT 2615.170 26.560 2615.490 26.620 ;
      LAYER via ;
        RECT 986.800 386.280 987.060 386.540 ;
        RECT 988.640 386.280 988.900 386.540 ;
        RECT 986.800 26.560 987.060 26.820 ;
        RECT 2615.200 26.560 2615.460 26.820 ;
      LAYER met2 ;
        RECT 989.910 400.250 990.190 404.000 ;
        RECT 988.700 400.110 990.190 400.250 ;
        RECT 988.700 386.570 988.840 400.110 ;
        RECT 989.910 400.000 990.190 400.110 ;
        RECT 986.800 386.250 987.060 386.570 ;
        RECT 988.640 386.250 988.900 386.570 ;
        RECT 986.860 26.850 987.000 386.250 ;
        RECT 986.800 26.530 987.060 26.850 ;
        RECT 2615.200 26.530 2615.460 26.850 ;
        RECT 2615.260 2.400 2615.400 26.530 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 993.670 26.420 993.990 26.480 ;
        RECT 2633.110 26.420 2633.430 26.480 ;
        RECT 993.670 26.280 2633.430 26.420 ;
        RECT 993.670 26.220 993.990 26.280 ;
        RECT 2633.110 26.220 2633.430 26.280 ;
      LAYER via ;
        RECT 993.700 26.220 993.960 26.480 ;
        RECT 2633.140 26.220 2633.400 26.480 ;
      LAYER met2 ;
        RECT 994.970 400.180 995.250 404.000 ;
        RECT 994.970 400.000 995.280 400.180 ;
        RECT 995.140 386.650 995.280 400.000 ;
        RECT 993.760 386.510 995.280 386.650 ;
        RECT 993.760 26.510 993.900 386.510 ;
        RECT 993.700 26.190 993.960 26.510 ;
        RECT 2633.140 26.190 2633.400 26.510 ;
        RECT 2633.200 2.400 2633.340 26.190 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.570 26.080 1000.890 26.140 ;
        RECT 2650.590 26.080 2650.910 26.140 ;
        RECT 1000.570 25.940 2650.910 26.080 ;
        RECT 1000.570 25.880 1000.890 25.940 ;
        RECT 2650.590 25.880 2650.910 25.940 ;
      LAYER via ;
        RECT 1000.600 25.880 1000.860 26.140 ;
        RECT 2650.620 25.880 2650.880 26.140 ;
      LAYER met2 ;
        RECT 1000.490 400.180 1000.770 404.000 ;
        RECT 1000.490 400.000 1000.800 400.180 ;
        RECT 1000.660 26.170 1000.800 400.000 ;
        RECT 1000.600 25.850 1000.860 26.170 ;
        RECT 2650.620 25.850 2650.880 26.170 ;
        RECT 2650.680 2.400 2650.820 25.850 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.030 386.480 1001.350 386.540 ;
        RECT 1004.710 386.480 1005.030 386.540 ;
        RECT 1001.030 386.340 1005.030 386.480 ;
        RECT 1001.030 386.280 1001.350 386.340 ;
        RECT 1004.710 386.280 1005.030 386.340 ;
        RECT 1001.030 25.740 1001.350 25.800 ;
        RECT 2668.530 25.740 2668.850 25.800 ;
        RECT 1001.030 25.600 2668.850 25.740 ;
        RECT 1001.030 25.540 1001.350 25.600 ;
        RECT 2668.530 25.540 2668.850 25.600 ;
      LAYER via ;
        RECT 1001.060 386.280 1001.320 386.540 ;
        RECT 1004.740 386.280 1005.000 386.540 ;
        RECT 1001.060 25.540 1001.320 25.800 ;
        RECT 2668.560 25.540 2668.820 25.800 ;
      LAYER met2 ;
        RECT 1006.010 400.250 1006.290 404.000 ;
        RECT 1004.800 400.110 1006.290 400.250 ;
        RECT 1004.800 386.570 1004.940 400.110 ;
        RECT 1006.010 400.000 1006.290 400.110 ;
        RECT 1001.060 386.250 1001.320 386.570 ;
        RECT 1004.740 386.250 1005.000 386.570 ;
        RECT 1001.120 25.830 1001.260 386.250 ;
        RECT 1001.060 25.510 1001.320 25.830 ;
        RECT 2668.560 25.510 2668.820 25.830 ;
        RECT 2668.620 2.400 2668.760 25.510 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.470 386.480 1007.790 386.540 ;
        RECT 1009.770 386.480 1010.090 386.540 ;
        RECT 1007.470 386.340 1010.090 386.480 ;
        RECT 1007.470 386.280 1007.790 386.340 ;
        RECT 1009.770 386.280 1010.090 386.340 ;
        RECT 1007.470 25.400 1007.790 25.460 ;
        RECT 2686.010 25.400 2686.330 25.460 ;
        RECT 1007.470 25.260 2686.330 25.400 ;
        RECT 1007.470 25.200 1007.790 25.260 ;
        RECT 2686.010 25.200 2686.330 25.260 ;
      LAYER via ;
        RECT 1007.500 386.280 1007.760 386.540 ;
        RECT 1009.800 386.280 1010.060 386.540 ;
        RECT 1007.500 25.200 1007.760 25.460 ;
        RECT 2686.040 25.200 2686.300 25.460 ;
      LAYER met2 ;
        RECT 1011.070 400.250 1011.350 404.000 ;
        RECT 1009.860 400.110 1011.350 400.250 ;
        RECT 1009.860 386.570 1010.000 400.110 ;
        RECT 1011.070 400.000 1011.350 400.110 ;
        RECT 1007.500 386.250 1007.760 386.570 ;
        RECT 1009.800 386.250 1010.060 386.570 ;
        RECT 1007.560 25.490 1007.700 386.250 ;
        RECT 1007.500 25.170 1007.760 25.490 ;
        RECT 2686.040 25.170 2686.300 25.490 ;
        RECT 2686.100 2.400 2686.240 25.170 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.370 386.480 1014.690 386.540 ;
        RECT 1015.750 386.480 1016.070 386.540 ;
        RECT 1014.370 386.340 1016.070 386.480 ;
        RECT 1014.370 386.280 1014.690 386.340 ;
        RECT 1015.750 386.280 1016.070 386.340 ;
        RECT 1014.370 25.060 1014.690 25.120 ;
        RECT 2703.950 25.060 2704.270 25.120 ;
        RECT 1014.370 24.920 2704.270 25.060 ;
        RECT 1014.370 24.860 1014.690 24.920 ;
        RECT 2703.950 24.860 2704.270 24.920 ;
      LAYER via ;
        RECT 1014.400 386.280 1014.660 386.540 ;
        RECT 1015.780 386.280 1016.040 386.540 ;
        RECT 1014.400 24.860 1014.660 25.120 ;
        RECT 2703.980 24.860 2704.240 25.120 ;
      LAYER met2 ;
        RECT 1016.590 400.250 1016.870 404.000 ;
        RECT 1015.840 400.110 1016.870 400.250 ;
        RECT 1015.840 386.570 1015.980 400.110 ;
        RECT 1016.590 400.000 1016.870 400.110 ;
        RECT 1014.400 386.250 1014.660 386.570 ;
        RECT 1015.780 386.250 1016.040 386.570 ;
        RECT 1014.460 25.150 1014.600 386.250 ;
        RECT 1014.400 24.830 1014.660 25.150 ;
        RECT 2703.980 24.830 2704.240 25.150 ;
        RECT 2704.040 2.400 2704.180 24.830 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.730 24.720 1022.050 24.780 ;
        RECT 2721.890 24.720 2722.210 24.780 ;
        RECT 1021.730 24.580 2722.210 24.720 ;
        RECT 1021.730 24.520 1022.050 24.580 ;
        RECT 2721.890 24.520 2722.210 24.580 ;
      LAYER via ;
        RECT 1021.760 24.520 1022.020 24.780 ;
        RECT 2721.920 24.520 2722.180 24.780 ;
      LAYER met2 ;
        RECT 1022.110 400.250 1022.390 404.000 ;
        RECT 1021.820 400.110 1022.390 400.250 ;
        RECT 1021.820 24.810 1021.960 400.110 ;
        RECT 1022.110 400.000 1022.390 400.110 ;
        RECT 1021.760 24.490 1022.020 24.810 ;
        RECT 2721.920 24.490 2722.180 24.810 ;
        RECT 2721.980 2.400 2722.120 24.490 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.270 386.480 1021.590 386.540 ;
        RECT 1025.870 386.480 1026.190 386.540 ;
        RECT 1021.270 386.340 1026.190 386.480 ;
        RECT 1021.270 386.280 1021.590 386.340 ;
        RECT 1025.870 386.280 1026.190 386.340 ;
        RECT 1021.270 24.380 1021.590 24.440 ;
        RECT 2739.370 24.380 2739.690 24.440 ;
        RECT 1021.270 24.240 2739.690 24.380 ;
        RECT 1021.270 24.180 1021.590 24.240 ;
        RECT 2739.370 24.180 2739.690 24.240 ;
      LAYER via ;
        RECT 1021.300 386.280 1021.560 386.540 ;
        RECT 1025.900 386.280 1026.160 386.540 ;
        RECT 1021.300 24.180 1021.560 24.440 ;
        RECT 2739.400 24.180 2739.660 24.440 ;
      LAYER met2 ;
        RECT 1027.170 400.250 1027.450 404.000 ;
        RECT 1025.960 400.110 1027.450 400.250 ;
        RECT 1025.960 386.570 1026.100 400.110 ;
        RECT 1027.170 400.000 1027.450 400.110 ;
        RECT 1021.300 386.250 1021.560 386.570 ;
        RECT 1025.900 386.250 1026.160 386.570 ;
        RECT 1021.360 24.470 1021.500 386.250 ;
        RECT 1021.300 24.150 1021.560 24.470 ;
        RECT 2739.400 24.150 2739.660 24.470 ;
        RECT 2739.460 2.400 2739.600 24.150 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 389.200 448.890 389.260 ;
        RECT 590.710 389.200 591.030 389.260 ;
        RECT 448.570 389.060 591.030 389.200 ;
        RECT 448.570 389.000 448.890 389.060 ;
        RECT 590.710 389.000 591.030 389.060 ;
        RECT 589.790 19.280 590.110 19.340 ;
        RECT 824.390 19.280 824.710 19.340 ;
        RECT 589.790 19.140 824.710 19.280 ;
        RECT 589.790 19.080 590.110 19.140 ;
        RECT 824.390 19.080 824.710 19.140 ;
      LAYER via ;
        RECT 448.600 389.000 448.860 389.260 ;
        RECT 590.740 389.000 591.000 389.260 ;
        RECT 589.820 19.080 590.080 19.340 ;
        RECT 824.420 19.080 824.680 19.340 ;
      LAYER met2 ;
        RECT 448.490 400.180 448.770 404.000 ;
        RECT 448.490 400.000 448.800 400.180 ;
        RECT 448.660 389.290 448.800 400.000 ;
        RECT 448.600 388.970 448.860 389.290 ;
        RECT 590.740 388.970 591.000 389.290 ;
        RECT 590.800 324.370 590.940 388.970 ;
        RECT 589.880 324.230 590.940 324.370 ;
        RECT 589.880 19.370 590.020 324.230 ;
        RECT 589.820 19.050 590.080 19.370 ;
        RECT 824.420 19.050 824.680 19.370 ;
        RECT 824.480 2.400 824.620 19.050 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.170 376.280 1028.490 376.340 ;
        RECT 1031.390 376.280 1031.710 376.340 ;
        RECT 1028.170 376.140 1031.710 376.280 ;
        RECT 1028.170 376.080 1028.490 376.140 ;
        RECT 1031.390 376.080 1031.710 376.140 ;
        RECT 1028.170 24.040 1028.490 24.100 ;
        RECT 2757.310 24.040 2757.630 24.100 ;
        RECT 1028.170 23.900 2757.630 24.040 ;
        RECT 1028.170 23.840 1028.490 23.900 ;
        RECT 2757.310 23.840 2757.630 23.900 ;
      LAYER via ;
        RECT 1028.200 376.080 1028.460 376.340 ;
        RECT 1031.420 376.080 1031.680 376.340 ;
        RECT 1028.200 23.840 1028.460 24.100 ;
        RECT 2757.340 23.840 2757.600 24.100 ;
      LAYER met2 ;
        RECT 1032.690 400.250 1032.970 404.000 ;
        RECT 1031.480 400.110 1032.970 400.250 ;
        RECT 1031.480 376.370 1031.620 400.110 ;
        RECT 1032.690 400.000 1032.970 400.110 ;
        RECT 1028.200 376.050 1028.460 376.370 ;
        RECT 1031.420 376.050 1031.680 376.370 ;
        RECT 1028.260 24.130 1028.400 376.050 ;
        RECT 1028.200 23.810 1028.460 24.130 ;
        RECT 2757.340 23.810 2757.600 24.130 ;
        RECT 2757.400 2.400 2757.540 23.810 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.070 392.940 1035.390 393.000 ;
        RECT 1038.290 392.940 1038.610 393.000 ;
        RECT 1035.070 392.800 1038.610 392.940 ;
        RECT 1035.070 392.740 1035.390 392.800 ;
        RECT 1038.290 392.740 1038.610 392.800 ;
      LAYER via ;
        RECT 1035.100 392.740 1035.360 393.000 ;
        RECT 1038.320 392.740 1038.580 393.000 ;
      LAYER met2 ;
        RECT 1038.210 400.180 1038.490 404.000 ;
        RECT 1038.210 400.000 1038.520 400.180 ;
        RECT 1038.380 393.030 1038.520 400.000 ;
        RECT 1035.100 392.710 1035.360 393.030 ;
        RECT 1038.320 392.710 1038.580 393.030 ;
        RECT 1035.160 24.325 1035.300 392.710 ;
        RECT 1035.090 23.955 1035.370 24.325 ;
        RECT 2774.810 23.955 2775.090 24.325 ;
        RECT 2774.880 2.400 2775.020 23.955 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
      LAYER via2 ;
        RECT 1035.090 24.000 1035.370 24.280 ;
        RECT 2774.810 24.000 2775.090 24.280 ;
      LAYER met3 ;
        RECT 1035.065 24.290 1035.395 24.305 ;
        RECT 2774.785 24.290 2775.115 24.305 ;
        RECT 1035.065 23.990 2775.115 24.290 ;
        RECT 1035.065 23.975 1035.395 23.990 ;
        RECT 2774.785 23.975 2775.115 23.990 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.890 107.340 1043.210 107.400 ;
        RECT 2787.670 107.340 2787.990 107.400 ;
        RECT 1042.890 107.200 2787.990 107.340 ;
        RECT 1042.890 107.140 1043.210 107.200 ;
        RECT 2787.670 107.140 2787.990 107.200 ;
      LAYER via ;
        RECT 1042.920 107.140 1043.180 107.400 ;
        RECT 2787.700 107.140 2787.960 107.400 ;
      LAYER met2 ;
        RECT 1043.270 400.250 1043.550 404.000 ;
        RECT 1042.980 400.110 1043.550 400.250 ;
        RECT 1042.980 107.430 1043.120 400.110 ;
        RECT 1043.270 400.000 1043.550 400.110 ;
        RECT 1042.920 107.110 1043.180 107.430 ;
        RECT 2787.700 107.110 2787.960 107.430 ;
        RECT 2787.760 82.870 2787.900 107.110 ;
        RECT 2787.760 82.730 2792.960 82.870 ;
        RECT 2792.820 2.400 2792.960 82.730 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.790 107.000 1050.110 107.060 ;
        RECT 2808.370 107.000 2808.690 107.060 ;
        RECT 1049.790 106.860 2808.690 107.000 ;
        RECT 1049.790 106.800 1050.110 106.860 ;
        RECT 2808.370 106.800 2808.690 106.860 ;
      LAYER via ;
        RECT 1049.820 106.800 1050.080 107.060 ;
        RECT 2808.400 106.800 2808.660 107.060 ;
      LAYER met2 ;
        RECT 1048.790 400.250 1049.070 404.000 ;
        RECT 1048.790 400.110 1050.020 400.250 ;
        RECT 1048.790 400.000 1049.070 400.110 ;
        RECT 1049.880 107.090 1050.020 400.110 ;
        RECT 1049.820 106.770 1050.080 107.090 ;
        RECT 2808.400 106.770 2808.660 107.090 ;
        RECT 2808.460 82.870 2808.600 106.770 ;
        RECT 2808.460 82.730 2810.440 82.870 ;
        RECT 2810.300 2.400 2810.440 82.730 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2822.170 17.580 2822.490 17.640 ;
        RECT 2826.310 17.580 2826.630 17.640 ;
        RECT 2822.170 17.440 2826.630 17.580 ;
        RECT 2822.170 17.380 2822.490 17.440 ;
        RECT 2826.310 17.380 2826.630 17.440 ;
      LAYER via ;
        RECT 2822.200 17.380 2822.460 17.640 ;
        RECT 2826.340 17.380 2826.600 17.640 ;
      LAYER met2 ;
        RECT 1054.310 400.250 1054.590 404.000 ;
        RECT 1053.100 400.110 1054.590 400.250 ;
        RECT 1053.100 324.370 1053.240 400.110 ;
        RECT 1054.310 400.000 1054.590 400.110 ;
        RECT 1050.340 324.230 1053.240 324.370 ;
        RECT 1050.340 107.285 1050.480 324.230 ;
        RECT 1050.270 106.915 1050.550 107.285 ;
        RECT 2822.190 106.915 2822.470 107.285 ;
        RECT 2822.260 17.670 2822.400 106.915 ;
        RECT 2822.200 17.350 2822.460 17.670 ;
        RECT 2826.340 17.350 2826.600 17.670 ;
        RECT 2826.400 1.770 2826.540 17.350 ;
        RECT 2828.030 1.770 2828.590 2.400 ;
        RECT 2826.400 1.630 2828.590 1.770 ;
        RECT 2828.030 -4.800 2828.590 1.630 ;
      LAYER via2 ;
        RECT 1050.270 106.960 1050.550 107.240 ;
        RECT 2822.190 106.960 2822.470 107.240 ;
      LAYER met3 ;
        RECT 1050.245 107.250 1050.575 107.265 ;
        RECT 2822.165 107.250 2822.495 107.265 ;
        RECT 1050.245 106.950 2822.495 107.250 ;
        RECT 1050.245 106.935 1050.575 106.950 ;
        RECT 2822.165 106.935 2822.495 106.950 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.770 376.280 1056.090 376.340 ;
        RECT 1058.070 376.280 1058.390 376.340 ;
        RECT 1055.770 376.140 1058.390 376.280 ;
        RECT 1055.770 376.080 1056.090 376.140 ;
        RECT 1058.070 376.080 1058.390 376.140 ;
        RECT 1055.770 31.860 1056.090 31.920 ;
        RECT 2845.630 31.860 2845.950 31.920 ;
        RECT 1055.770 31.720 2845.950 31.860 ;
        RECT 1055.770 31.660 1056.090 31.720 ;
        RECT 2845.630 31.660 2845.950 31.720 ;
      LAYER via ;
        RECT 1055.800 376.080 1056.060 376.340 ;
        RECT 1058.100 376.080 1058.360 376.340 ;
        RECT 1055.800 31.660 1056.060 31.920 ;
        RECT 2845.660 31.660 2845.920 31.920 ;
      LAYER met2 ;
        RECT 1059.370 400.250 1059.650 404.000 ;
        RECT 1058.160 400.110 1059.650 400.250 ;
        RECT 1058.160 376.370 1058.300 400.110 ;
        RECT 1059.370 400.000 1059.650 400.110 ;
        RECT 1055.800 376.050 1056.060 376.370 ;
        RECT 1058.100 376.050 1058.360 376.370 ;
        RECT 1055.860 31.950 1056.000 376.050 ;
        RECT 1055.800 31.630 1056.060 31.950 ;
        RECT 2845.660 31.630 2845.920 31.950 ;
        RECT 2845.720 2.400 2845.860 31.630 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1062.670 376.280 1062.990 376.340 ;
        RECT 1064.050 376.280 1064.370 376.340 ;
        RECT 1062.670 376.140 1064.370 376.280 ;
        RECT 1062.670 376.080 1062.990 376.140 ;
        RECT 1064.050 376.080 1064.370 376.140 ;
        RECT 1062.670 31.520 1062.990 31.580 ;
        RECT 2863.570 31.520 2863.890 31.580 ;
        RECT 1062.670 31.380 2863.890 31.520 ;
        RECT 1062.670 31.320 1062.990 31.380 ;
        RECT 2863.570 31.320 2863.890 31.380 ;
      LAYER via ;
        RECT 1062.700 376.080 1062.960 376.340 ;
        RECT 1064.080 376.080 1064.340 376.340 ;
        RECT 1062.700 31.320 1062.960 31.580 ;
        RECT 2863.600 31.320 2863.860 31.580 ;
      LAYER met2 ;
        RECT 1064.890 400.250 1065.170 404.000 ;
        RECT 1064.140 400.110 1065.170 400.250 ;
        RECT 1064.140 376.370 1064.280 400.110 ;
        RECT 1064.890 400.000 1065.170 400.110 ;
        RECT 1062.700 376.050 1062.960 376.370 ;
        RECT 1064.080 376.050 1064.340 376.370 ;
        RECT 1062.760 31.610 1062.900 376.050 ;
        RECT 1062.700 31.290 1062.960 31.610 ;
        RECT 2863.600 31.290 2863.860 31.610 ;
        RECT 2863.660 2.400 2863.800 31.290 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.570 31.180 1069.890 31.240 ;
        RECT 2881.510 31.180 2881.830 31.240 ;
        RECT 1069.570 31.040 2881.830 31.180 ;
        RECT 1069.570 30.980 1069.890 31.040 ;
        RECT 2881.510 30.980 2881.830 31.040 ;
      LAYER via ;
        RECT 1069.600 30.980 1069.860 31.240 ;
        RECT 2881.540 30.980 2881.800 31.240 ;
      LAYER met2 ;
        RECT 1069.950 400.250 1070.230 404.000 ;
        RECT 1069.660 400.110 1070.230 400.250 ;
        RECT 1069.660 31.270 1069.800 400.110 ;
        RECT 1069.950 400.000 1070.230 400.110 ;
        RECT 1069.600 30.950 1069.860 31.270 ;
        RECT 2881.540 30.950 2881.800 31.270 ;
        RECT 2881.600 2.400 2881.740 30.950 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 385.800 449.350 385.860 ;
        RECT 452.710 385.800 453.030 385.860 ;
        RECT 449.030 385.660 453.030 385.800 ;
        RECT 449.030 385.600 449.350 385.660 ;
        RECT 452.710 385.600 453.030 385.660 ;
        RECT 449.030 40.360 449.350 40.420 ;
        RECT 596.230 40.360 596.550 40.420 ;
        RECT 449.030 40.220 596.550 40.360 ;
        RECT 449.030 40.160 449.350 40.220 ;
        RECT 596.230 40.160 596.550 40.220 ;
        RECT 596.230 18.600 596.550 18.660 ;
        RECT 841.870 18.600 842.190 18.660 ;
        RECT 596.230 18.460 842.190 18.600 ;
        RECT 596.230 18.400 596.550 18.460 ;
        RECT 841.870 18.400 842.190 18.460 ;
      LAYER via ;
        RECT 449.060 385.600 449.320 385.860 ;
        RECT 452.740 385.600 453.000 385.860 ;
        RECT 449.060 40.160 449.320 40.420 ;
        RECT 596.260 40.160 596.520 40.420 ;
        RECT 596.260 18.400 596.520 18.660 ;
        RECT 841.900 18.400 842.160 18.660 ;
      LAYER met2 ;
        RECT 454.010 400.250 454.290 404.000 ;
        RECT 452.800 400.110 454.290 400.250 ;
        RECT 452.800 385.890 452.940 400.110 ;
        RECT 454.010 400.000 454.290 400.110 ;
        RECT 449.060 385.570 449.320 385.890 ;
        RECT 452.740 385.570 453.000 385.890 ;
        RECT 449.120 40.450 449.260 385.570 ;
        RECT 449.060 40.130 449.320 40.450 ;
        RECT 596.260 40.130 596.520 40.450 ;
        RECT 596.320 18.690 596.460 40.130 ;
        RECT 596.260 18.370 596.520 18.690 ;
        RECT 841.900 18.370 842.160 18.690 ;
        RECT 841.960 2.400 842.100 18.370 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 459.610 388.860 459.930 388.920 ;
        RECT 596.690 388.860 597.010 388.920 ;
        RECT 459.610 388.720 597.010 388.860 ;
        RECT 459.610 388.660 459.930 388.720 ;
        RECT 596.690 388.660 597.010 388.720 ;
        RECT 596.690 18.260 597.010 18.320 ;
        RECT 859.810 18.260 860.130 18.320 ;
        RECT 596.690 18.120 860.130 18.260 ;
        RECT 596.690 18.060 597.010 18.120 ;
        RECT 859.810 18.060 860.130 18.120 ;
      LAYER via ;
        RECT 459.640 388.660 459.900 388.920 ;
        RECT 596.720 388.660 596.980 388.920 ;
        RECT 596.720 18.060 596.980 18.320 ;
        RECT 859.840 18.060 860.100 18.320 ;
      LAYER met2 ;
        RECT 459.530 400.180 459.810 404.000 ;
        RECT 459.530 400.000 459.840 400.180 ;
        RECT 459.700 388.950 459.840 400.000 ;
        RECT 459.640 388.630 459.900 388.950 ;
        RECT 596.720 388.630 596.980 388.950 ;
        RECT 596.780 18.350 596.920 388.630 ;
        RECT 596.720 18.030 596.980 18.350 ;
        RECT 859.840 18.030 860.100 18.350 ;
        RECT 859.900 2.400 860.040 18.030 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 464.670 388.520 464.990 388.580 ;
        RECT 603.590 388.520 603.910 388.580 ;
        RECT 464.670 388.380 603.910 388.520 ;
        RECT 464.670 388.320 464.990 388.380 ;
        RECT 603.590 388.320 603.910 388.380 ;
        RECT 603.590 17.920 603.910 17.980 ;
        RECT 877.290 17.920 877.610 17.980 ;
        RECT 603.590 17.780 877.610 17.920 ;
        RECT 603.590 17.720 603.910 17.780 ;
        RECT 877.290 17.720 877.610 17.780 ;
      LAYER via ;
        RECT 464.700 388.320 464.960 388.580 ;
        RECT 603.620 388.320 603.880 388.580 ;
        RECT 603.620 17.720 603.880 17.980 ;
        RECT 877.320 17.720 877.580 17.980 ;
      LAYER met2 ;
        RECT 464.590 400.180 464.870 404.000 ;
        RECT 464.590 400.000 464.900 400.180 ;
        RECT 464.760 388.610 464.900 400.000 ;
        RECT 464.700 388.290 464.960 388.610 ;
        RECT 603.620 388.290 603.880 388.610 ;
        RECT 603.680 18.010 603.820 388.290 ;
        RECT 603.620 17.690 603.880 18.010 ;
        RECT 877.320 17.690 877.580 18.010 ;
        RECT 877.380 2.400 877.520 17.690 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 26.420 469.590 26.480 ;
        RECT 895.230 26.420 895.550 26.480 ;
        RECT 469.270 26.280 895.550 26.420 ;
        RECT 469.270 26.220 469.590 26.280 ;
        RECT 895.230 26.220 895.550 26.280 ;
      LAYER via ;
        RECT 469.300 26.220 469.560 26.480 ;
        RECT 895.260 26.220 895.520 26.480 ;
      LAYER met2 ;
        RECT 470.110 400.250 470.390 404.000 ;
        RECT 469.360 400.110 470.390 400.250 ;
        RECT 469.360 26.510 469.500 400.110 ;
        RECT 470.110 400.000 470.390 400.110 ;
        RECT 469.300 26.190 469.560 26.510 ;
        RECT 895.260 26.190 895.520 26.510 ;
        RECT 895.320 2.400 895.460 26.190 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.730 386.140 470.050 386.200 ;
        RECT 474.330 386.140 474.650 386.200 ;
        RECT 469.730 386.000 474.650 386.140 ;
        RECT 469.730 385.940 470.050 386.000 ;
        RECT 474.330 385.940 474.650 386.000 ;
        RECT 469.730 26.080 470.050 26.140 ;
        RECT 912.710 26.080 913.030 26.140 ;
        RECT 469.730 25.940 913.030 26.080 ;
        RECT 469.730 25.880 470.050 25.940 ;
        RECT 912.710 25.880 913.030 25.940 ;
      LAYER via ;
        RECT 469.760 385.940 470.020 386.200 ;
        RECT 474.360 385.940 474.620 386.200 ;
        RECT 469.760 25.880 470.020 26.140 ;
        RECT 912.740 25.880 913.000 26.140 ;
      LAYER met2 ;
        RECT 475.170 400.250 475.450 404.000 ;
        RECT 474.420 400.110 475.450 400.250 ;
        RECT 474.420 386.230 474.560 400.110 ;
        RECT 475.170 400.000 475.450 400.110 ;
        RECT 469.760 385.910 470.020 386.230 ;
        RECT 474.360 385.910 474.620 386.230 ;
        RECT 469.820 26.170 469.960 385.910 ;
        RECT 469.760 25.850 470.020 26.170 ;
        RECT 912.740 25.850 913.000 26.170 ;
        RECT 912.800 2.400 912.940 25.850 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 25.740 476.490 25.800 ;
        RECT 930.650 25.740 930.970 25.800 ;
        RECT 476.170 25.600 930.970 25.740 ;
        RECT 476.170 25.540 476.490 25.600 ;
        RECT 930.650 25.540 930.970 25.600 ;
      LAYER via ;
        RECT 476.200 25.540 476.460 25.800 ;
        RECT 930.680 25.540 930.940 25.800 ;
      LAYER met2 ;
        RECT 480.690 400.250 480.970 404.000 ;
        RECT 479.480 400.110 480.970 400.250 ;
        RECT 479.480 386.650 479.620 400.110 ;
        RECT 480.690 400.000 480.970 400.110 ;
        RECT 476.260 386.510 479.620 386.650 ;
        RECT 476.260 25.830 476.400 386.510 ;
        RECT 476.200 25.510 476.460 25.830 ;
        RECT 930.680 25.510 930.940 25.830 ;
        RECT 930.740 2.400 930.880 25.510 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 386.480 483.390 386.540 ;
        RECT 484.910 386.480 485.230 386.540 ;
        RECT 483.070 386.340 485.230 386.480 ;
        RECT 483.070 386.280 483.390 386.340 ;
        RECT 484.910 386.280 485.230 386.340 ;
        RECT 483.070 25.400 483.390 25.460 ;
        RECT 948.590 25.400 948.910 25.460 ;
        RECT 483.070 25.260 948.910 25.400 ;
        RECT 483.070 25.200 483.390 25.260 ;
        RECT 948.590 25.200 948.910 25.260 ;
      LAYER via ;
        RECT 483.100 386.280 483.360 386.540 ;
        RECT 484.940 386.280 485.200 386.540 ;
        RECT 483.100 25.200 483.360 25.460 ;
        RECT 948.620 25.200 948.880 25.460 ;
      LAYER met2 ;
        RECT 486.210 400.250 486.490 404.000 ;
        RECT 485.000 400.110 486.490 400.250 ;
        RECT 485.000 386.570 485.140 400.110 ;
        RECT 486.210 400.000 486.490 400.110 ;
        RECT 483.100 386.250 483.360 386.570 ;
        RECT 484.940 386.250 485.200 386.570 ;
        RECT 483.160 25.490 483.300 386.250 ;
        RECT 483.100 25.170 483.360 25.490 ;
        RECT 948.620 25.170 948.880 25.490 ;
        RECT 948.680 2.400 948.820 25.170 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 386.480 490.290 386.540 ;
        RECT 491.350 386.480 491.670 386.540 ;
        RECT 489.970 386.340 491.670 386.480 ;
        RECT 489.970 386.280 490.290 386.340 ;
        RECT 491.350 386.280 491.670 386.340 ;
        RECT 489.970 25.060 490.290 25.120 ;
        RECT 966.070 25.060 966.390 25.120 ;
        RECT 489.970 24.920 966.390 25.060 ;
        RECT 489.970 24.860 490.290 24.920 ;
        RECT 966.070 24.860 966.390 24.920 ;
      LAYER via ;
        RECT 490.000 386.280 490.260 386.540 ;
        RECT 491.380 386.280 491.640 386.540 ;
        RECT 490.000 24.860 490.260 25.120 ;
        RECT 966.100 24.860 966.360 25.120 ;
      LAYER met2 ;
        RECT 491.270 400.180 491.550 404.000 ;
        RECT 491.270 400.000 491.580 400.180 ;
        RECT 491.440 386.570 491.580 400.000 ;
        RECT 490.000 386.250 490.260 386.570 ;
        RECT 491.380 386.250 491.640 386.570 ;
        RECT 490.060 25.150 490.200 386.250 ;
        RECT 490.000 24.830 490.260 25.150 ;
        RECT 966.100 24.830 966.360 25.150 ;
        RECT 966.160 2.400 966.300 24.830 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.490 376.280 1070.810 376.340 ;
        RECT 1074.170 376.280 1074.490 376.340 ;
        RECT 1070.490 376.140 1074.490 376.280 ;
        RECT 1070.490 376.080 1070.810 376.140 ;
        RECT 1074.170 376.080 1074.490 376.140 ;
        RECT 831.290 28.460 831.610 28.520 ;
        RECT 1070.490 28.460 1070.810 28.520 ;
        RECT 831.290 28.320 1070.810 28.460 ;
        RECT 831.290 28.260 831.610 28.320 ;
        RECT 1070.490 28.260 1070.810 28.320 ;
        RECT 641.770 20.640 642.090 20.700 ;
        RECT 646.830 20.640 647.150 20.700 ;
        RECT 831.290 20.640 831.610 20.700 ;
        RECT 641.770 20.500 831.610 20.640 ;
        RECT 641.770 20.440 642.090 20.500 ;
        RECT 646.830 20.440 647.150 20.500 ;
        RECT 831.290 20.440 831.610 20.500 ;
      LAYER via ;
        RECT 1070.520 376.080 1070.780 376.340 ;
        RECT 1074.200 376.080 1074.460 376.340 ;
        RECT 831.320 28.260 831.580 28.520 ;
        RECT 1070.520 28.260 1070.780 28.520 ;
        RECT 641.800 20.440 642.060 20.700 ;
        RECT 646.860 20.440 647.120 20.700 ;
        RECT 831.320 20.440 831.580 20.700 ;
      LAYER met2 ;
        RECT 395.130 400.930 395.410 404.000 ;
        RECT 395.130 400.790 396.360 400.930 ;
        RECT 395.130 400.000 395.410 400.790 ;
        RECT 396.220 351.970 396.360 400.790 ;
        RECT 1075.470 400.250 1075.750 404.000 ;
        RECT 1074.260 400.110 1075.750 400.250 ;
        RECT 1074.260 376.370 1074.400 400.110 ;
        RECT 1075.470 400.000 1075.750 400.110 ;
        RECT 1070.520 376.050 1070.780 376.370 ;
        RECT 1074.200 376.050 1074.460 376.370 ;
        RECT 395.300 351.830 396.360 351.970 ;
        RECT 395.300 24.325 395.440 351.830 ;
        RECT 1070.580 28.550 1070.720 376.050 ;
        RECT 831.320 28.230 831.580 28.550 ;
        RECT 1070.520 28.230 1070.780 28.550 ;
        RECT 395.230 23.955 395.510 24.325 ;
        RECT 641.790 23.955 642.070 24.325 ;
        RECT 641.860 20.730 642.000 23.955 ;
        RECT 831.380 20.730 831.520 28.230 ;
        RECT 641.800 20.410 642.060 20.730 ;
        RECT 646.860 20.410 647.120 20.730 ;
        RECT 831.320 20.410 831.580 20.730 ;
        RECT 646.920 2.400 647.060 20.410 ;
        RECT 646.710 -4.800 647.270 2.400 ;
      LAYER via2 ;
        RECT 395.230 24.000 395.510 24.280 ;
        RECT 641.790 24.000 642.070 24.280 ;
      LAYER met3 ;
        RECT 395.205 24.290 395.535 24.305 ;
        RECT 641.765 24.290 642.095 24.305 ;
        RECT 395.205 23.990 642.095 24.290 ;
        RECT 395.205 23.975 395.535 23.990 ;
        RECT 641.765 23.975 642.095 23.990 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 24.720 497.190 24.780 ;
        RECT 984.010 24.720 984.330 24.780 ;
        RECT 496.870 24.580 984.330 24.720 ;
        RECT 496.870 24.520 497.190 24.580 ;
        RECT 984.010 24.520 984.330 24.580 ;
      LAYER via ;
        RECT 496.900 24.520 497.160 24.780 ;
        RECT 984.040 24.520 984.300 24.780 ;
      LAYER met2 ;
        RECT 496.790 400.180 497.070 404.000 ;
        RECT 496.790 400.000 497.100 400.180 ;
        RECT 496.960 24.810 497.100 400.000 ;
        RECT 496.900 24.490 497.160 24.810 ;
        RECT 984.040 24.490 984.300 24.810 ;
        RECT 984.100 2.400 984.240 24.490 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 386.480 497.650 386.540 ;
        RECT 501.010 386.480 501.330 386.540 ;
        RECT 497.330 386.340 501.330 386.480 ;
        RECT 497.330 386.280 497.650 386.340 ;
        RECT 501.010 386.280 501.330 386.340 ;
        RECT 497.330 24.380 497.650 24.440 ;
        RECT 1001.490 24.380 1001.810 24.440 ;
        RECT 497.330 24.240 1001.810 24.380 ;
        RECT 497.330 24.180 497.650 24.240 ;
        RECT 1001.490 24.180 1001.810 24.240 ;
      LAYER via ;
        RECT 497.360 386.280 497.620 386.540 ;
        RECT 501.040 386.280 501.300 386.540 ;
        RECT 497.360 24.180 497.620 24.440 ;
        RECT 1001.520 24.180 1001.780 24.440 ;
      LAYER met2 ;
        RECT 502.310 400.250 502.590 404.000 ;
        RECT 501.100 400.110 502.590 400.250 ;
        RECT 501.100 386.570 501.240 400.110 ;
        RECT 502.310 400.000 502.590 400.110 ;
        RECT 497.360 386.250 497.620 386.570 ;
        RECT 501.040 386.250 501.300 386.570 ;
        RECT 497.420 24.470 497.560 386.250 ;
        RECT 497.360 24.150 497.620 24.470 ;
        RECT 1001.520 24.150 1001.780 24.470 ;
        RECT 1001.580 2.400 1001.720 24.150 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 386.480 504.090 386.540 ;
        RECT 506.070 386.480 506.390 386.540 ;
        RECT 503.770 386.340 506.390 386.480 ;
        RECT 503.770 386.280 504.090 386.340 ;
        RECT 506.070 386.280 506.390 386.340 ;
        RECT 503.770 24.040 504.090 24.100 ;
        RECT 1019.430 24.040 1019.750 24.100 ;
        RECT 503.770 23.900 1019.750 24.040 ;
        RECT 503.770 23.840 504.090 23.900 ;
        RECT 1019.430 23.840 1019.750 23.900 ;
      LAYER via ;
        RECT 503.800 386.280 504.060 386.540 ;
        RECT 506.100 386.280 506.360 386.540 ;
        RECT 503.800 23.840 504.060 24.100 ;
        RECT 1019.460 23.840 1019.720 24.100 ;
      LAYER met2 ;
        RECT 507.370 400.250 507.650 404.000 ;
        RECT 506.160 400.110 507.650 400.250 ;
        RECT 506.160 386.570 506.300 400.110 ;
        RECT 507.370 400.000 507.650 400.110 ;
        RECT 503.800 386.250 504.060 386.570 ;
        RECT 506.100 386.250 506.360 386.570 ;
        RECT 503.860 24.130 504.000 386.250 ;
        RECT 503.800 23.810 504.060 24.130 ;
        RECT 1019.460 23.810 1019.720 24.130 ;
        RECT 1019.520 2.400 1019.660 23.810 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 386.140 510.990 386.200 ;
        RECT 512.510 386.140 512.830 386.200 ;
        RECT 510.670 386.000 512.830 386.140 ;
        RECT 510.670 385.940 510.990 386.000 ;
        RECT 512.510 385.940 512.830 386.000 ;
      LAYER via ;
        RECT 510.700 385.940 510.960 386.200 ;
        RECT 512.540 385.940 512.800 386.200 ;
      LAYER met2 ;
        RECT 512.890 400.250 513.170 404.000 ;
        RECT 512.600 400.110 513.170 400.250 ;
        RECT 512.600 386.230 512.740 400.110 ;
        RECT 512.890 400.000 513.170 400.110 ;
        RECT 510.700 385.910 510.960 386.230 ;
        RECT 512.540 385.910 512.800 386.230 ;
        RECT 510.760 25.685 510.900 385.910 ;
        RECT 510.690 25.315 510.970 25.685 ;
        RECT 1036.930 25.315 1037.210 25.685 ;
        RECT 1037.000 2.400 1037.140 25.315 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
      LAYER via2 ;
        RECT 510.690 25.360 510.970 25.640 ;
        RECT 1036.930 25.360 1037.210 25.640 ;
      LAYER met3 ;
        RECT 510.665 25.650 510.995 25.665 ;
        RECT 1036.905 25.650 1037.235 25.665 ;
        RECT 510.665 25.350 1037.235 25.650 ;
        RECT 510.665 25.335 510.995 25.350 ;
        RECT 1036.905 25.335 1037.235 25.350 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.410 400.250 518.690 404.000 ;
        RECT 517.660 400.110 518.690 400.250 ;
        RECT 517.660 25.005 517.800 400.110 ;
        RECT 518.410 400.000 518.690 400.110 ;
        RECT 517.590 24.635 517.870 25.005 ;
        RECT 1054.870 24.635 1055.150 25.005 ;
        RECT 1054.940 2.400 1055.080 24.635 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
      LAYER via2 ;
        RECT 517.590 24.680 517.870 24.960 ;
        RECT 1054.870 24.680 1055.150 24.960 ;
      LAYER met3 ;
        RECT 517.565 24.970 517.895 24.985 ;
        RECT 1054.845 24.970 1055.175 24.985 ;
        RECT 517.565 24.670 1055.175 24.970 ;
        RECT 517.565 24.655 517.895 24.670 ;
        RECT 1054.845 24.655 1055.175 24.670 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.490 105.300 518.810 105.360 ;
        RECT 1070.950 105.300 1071.270 105.360 ;
        RECT 518.490 105.160 1071.270 105.300 ;
        RECT 518.490 105.100 518.810 105.160 ;
        RECT 1070.950 105.100 1071.270 105.160 ;
      LAYER via ;
        RECT 518.520 105.100 518.780 105.360 ;
        RECT 1070.980 105.100 1071.240 105.360 ;
      LAYER met2 ;
        RECT 523.470 400.250 523.750 404.000 ;
        RECT 522.260 400.110 523.750 400.250 ;
        RECT 522.260 324.370 522.400 400.110 ;
        RECT 523.470 400.000 523.750 400.110 ;
        RECT 518.580 324.230 522.400 324.370 ;
        RECT 518.580 105.390 518.720 324.230 ;
        RECT 518.520 105.070 518.780 105.390 ;
        RECT 1070.980 105.070 1071.240 105.390 ;
        RECT 1071.040 82.870 1071.180 105.070 ;
        RECT 1071.040 82.730 1072.560 82.870 ;
        RECT 1072.420 2.400 1072.560 82.730 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 529.070 390.560 529.390 390.620 ;
        RECT 756.770 390.560 757.090 390.620 ;
        RECT 529.070 390.420 757.090 390.560 ;
        RECT 529.070 390.360 529.390 390.420 ;
        RECT 756.770 390.360 757.090 390.420 ;
        RECT 755.850 29.140 756.170 29.200 ;
        RECT 1090.730 29.140 1091.050 29.200 ;
        RECT 755.850 29.000 1091.050 29.140 ;
        RECT 755.850 28.940 756.170 29.000 ;
        RECT 1090.730 28.940 1091.050 29.000 ;
      LAYER via ;
        RECT 529.100 390.360 529.360 390.620 ;
        RECT 756.800 390.360 757.060 390.620 ;
        RECT 755.880 28.940 756.140 29.200 ;
        RECT 1090.760 28.940 1091.020 29.200 ;
      LAYER met2 ;
        RECT 528.990 400.180 529.270 404.000 ;
        RECT 528.990 400.000 529.300 400.180 ;
        RECT 529.160 390.650 529.300 400.000 ;
        RECT 529.100 390.330 529.360 390.650 ;
        RECT 756.800 390.330 757.060 390.650 ;
        RECT 756.860 324.370 757.000 390.330 ;
        RECT 755.940 324.230 757.000 324.370 ;
        RECT 755.940 29.230 756.080 324.230 ;
        RECT 755.880 28.910 756.140 29.230 ;
        RECT 1090.760 28.910 1091.020 29.230 ;
        RECT 1090.820 14.690 1090.960 28.910 ;
        RECT 1090.360 14.550 1090.960 14.690 ;
        RECT 1090.360 2.400 1090.500 14.550 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 569.090 393.280 569.410 393.340 ;
        RECT 639.470 393.280 639.790 393.340 ;
        RECT 569.090 393.140 639.790 393.280 ;
        RECT 569.090 393.080 569.410 393.140 ;
        RECT 639.470 393.080 639.790 393.140 ;
        RECT 534.590 388.180 534.910 388.240 ;
        RECT 569.090 388.180 569.410 388.240 ;
        RECT 534.590 388.040 569.410 388.180 ;
        RECT 534.590 387.980 534.910 388.040 ;
        RECT 569.090 387.980 569.410 388.040 ;
        RECT 638.550 29.480 638.870 29.540 ;
        RECT 1107.750 29.480 1108.070 29.540 ;
        RECT 638.550 29.340 1108.070 29.480 ;
        RECT 638.550 29.280 638.870 29.340 ;
        RECT 1107.750 29.280 1108.070 29.340 ;
      LAYER via ;
        RECT 569.120 393.080 569.380 393.340 ;
        RECT 639.500 393.080 639.760 393.340 ;
        RECT 534.620 387.980 534.880 388.240 ;
        RECT 569.120 387.980 569.380 388.240 ;
        RECT 638.580 29.280 638.840 29.540 ;
        RECT 1107.780 29.280 1108.040 29.540 ;
      LAYER met2 ;
        RECT 534.510 400.180 534.790 404.000 ;
        RECT 534.510 400.000 534.820 400.180 ;
        RECT 534.680 388.270 534.820 400.000 ;
        RECT 569.120 393.050 569.380 393.370 ;
        RECT 639.500 393.050 639.760 393.370 ;
        RECT 569.180 388.270 569.320 393.050 ;
        RECT 534.620 387.950 534.880 388.270 ;
        RECT 569.120 387.950 569.380 388.270 ;
        RECT 639.560 324.370 639.700 393.050 ;
        RECT 638.640 324.230 639.700 324.370 ;
        RECT 638.640 29.570 638.780 324.230 ;
        RECT 638.580 29.250 638.840 29.570 ;
        RECT 1107.780 29.250 1108.040 29.570 ;
        RECT 1107.840 2.400 1107.980 29.250 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 29.820 538.590 29.880 ;
        RECT 1125.690 29.820 1126.010 29.880 ;
        RECT 538.270 29.680 1126.010 29.820 ;
        RECT 538.270 29.620 538.590 29.680 ;
        RECT 1125.690 29.620 1126.010 29.680 ;
      LAYER via ;
        RECT 538.300 29.620 538.560 29.880 ;
        RECT 1125.720 29.620 1125.980 29.880 ;
      LAYER met2 ;
        RECT 539.570 400.250 539.850 404.000 ;
        RECT 538.360 400.110 539.850 400.250 ;
        RECT 538.360 29.910 538.500 400.110 ;
        RECT 539.570 400.000 539.850 400.110 ;
        RECT 538.300 29.590 538.560 29.910 ;
        RECT 1125.720 29.590 1125.980 29.910 ;
        RECT 1125.780 2.400 1125.920 29.590 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 30.160 545.490 30.220 ;
        RECT 1143.630 30.160 1143.950 30.220 ;
        RECT 545.170 30.020 1143.950 30.160 ;
        RECT 545.170 29.960 545.490 30.020 ;
        RECT 1143.630 29.960 1143.950 30.020 ;
      LAYER via ;
        RECT 545.200 29.960 545.460 30.220 ;
        RECT 1143.660 29.960 1143.920 30.220 ;
      LAYER met2 ;
        RECT 545.090 400.180 545.370 404.000 ;
        RECT 545.090 400.000 545.400 400.180 ;
        RECT 545.260 30.250 545.400 400.000 ;
        RECT 545.200 29.930 545.460 30.250 ;
        RECT 1143.660 29.930 1143.920 30.250 ;
        RECT 1143.720 2.400 1143.860 29.930 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.730 23.360 401.050 23.420 ;
        RECT 664.770 23.360 665.090 23.420 ;
        RECT 400.730 23.220 665.090 23.360 ;
        RECT 400.730 23.160 401.050 23.220 ;
        RECT 664.770 23.160 665.090 23.220 ;
      LAYER via ;
        RECT 400.760 23.160 401.020 23.420 ;
        RECT 664.800 23.160 665.060 23.420 ;
      LAYER met2 ;
        RECT 400.190 400.250 400.470 404.000 ;
        RECT 400.190 400.110 400.960 400.250 ;
        RECT 400.190 400.000 400.470 400.110 ;
        RECT 400.820 23.450 400.960 400.110 ;
        RECT 400.760 23.130 401.020 23.450 ;
        RECT 664.800 23.130 665.060 23.450 ;
        RECT 664.860 2.400 665.000 23.130 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.630 375.940 545.950 376.000 ;
        RECT 549.310 375.940 549.630 376.000 ;
        RECT 545.630 375.800 549.630 375.940 ;
        RECT 545.630 375.740 545.950 375.800 ;
        RECT 549.310 375.740 549.630 375.800 ;
        RECT 545.630 30.500 545.950 30.560 ;
        RECT 1161.110 30.500 1161.430 30.560 ;
        RECT 545.630 30.360 1161.430 30.500 ;
        RECT 545.630 30.300 545.950 30.360 ;
        RECT 1161.110 30.300 1161.430 30.360 ;
      LAYER via ;
        RECT 545.660 375.740 545.920 376.000 ;
        RECT 549.340 375.740 549.600 376.000 ;
        RECT 545.660 30.300 545.920 30.560 ;
        RECT 1161.140 30.300 1161.400 30.560 ;
      LAYER met2 ;
        RECT 550.610 400.250 550.890 404.000 ;
        RECT 549.400 400.110 550.890 400.250 ;
        RECT 549.400 376.030 549.540 400.110 ;
        RECT 550.610 400.000 550.890 400.110 ;
        RECT 545.660 375.710 545.920 376.030 ;
        RECT 549.340 375.710 549.600 376.030 ;
        RECT 545.720 30.590 545.860 375.710 ;
        RECT 545.660 30.270 545.920 30.590 ;
        RECT 1161.140 30.270 1161.400 30.590 ;
        RECT 1161.200 2.400 1161.340 30.270 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 375.940 552.390 376.000 ;
        RECT 554.370 375.940 554.690 376.000 ;
        RECT 552.070 375.800 554.690 375.940 ;
        RECT 552.070 375.740 552.390 375.800 ;
        RECT 554.370 375.740 554.690 375.800 ;
        RECT 552.070 34.240 552.390 34.300 ;
        RECT 1179.050 34.240 1179.370 34.300 ;
        RECT 552.070 34.100 1179.370 34.240 ;
        RECT 552.070 34.040 552.390 34.100 ;
        RECT 1179.050 34.040 1179.370 34.100 ;
      LAYER via ;
        RECT 552.100 375.740 552.360 376.000 ;
        RECT 554.400 375.740 554.660 376.000 ;
        RECT 552.100 34.040 552.360 34.300 ;
        RECT 1179.080 34.040 1179.340 34.300 ;
      LAYER met2 ;
        RECT 555.670 400.250 555.950 404.000 ;
        RECT 554.460 400.110 555.950 400.250 ;
        RECT 554.460 376.030 554.600 400.110 ;
        RECT 555.670 400.000 555.950 400.110 ;
        RECT 552.100 375.710 552.360 376.030 ;
        RECT 554.400 375.710 554.660 376.030 ;
        RECT 552.160 34.330 552.300 375.710 ;
        RECT 552.100 34.010 552.360 34.330 ;
        RECT 1179.080 34.010 1179.340 34.330 ;
        RECT 1179.140 2.400 1179.280 34.010 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 378.320 559.290 378.380 ;
        RECT 559.890 378.320 560.210 378.380 ;
        RECT 558.970 378.180 560.210 378.320 ;
        RECT 558.970 378.120 559.290 378.180 ;
        RECT 559.890 378.120 560.210 378.180 ;
        RECT 558.970 33.900 559.290 33.960 ;
        RECT 1196.530 33.900 1196.850 33.960 ;
        RECT 558.970 33.760 1196.850 33.900 ;
        RECT 558.970 33.700 559.290 33.760 ;
        RECT 1196.530 33.700 1196.850 33.760 ;
      LAYER via ;
        RECT 559.000 378.120 559.260 378.380 ;
        RECT 559.920 378.120 560.180 378.380 ;
        RECT 559.000 33.700 559.260 33.960 ;
        RECT 1196.560 33.700 1196.820 33.960 ;
      LAYER met2 ;
        RECT 561.190 400.250 561.470 404.000 ;
        RECT 559.980 400.110 561.470 400.250 ;
        RECT 559.980 378.410 560.120 400.110 ;
        RECT 561.190 400.000 561.470 400.110 ;
        RECT 559.000 378.090 559.260 378.410 ;
        RECT 559.920 378.090 560.180 378.410 ;
        RECT 559.060 33.990 559.200 378.090 ;
        RECT 559.000 33.670 559.260 33.990 ;
        RECT 1196.560 33.670 1196.820 33.990 ;
        RECT 1196.620 2.400 1196.760 33.670 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.330 33.560 566.650 33.620 ;
        RECT 1214.930 33.560 1215.250 33.620 ;
        RECT 566.330 33.420 1215.250 33.560 ;
        RECT 566.330 33.360 566.650 33.420 ;
        RECT 1214.930 33.360 1215.250 33.420 ;
      LAYER via ;
        RECT 566.360 33.360 566.620 33.620 ;
        RECT 1214.960 33.360 1215.220 33.620 ;
      LAYER met2 ;
        RECT 566.710 400.250 566.990 404.000 ;
        RECT 566.420 400.110 566.990 400.250 ;
        RECT 566.420 33.650 566.560 400.110 ;
        RECT 566.710 400.000 566.990 400.110 ;
        RECT 566.360 33.330 566.620 33.650 ;
        RECT 1214.960 33.330 1215.220 33.650 ;
        RECT 1215.020 14.690 1215.160 33.330 ;
        RECT 1214.560 14.550 1215.160 14.690 ;
        RECT 1214.560 2.400 1214.700 14.550 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 376.280 566.190 376.340 ;
        RECT 570.470 376.280 570.790 376.340 ;
        RECT 565.870 376.140 570.790 376.280 ;
        RECT 565.870 376.080 566.190 376.140 ;
        RECT 570.470 376.080 570.790 376.140 ;
        RECT 565.870 33.220 566.190 33.280 ;
        RECT 1231.950 33.220 1232.270 33.280 ;
        RECT 565.870 33.080 1232.270 33.220 ;
        RECT 565.870 33.020 566.190 33.080 ;
        RECT 1231.950 33.020 1232.270 33.080 ;
      LAYER via ;
        RECT 565.900 376.080 566.160 376.340 ;
        RECT 570.500 376.080 570.760 376.340 ;
        RECT 565.900 33.020 566.160 33.280 ;
        RECT 1231.980 33.020 1232.240 33.280 ;
      LAYER met2 ;
        RECT 571.770 400.250 572.050 404.000 ;
        RECT 570.560 400.110 572.050 400.250 ;
        RECT 570.560 376.370 570.700 400.110 ;
        RECT 571.770 400.000 572.050 400.110 ;
        RECT 565.900 376.050 566.160 376.370 ;
        RECT 570.500 376.050 570.760 376.370 ;
        RECT 565.960 33.310 566.100 376.050 ;
        RECT 565.900 32.990 566.160 33.310 ;
        RECT 1231.980 32.990 1232.240 33.310 ;
        RECT 1232.040 2.400 1232.180 32.990 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 375.940 573.090 376.000 ;
        RECT 575.990 375.940 576.310 376.000 ;
        RECT 572.770 375.800 576.310 375.940 ;
        RECT 572.770 375.740 573.090 375.800 ;
        RECT 575.990 375.740 576.310 375.800 ;
        RECT 572.770 32.880 573.090 32.940 ;
        RECT 1249.890 32.880 1250.210 32.940 ;
        RECT 572.770 32.740 1250.210 32.880 ;
        RECT 572.770 32.680 573.090 32.740 ;
        RECT 1249.890 32.680 1250.210 32.740 ;
      LAYER via ;
        RECT 572.800 375.740 573.060 376.000 ;
        RECT 576.020 375.740 576.280 376.000 ;
        RECT 572.800 32.680 573.060 32.940 ;
        RECT 1249.920 32.680 1250.180 32.940 ;
      LAYER met2 ;
        RECT 577.290 400.250 577.570 404.000 ;
        RECT 576.080 400.110 577.570 400.250 ;
        RECT 576.080 376.030 576.220 400.110 ;
        RECT 577.290 400.000 577.570 400.110 ;
        RECT 572.800 375.710 573.060 376.030 ;
        RECT 576.020 375.710 576.280 376.030 ;
        RECT 572.860 32.970 573.000 375.710 ;
        RECT 572.800 32.650 573.060 32.970 ;
        RECT 1249.920 32.650 1250.180 32.970 ;
        RECT 1249.980 2.400 1250.120 32.650 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.670 376.280 579.990 376.340 ;
        RECT 581.510 376.280 581.830 376.340 ;
        RECT 579.670 376.140 581.830 376.280 ;
        RECT 579.670 376.080 579.990 376.140 ;
        RECT 581.510 376.080 581.830 376.140 ;
        RECT 579.670 32.540 579.990 32.600 ;
        RECT 1267.370 32.540 1267.690 32.600 ;
        RECT 579.670 32.400 1267.690 32.540 ;
        RECT 579.670 32.340 579.990 32.400 ;
        RECT 1267.370 32.340 1267.690 32.400 ;
      LAYER via ;
        RECT 579.700 376.080 579.960 376.340 ;
        RECT 581.540 376.080 581.800 376.340 ;
        RECT 579.700 32.340 579.960 32.600 ;
        RECT 1267.400 32.340 1267.660 32.600 ;
      LAYER met2 ;
        RECT 582.350 400.250 582.630 404.000 ;
        RECT 581.600 400.110 582.630 400.250 ;
        RECT 581.600 376.370 581.740 400.110 ;
        RECT 582.350 400.000 582.630 400.110 ;
        RECT 579.700 376.050 579.960 376.370 ;
        RECT 581.540 376.050 581.800 376.370 ;
        RECT 579.760 32.630 579.900 376.050 ;
        RECT 579.700 32.310 579.960 32.630 ;
        RECT 1267.400 32.310 1267.660 32.630 ;
        RECT 1267.460 2.400 1267.600 32.310 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 32.200 586.890 32.260 ;
        RECT 1285.310 32.200 1285.630 32.260 ;
        RECT 586.570 32.060 1285.630 32.200 ;
        RECT 586.570 32.000 586.890 32.060 ;
        RECT 1285.310 32.000 1285.630 32.060 ;
      LAYER via ;
        RECT 586.600 32.000 586.860 32.260 ;
        RECT 1285.340 32.000 1285.600 32.260 ;
      LAYER met2 ;
        RECT 587.870 400.250 588.150 404.000 ;
        RECT 586.660 400.110 588.150 400.250 ;
        RECT 586.660 32.290 586.800 400.110 ;
        RECT 587.870 400.000 588.150 400.110 ;
        RECT 586.600 31.970 586.860 32.290 ;
        RECT 1285.340 31.970 1285.600 32.290 ;
        RECT 1285.400 2.400 1285.540 31.970 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 376.280 593.790 376.340 ;
        RECT 594.390 376.280 594.710 376.340 ;
        RECT 593.470 376.140 594.710 376.280 ;
        RECT 593.470 376.080 593.790 376.140 ;
        RECT 594.390 376.080 594.710 376.140 ;
      LAYER via ;
        RECT 593.500 376.080 593.760 376.340 ;
        RECT 594.420 376.080 594.680 376.340 ;
      LAYER met2 ;
        RECT 593.390 400.180 593.670 404.000 ;
        RECT 593.390 400.000 593.700 400.180 ;
        RECT 593.560 376.370 593.700 400.000 ;
        RECT 593.500 376.050 593.760 376.370 ;
        RECT 594.420 376.050 594.680 376.370 ;
        RECT 594.480 31.805 594.620 376.050 ;
        RECT 594.410 31.435 594.690 31.805 ;
        RECT 1303.270 31.435 1303.550 31.805 ;
        RECT 1303.340 2.400 1303.480 31.435 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
      LAYER via2 ;
        RECT 594.410 31.480 594.690 31.760 ;
        RECT 1303.270 31.480 1303.550 31.760 ;
      LAYER met3 ;
        RECT 594.385 31.770 594.715 31.785 ;
        RECT 1303.245 31.770 1303.575 31.785 ;
        RECT 594.385 31.470 1303.575 31.770 ;
        RECT 594.385 31.455 594.715 31.470 ;
        RECT 1303.245 31.455 1303.575 31.470 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 375.600 593.790 375.660 ;
        RECT 597.610 375.600 597.930 375.660 ;
        RECT 593.470 375.460 597.930 375.600 ;
        RECT 593.470 375.400 593.790 375.460 ;
        RECT 597.610 375.400 597.930 375.460 ;
      LAYER via ;
        RECT 593.500 375.400 593.760 375.660 ;
        RECT 597.640 375.400 597.900 375.660 ;
      LAYER met2 ;
        RECT 598.450 400.250 598.730 404.000 ;
        RECT 597.700 400.110 598.730 400.250 ;
        RECT 597.700 375.690 597.840 400.110 ;
        RECT 598.450 400.000 598.730 400.110 ;
        RECT 593.500 375.370 593.760 375.690 ;
        RECT 597.640 375.370 597.900 375.690 ;
        RECT 593.560 31.125 593.700 375.370 ;
        RECT 593.490 30.755 593.770 31.125 ;
        RECT 1320.750 30.755 1321.030 31.125 ;
        RECT 1320.820 2.400 1320.960 30.755 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
      LAYER via2 ;
        RECT 593.490 30.800 593.770 31.080 ;
        RECT 1320.750 30.800 1321.030 31.080 ;
      LAYER met3 ;
        RECT 593.465 31.090 593.795 31.105 ;
        RECT 1320.725 31.090 1321.055 31.105 ;
        RECT 593.465 30.790 1321.055 31.090 ;
        RECT 593.465 30.775 593.795 30.790 ;
        RECT 1320.725 30.775 1321.055 30.790 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 386.480 400.590 386.540 ;
        RECT 404.410 386.480 404.730 386.540 ;
        RECT 400.270 386.340 404.730 386.480 ;
        RECT 400.270 386.280 400.590 386.340 ;
        RECT 404.410 386.280 404.730 386.340 ;
        RECT 400.270 22.680 400.590 22.740 ;
        RECT 682.250 22.680 682.570 22.740 ;
        RECT 400.270 22.540 682.570 22.680 ;
        RECT 400.270 22.480 400.590 22.540 ;
        RECT 682.250 22.480 682.570 22.540 ;
      LAYER via ;
        RECT 400.300 386.280 400.560 386.540 ;
        RECT 404.440 386.280 404.700 386.540 ;
        RECT 400.300 22.480 400.560 22.740 ;
        RECT 682.280 22.480 682.540 22.740 ;
      LAYER met2 ;
        RECT 405.710 400.250 405.990 404.000 ;
        RECT 404.500 400.110 405.990 400.250 ;
        RECT 404.500 386.570 404.640 400.110 ;
        RECT 405.710 400.000 405.990 400.110 ;
        RECT 400.300 386.250 400.560 386.570 ;
        RECT 404.440 386.250 404.700 386.570 ;
        RECT 400.360 22.770 400.500 386.250 ;
        RECT 400.300 22.450 400.560 22.770 ;
        RECT 682.280 22.450 682.540 22.770 ;
        RECT 682.340 2.400 682.480 22.450 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 105.640 602.070 105.700 ;
        RECT 1338.670 105.640 1338.990 105.700 ;
        RECT 601.750 105.500 1338.990 105.640 ;
        RECT 601.750 105.440 602.070 105.500 ;
        RECT 1338.670 105.440 1338.990 105.500 ;
      LAYER via ;
        RECT 601.780 105.440 602.040 105.700 ;
        RECT 1338.700 105.440 1338.960 105.700 ;
      LAYER met2 ;
        RECT 603.970 400.250 604.250 404.000 ;
        RECT 602.760 400.110 604.250 400.250 ;
        RECT 602.760 324.370 602.900 400.110 ;
        RECT 603.970 400.000 604.250 400.110 ;
        RECT 601.840 324.230 602.900 324.370 ;
        RECT 601.840 105.730 601.980 324.230 ;
        RECT 601.780 105.410 602.040 105.730 ;
        RECT 1338.700 105.410 1338.960 105.730 ;
        RECT 1338.760 2.400 1338.900 105.410 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.650 105.980 608.970 106.040 ;
        RECT 1352.470 105.980 1352.790 106.040 ;
        RECT 608.650 105.840 1352.790 105.980 ;
        RECT 608.650 105.780 608.970 105.840 ;
        RECT 1352.470 105.780 1352.790 105.840 ;
      LAYER via ;
        RECT 608.680 105.780 608.940 106.040 ;
        RECT 1352.500 105.780 1352.760 106.040 ;
      LAYER met2 ;
        RECT 609.490 400.250 609.770 404.000 ;
        RECT 608.740 400.110 609.770 400.250 ;
        RECT 608.740 106.070 608.880 400.110 ;
        RECT 609.490 400.000 609.770 400.110 ;
        RECT 608.680 105.750 608.940 106.070 ;
        RECT 1352.500 105.750 1352.760 106.070 ;
        RECT 1352.560 82.870 1352.700 105.750 ;
        RECT 1352.560 82.730 1354.080 82.870 ;
        RECT 1353.940 1.770 1354.080 82.730 ;
        RECT 1356.030 1.770 1356.590 2.400 ;
        RECT 1353.940 1.630 1356.590 1.770 ;
        RECT 1356.030 -4.800 1356.590 1.630 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.550 106.320 615.870 106.380 ;
        RECT 1373.170 106.320 1373.490 106.380 ;
        RECT 615.550 106.180 1373.490 106.320 ;
        RECT 615.550 106.120 615.870 106.180 ;
        RECT 1373.170 106.120 1373.490 106.180 ;
      LAYER via ;
        RECT 615.580 106.120 615.840 106.380 ;
        RECT 1373.200 106.120 1373.460 106.380 ;
      LAYER met2 ;
        RECT 614.550 400.250 614.830 404.000 ;
        RECT 614.550 400.110 616.240 400.250 ;
        RECT 614.550 400.000 614.830 400.110 ;
        RECT 616.100 351.970 616.240 400.110 ;
        RECT 616.100 351.830 616.700 351.970 ;
        RECT 616.560 324.370 616.700 351.830 ;
        RECT 615.640 324.230 616.700 324.370 ;
        RECT 615.640 106.410 615.780 324.230 ;
        RECT 615.580 106.090 615.840 106.410 ;
        RECT 1373.200 106.090 1373.460 106.410 ;
        RECT 1373.260 82.870 1373.400 106.090 ;
        RECT 1373.260 82.730 1374.320 82.870 ;
        RECT 1374.180 2.400 1374.320 82.730 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 376.280 615.410 376.340 ;
        RECT 618.770 376.280 619.090 376.340 ;
        RECT 615.090 376.140 619.090 376.280 ;
        RECT 615.090 376.080 615.410 376.140 ;
        RECT 618.770 376.080 619.090 376.140 ;
        RECT 615.090 106.660 615.410 106.720 ;
        RECT 1386.970 106.660 1387.290 106.720 ;
        RECT 615.090 106.520 1387.290 106.660 ;
        RECT 615.090 106.460 615.410 106.520 ;
        RECT 1386.970 106.460 1387.290 106.520 ;
      LAYER via ;
        RECT 615.120 376.080 615.380 376.340 ;
        RECT 618.800 376.080 619.060 376.340 ;
        RECT 615.120 106.460 615.380 106.720 ;
        RECT 1387.000 106.460 1387.260 106.720 ;
      LAYER met2 ;
        RECT 620.070 400.250 620.350 404.000 ;
        RECT 618.860 400.110 620.350 400.250 ;
        RECT 618.860 376.370 619.000 400.110 ;
        RECT 620.070 400.000 620.350 400.110 ;
        RECT 615.120 376.050 615.380 376.370 ;
        RECT 618.800 376.050 619.060 376.370 ;
        RECT 615.180 106.750 615.320 376.050 ;
        RECT 615.120 106.430 615.380 106.750 ;
        RECT 1387.000 106.430 1387.260 106.750 ;
        RECT 1387.060 82.870 1387.200 106.430 ;
        RECT 1387.060 82.730 1391.800 82.870 ;
        RECT 1391.660 2.400 1391.800 82.730 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 110.400 622.770 110.460 ;
        RECT 1407.670 110.400 1407.990 110.460 ;
        RECT 622.450 110.260 1407.990 110.400 ;
        RECT 622.450 110.200 622.770 110.260 ;
        RECT 1407.670 110.200 1407.990 110.260 ;
      LAYER via ;
        RECT 622.480 110.200 622.740 110.460 ;
        RECT 1407.700 110.200 1407.960 110.460 ;
      LAYER met2 ;
        RECT 625.590 400.250 625.870 404.000 ;
        RECT 624.380 400.110 625.870 400.250 ;
        RECT 624.380 324.370 624.520 400.110 ;
        RECT 625.590 400.000 625.870 400.110 ;
        RECT 622.540 324.230 624.520 324.370 ;
        RECT 622.540 110.490 622.680 324.230 ;
        RECT 622.480 110.170 622.740 110.490 ;
        RECT 1407.700 110.170 1407.960 110.490 ;
        RECT 1407.760 1.770 1407.900 110.170 ;
        RECT 1409.390 1.770 1409.950 2.400 ;
        RECT 1407.760 1.630 1409.950 1.770 ;
        RECT 1409.390 -4.800 1409.950 1.630 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.970 376.280 628.290 376.340 ;
        RECT 629.810 376.280 630.130 376.340 ;
        RECT 627.970 376.140 630.130 376.280 ;
        RECT 627.970 376.080 628.290 376.140 ;
        RECT 629.810 376.080 630.130 376.140 ;
        RECT 627.970 36.280 628.290 36.340 ;
        RECT 1426.990 36.280 1427.310 36.340 ;
        RECT 627.970 36.140 1427.310 36.280 ;
        RECT 627.970 36.080 628.290 36.140 ;
        RECT 1426.990 36.080 1427.310 36.140 ;
      LAYER via ;
        RECT 628.000 376.080 628.260 376.340 ;
        RECT 629.840 376.080 630.100 376.340 ;
        RECT 628.000 36.080 628.260 36.340 ;
        RECT 1427.020 36.080 1427.280 36.340 ;
      LAYER met2 ;
        RECT 630.650 400.250 630.930 404.000 ;
        RECT 629.900 400.110 630.930 400.250 ;
        RECT 629.900 376.370 630.040 400.110 ;
        RECT 630.650 400.000 630.930 400.110 ;
        RECT 628.000 376.050 628.260 376.370 ;
        RECT 629.840 376.050 630.100 376.370 ;
        RECT 628.060 36.370 628.200 376.050 ;
        RECT 628.000 36.050 628.260 36.370 ;
        RECT 1427.020 36.050 1427.280 36.370 ;
        RECT 1427.080 2.400 1427.220 36.050 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.870 36.620 635.190 36.680 ;
        RECT 1444.930 36.620 1445.250 36.680 ;
        RECT 634.870 36.480 1445.250 36.620 ;
        RECT 634.870 36.420 635.190 36.480 ;
        RECT 1444.930 36.420 1445.250 36.480 ;
      LAYER via ;
        RECT 634.900 36.420 635.160 36.680 ;
        RECT 1444.960 36.420 1445.220 36.680 ;
      LAYER met2 ;
        RECT 636.170 400.250 636.450 404.000 ;
        RECT 634.960 400.110 636.450 400.250 ;
        RECT 634.960 36.710 635.100 400.110 ;
        RECT 636.170 400.000 636.450 400.110 ;
        RECT 634.900 36.390 635.160 36.710 ;
        RECT 1444.960 36.390 1445.220 36.710 ;
        RECT 1445.020 2.400 1445.160 36.390 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.230 36.960 642.550 37.020 ;
        RECT 1462.870 36.960 1463.190 37.020 ;
        RECT 642.230 36.820 1463.190 36.960 ;
        RECT 642.230 36.760 642.550 36.820 ;
        RECT 1462.870 36.760 1463.190 36.820 ;
      LAYER via ;
        RECT 642.260 36.760 642.520 37.020 ;
        RECT 1462.900 36.760 1463.160 37.020 ;
      LAYER met2 ;
        RECT 641.690 400.250 641.970 404.000 ;
        RECT 641.690 400.110 642.460 400.250 ;
        RECT 641.690 400.000 641.970 400.110 ;
        RECT 642.320 37.050 642.460 400.110 ;
        RECT 642.260 36.730 642.520 37.050 ;
        RECT 1462.900 36.730 1463.160 37.050 ;
        RECT 1462.960 2.400 1463.100 36.730 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 376.280 642.090 376.340 ;
        RECT 645.450 376.280 645.770 376.340 ;
        RECT 641.770 376.140 645.770 376.280 ;
        RECT 641.770 376.080 642.090 376.140 ;
        RECT 645.450 376.080 645.770 376.140 ;
        RECT 641.770 37.300 642.090 37.360 ;
        RECT 1480.350 37.300 1480.670 37.360 ;
        RECT 641.770 37.160 1480.670 37.300 ;
        RECT 641.770 37.100 642.090 37.160 ;
        RECT 1480.350 37.100 1480.670 37.160 ;
      LAYER via ;
        RECT 641.800 376.080 642.060 376.340 ;
        RECT 645.480 376.080 645.740 376.340 ;
        RECT 641.800 37.100 642.060 37.360 ;
        RECT 1480.380 37.100 1480.640 37.360 ;
      LAYER met2 ;
        RECT 646.750 400.250 647.030 404.000 ;
        RECT 645.540 400.110 647.030 400.250 ;
        RECT 645.540 376.370 645.680 400.110 ;
        RECT 646.750 400.000 647.030 400.110 ;
        RECT 641.800 376.050 642.060 376.370 ;
        RECT 645.480 376.050 645.740 376.370 ;
        RECT 641.860 37.390 642.000 376.050 ;
        RECT 641.800 37.070 642.060 37.390 ;
        RECT 1480.380 37.070 1480.640 37.390 ;
        RECT 1480.440 2.400 1480.580 37.070 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 375.600 648.990 375.660 ;
        RECT 650.970 375.600 651.290 375.660 ;
        RECT 648.670 375.460 651.290 375.600 ;
        RECT 648.670 375.400 648.990 375.460 ;
        RECT 650.970 375.400 651.290 375.460 ;
        RECT 648.670 37.640 648.990 37.700 ;
        RECT 1498.290 37.640 1498.610 37.700 ;
        RECT 648.670 37.500 1498.610 37.640 ;
        RECT 648.670 37.440 648.990 37.500 ;
        RECT 1498.290 37.440 1498.610 37.500 ;
      LAYER via ;
        RECT 648.700 375.400 648.960 375.660 ;
        RECT 651.000 375.400 651.260 375.660 ;
        RECT 648.700 37.440 648.960 37.700 ;
        RECT 1498.320 37.440 1498.580 37.700 ;
      LAYER met2 ;
        RECT 652.270 400.250 652.550 404.000 ;
        RECT 651.060 400.110 652.550 400.250 ;
        RECT 651.060 375.690 651.200 400.110 ;
        RECT 652.270 400.000 652.550 400.110 ;
        RECT 648.700 375.370 648.960 375.690 ;
        RECT 651.000 375.370 651.260 375.690 ;
        RECT 648.760 37.730 648.900 375.370 ;
        RECT 648.700 37.410 648.960 37.730 ;
        RECT 1498.320 37.410 1498.580 37.730 ;
        RECT 1498.380 2.400 1498.520 37.410 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 375.940 407.490 376.000 ;
        RECT 409.930 375.940 410.250 376.000 ;
        RECT 407.170 375.800 410.250 375.940 ;
        RECT 407.170 375.740 407.490 375.800 ;
        RECT 409.930 375.740 410.250 375.800 ;
        RECT 407.170 23.700 407.490 23.760 ;
        RECT 700.190 23.700 700.510 23.760 ;
        RECT 407.170 23.560 700.510 23.700 ;
        RECT 407.170 23.500 407.490 23.560 ;
        RECT 700.190 23.500 700.510 23.560 ;
      LAYER via ;
        RECT 407.200 375.740 407.460 376.000 ;
        RECT 409.960 375.740 410.220 376.000 ;
        RECT 407.200 23.500 407.460 23.760 ;
        RECT 700.220 23.500 700.480 23.760 ;
      LAYER met2 ;
        RECT 411.230 400.250 411.510 404.000 ;
        RECT 410.020 400.110 411.510 400.250 ;
        RECT 410.020 376.030 410.160 400.110 ;
        RECT 411.230 400.000 411.510 400.110 ;
        RECT 407.200 375.710 407.460 376.030 ;
        RECT 409.960 375.710 410.220 376.030 ;
        RECT 407.260 23.790 407.400 375.710 ;
        RECT 407.200 23.470 407.460 23.790 ;
        RECT 700.220 23.470 700.480 23.790 ;
        RECT 700.280 2.400 700.420 23.470 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 655.570 399.740 655.890 399.800 ;
        RECT 656.490 399.740 656.810 399.800 ;
        RECT 655.570 399.600 656.810 399.740 ;
        RECT 655.570 399.540 655.890 399.600 ;
        RECT 656.490 399.540 656.810 399.600 ;
        RECT 655.570 41.380 655.890 41.440 ;
        RECT 1515.770 41.380 1516.090 41.440 ;
        RECT 655.570 41.240 1516.090 41.380 ;
        RECT 655.570 41.180 655.890 41.240 ;
        RECT 1515.770 41.180 1516.090 41.240 ;
      LAYER via ;
        RECT 655.600 399.540 655.860 399.800 ;
        RECT 656.520 399.540 656.780 399.800 ;
        RECT 655.600 41.180 655.860 41.440 ;
        RECT 1515.800 41.180 1516.060 41.440 ;
      LAYER met2 ;
        RECT 657.790 400.250 658.070 404.000 ;
        RECT 656.580 400.110 658.070 400.250 ;
        RECT 656.580 399.830 656.720 400.110 ;
        RECT 657.790 400.000 658.070 400.110 ;
        RECT 655.600 399.510 655.860 399.830 ;
        RECT 656.520 399.510 656.780 399.830 ;
        RECT 655.660 41.470 655.800 399.510 ;
        RECT 655.600 41.150 655.860 41.470 ;
        RECT 1515.800 41.150 1516.060 41.470 ;
        RECT 1515.860 2.400 1516.000 41.150 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 41.040 662.790 41.100 ;
        RECT 1533.710 41.040 1534.030 41.100 ;
        RECT 662.470 40.900 1534.030 41.040 ;
        RECT 662.470 40.840 662.790 40.900 ;
        RECT 1533.710 40.840 1534.030 40.900 ;
      LAYER via ;
        RECT 662.500 40.840 662.760 41.100 ;
        RECT 1533.740 40.840 1534.000 41.100 ;
      LAYER met2 ;
        RECT 662.850 400.250 663.130 404.000 ;
        RECT 662.560 400.110 663.130 400.250 ;
        RECT 662.560 41.130 662.700 400.110 ;
        RECT 662.850 400.000 663.130 400.110 ;
        RECT 662.500 40.810 662.760 41.130 ;
        RECT 1533.740 40.810 1534.000 41.130 ;
        RECT 1533.800 2.400 1533.940 40.810 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.930 376.280 663.250 376.340 ;
        RECT 667.070 376.280 667.390 376.340 ;
        RECT 662.930 376.140 667.390 376.280 ;
        RECT 662.930 376.080 663.250 376.140 ;
        RECT 667.070 376.080 667.390 376.140 ;
        RECT 662.930 40.700 663.250 40.760 ;
        RECT 1551.190 40.700 1551.510 40.760 ;
        RECT 662.930 40.560 1551.510 40.700 ;
        RECT 662.930 40.500 663.250 40.560 ;
        RECT 1551.190 40.500 1551.510 40.560 ;
      LAYER via ;
        RECT 662.960 376.080 663.220 376.340 ;
        RECT 667.100 376.080 667.360 376.340 ;
        RECT 662.960 40.500 663.220 40.760 ;
        RECT 1551.220 40.500 1551.480 40.760 ;
      LAYER met2 ;
        RECT 668.370 400.250 668.650 404.000 ;
        RECT 667.160 400.110 668.650 400.250 ;
        RECT 667.160 376.370 667.300 400.110 ;
        RECT 668.370 400.000 668.650 400.110 ;
        RECT 662.960 376.050 663.220 376.370 ;
        RECT 667.100 376.050 667.360 376.370 ;
        RECT 663.020 40.790 663.160 376.050 ;
        RECT 662.960 40.470 663.220 40.790 ;
        RECT 1551.220 40.470 1551.480 40.790 ;
        RECT 1551.280 2.400 1551.420 40.470 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.370 375.940 669.690 376.000 ;
        RECT 672.590 375.940 672.910 376.000 ;
        RECT 669.370 375.800 672.910 375.940 ;
        RECT 669.370 375.740 669.690 375.800 ;
        RECT 672.590 375.740 672.910 375.800 ;
        RECT 669.370 40.360 669.690 40.420 ;
        RECT 1569.130 40.360 1569.450 40.420 ;
        RECT 669.370 40.220 1569.450 40.360 ;
        RECT 669.370 40.160 669.690 40.220 ;
        RECT 1569.130 40.160 1569.450 40.220 ;
      LAYER via ;
        RECT 669.400 375.740 669.660 376.000 ;
        RECT 672.620 375.740 672.880 376.000 ;
        RECT 669.400 40.160 669.660 40.420 ;
        RECT 1569.160 40.160 1569.420 40.420 ;
      LAYER met2 ;
        RECT 673.430 400.250 673.710 404.000 ;
        RECT 672.680 400.110 673.710 400.250 ;
        RECT 672.680 376.030 672.820 400.110 ;
        RECT 673.430 400.000 673.710 400.110 ;
        RECT 669.400 375.710 669.660 376.030 ;
        RECT 672.620 375.710 672.880 376.030 ;
        RECT 669.460 40.450 669.600 375.710 ;
        RECT 669.400 40.130 669.660 40.450 ;
        RECT 1569.160 40.130 1569.420 40.450 ;
        RECT 1569.220 2.400 1569.360 40.130 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.270 376.280 676.590 376.340 ;
        RECT 677.650 376.280 677.970 376.340 ;
        RECT 676.270 376.140 677.970 376.280 ;
        RECT 676.270 376.080 676.590 376.140 ;
        RECT 677.650 376.080 677.970 376.140 ;
        RECT 676.270 40.020 676.590 40.080 ;
        RECT 1586.610 40.020 1586.930 40.080 ;
        RECT 676.270 39.880 1586.930 40.020 ;
        RECT 676.270 39.820 676.590 39.880 ;
        RECT 1586.610 39.820 1586.930 39.880 ;
      LAYER via ;
        RECT 676.300 376.080 676.560 376.340 ;
        RECT 677.680 376.080 677.940 376.340 ;
        RECT 676.300 39.820 676.560 40.080 ;
        RECT 1586.640 39.820 1586.900 40.080 ;
      LAYER met2 ;
        RECT 678.950 400.250 679.230 404.000 ;
        RECT 677.740 400.110 679.230 400.250 ;
        RECT 677.740 376.370 677.880 400.110 ;
        RECT 678.950 400.000 679.230 400.110 ;
        RECT 676.300 376.050 676.560 376.370 ;
        RECT 677.680 376.050 677.940 376.370 ;
        RECT 676.360 40.110 676.500 376.050 ;
        RECT 676.300 39.790 676.560 40.110 ;
        RECT 1586.640 39.790 1586.900 40.110 ;
        RECT 1586.700 2.400 1586.840 39.790 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.170 39.680 683.490 39.740 ;
        RECT 1604.550 39.680 1604.870 39.740 ;
        RECT 683.170 39.540 1604.870 39.680 ;
        RECT 683.170 39.480 683.490 39.540 ;
        RECT 1604.550 39.480 1604.870 39.540 ;
      LAYER via ;
        RECT 683.200 39.480 683.460 39.740 ;
        RECT 1604.580 39.480 1604.840 39.740 ;
      LAYER met2 ;
        RECT 684.470 400.250 684.750 404.000 ;
        RECT 683.260 400.110 684.750 400.250 ;
        RECT 683.260 39.770 683.400 400.110 ;
        RECT 684.470 400.000 684.750 400.110 ;
        RECT 683.200 39.450 683.460 39.770 ;
        RECT 1604.580 39.450 1604.840 39.770 ;
        RECT 1604.640 2.400 1604.780 39.450 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 376.280 683.950 376.340 ;
        RECT 688.690 376.280 689.010 376.340 ;
        RECT 683.630 376.140 689.010 376.280 ;
        RECT 683.630 376.080 683.950 376.140 ;
        RECT 688.690 376.080 689.010 376.140 ;
        RECT 683.630 39.340 683.950 39.400 ;
        RECT 1622.030 39.340 1622.350 39.400 ;
        RECT 683.630 39.200 1622.350 39.340 ;
        RECT 683.630 39.140 683.950 39.200 ;
        RECT 1622.030 39.140 1622.350 39.200 ;
      LAYER via ;
        RECT 683.660 376.080 683.920 376.340 ;
        RECT 688.720 376.080 688.980 376.340 ;
        RECT 683.660 39.140 683.920 39.400 ;
        RECT 1622.060 39.140 1622.320 39.400 ;
      LAYER met2 ;
        RECT 689.530 400.250 689.810 404.000 ;
        RECT 688.780 400.110 689.810 400.250 ;
        RECT 688.780 376.370 688.920 400.110 ;
        RECT 689.530 400.000 689.810 400.110 ;
        RECT 683.660 376.050 683.920 376.370 ;
        RECT 688.720 376.050 688.980 376.370 ;
        RECT 683.720 39.430 683.860 376.050 ;
        RECT 683.660 39.110 683.920 39.430 ;
        RECT 1622.060 39.110 1622.320 39.430 ;
        RECT 1622.120 2.400 1622.260 39.110 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.070 373.220 690.390 373.280 ;
        RECT 693.750 373.220 694.070 373.280 ;
        RECT 690.070 373.080 694.070 373.220 ;
        RECT 690.070 373.020 690.390 373.080 ;
        RECT 693.750 373.020 694.070 373.080 ;
        RECT 690.070 39.000 690.390 39.060 ;
        RECT 1639.970 39.000 1640.290 39.060 ;
        RECT 690.070 38.860 1640.290 39.000 ;
        RECT 690.070 38.800 690.390 38.860 ;
        RECT 1639.970 38.800 1640.290 38.860 ;
      LAYER via ;
        RECT 690.100 373.020 690.360 373.280 ;
        RECT 693.780 373.020 694.040 373.280 ;
        RECT 690.100 38.800 690.360 39.060 ;
        RECT 1640.000 38.800 1640.260 39.060 ;
      LAYER met2 ;
        RECT 695.050 400.250 695.330 404.000 ;
        RECT 693.840 400.110 695.330 400.250 ;
        RECT 693.840 373.310 693.980 400.110 ;
        RECT 695.050 400.000 695.330 400.110 ;
        RECT 690.100 372.990 690.360 373.310 ;
        RECT 693.780 372.990 694.040 373.310 ;
        RECT 690.160 39.090 690.300 372.990 ;
        RECT 690.100 38.770 690.360 39.090 ;
        RECT 1640.000 38.770 1640.260 39.090 ;
        RECT 1640.060 2.400 1640.200 38.770 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.970 386.140 697.290 386.200 ;
        RECT 699.270 386.140 699.590 386.200 ;
        RECT 696.970 386.000 699.590 386.140 ;
        RECT 696.970 385.940 697.290 386.000 ;
        RECT 699.270 385.940 699.590 386.000 ;
        RECT 696.970 38.660 697.290 38.720 ;
        RECT 1657.910 38.660 1658.230 38.720 ;
        RECT 696.970 38.520 1658.230 38.660 ;
        RECT 696.970 38.460 697.290 38.520 ;
        RECT 1657.910 38.460 1658.230 38.520 ;
      LAYER via ;
        RECT 697.000 385.940 697.260 386.200 ;
        RECT 699.300 385.940 699.560 386.200 ;
        RECT 697.000 38.460 697.260 38.720 ;
        RECT 1657.940 38.460 1658.200 38.720 ;
      LAYER met2 ;
        RECT 700.570 400.250 700.850 404.000 ;
        RECT 699.360 400.110 700.850 400.250 ;
        RECT 699.360 386.230 699.500 400.110 ;
        RECT 700.570 400.000 700.850 400.110 ;
        RECT 697.000 385.910 697.260 386.230 ;
        RECT 699.300 385.910 699.560 386.230 ;
        RECT 697.060 38.750 697.200 385.910 ;
        RECT 697.000 38.430 697.260 38.750 ;
        RECT 1657.940 38.430 1658.200 38.750 ;
        RECT 1658.000 2.400 1658.140 38.430 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.870 38.320 704.190 38.380 ;
        RECT 1675.390 38.320 1675.710 38.380 ;
        RECT 703.870 38.180 1675.710 38.320 ;
        RECT 703.870 38.120 704.190 38.180 ;
        RECT 1675.390 38.120 1675.710 38.180 ;
      LAYER via ;
        RECT 703.900 38.120 704.160 38.380 ;
        RECT 1675.420 38.120 1675.680 38.380 ;
      LAYER met2 ;
        RECT 705.630 400.250 705.910 404.000 ;
        RECT 704.420 400.110 705.910 400.250 ;
        RECT 704.420 386.470 704.560 400.110 ;
        RECT 705.630 400.000 705.910 400.110 ;
        RECT 703.960 386.330 704.560 386.470 ;
        RECT 703.960 38.410 704.100 386.330 ;
        RECT 703.900 38.090 704.160 38.410 ;
        RECT 1675.420 38.090 1675.680 38.410 ;
        RECT 1675.480 2.400 1675.620 38.090 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 387.160 414.390 387.220 ;
        RECT 414.990 387.160 415.310 387.220 ;
        RECT 414.070 387.020 415.310 387.160 ;
        RECT 414.070 386.960 414.390 387.020 ;
        RECT 414.990 386.960 415.310 387.020 ;
        RECT 414.070 27.440 414.390 27.500 ;
        RECT 717.670 27.440 717.990 27.500 ;
        RECT 414.070 27.300 717.990 27.440 ;
        RECT 414.070 27.240 414.390 27.300 ;
        RECT 717.670 27.240 717.990 27.300 ;
      LAYER via ;
        RECT 414.100 386.960 414.360 387.220 ;
        RECT 415.020 386.960 415.280 387.220 ;
        RECT 414.100 27.240 414.360 27.500 ;
        RECT 717.700 27.240 717.960 27.500 ;
      LAYER met2 ;
        RECT 416.290 400.250 416.570 404.000 ;
        RECT 415.080 400.110 416.570 400.250 ;
        RECT 415.080 387.250 415.220 400.110 ;
        RECT 416.290 400.000 416.570 400.110 ;
        RECT 414.100 386.930 414.360 387.250 ;
        RECT 415.020 386.930 415.280 387.250 ;
        RECT 414.160 27.530 414.300 386.930 ;
        RECT 414.100 27.210 414.360 27.530 ;
        RECT 717.700 27.210 717.960 27.530 ;
        RECT 717.760 2.400 717.900 27.210 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.230 37.980 711.550 38.040 ;
        RECT 1693.330 37.980 1693.650 38.040 ;
        RECT 711.230 37.840 1693.650 37.980 ;
        RECT 711.230 37.780 711.550 37.840 ;
        RECT 1693.330 37.780 1693.650 37.840 ;
      LAYER via ;
        RECT 711.260 37.780 711.520 38.040 ;
        RECT 1693.360 37.780 1693.620 38.040 ;
      LAYER met2 ;
        RECT 711.150 400.180 711.430 404.000 ;
        RECT 711.150 400.000 711.460 400.180 ;
        RECT 711.320 38.070 711.460 400.000 ;
        RECT 711.260 37.750 711.520 38.070 ;
        RECT 1693.360 37.750 1693.620 38.070 ;
        RECT 1693.420 2.400 1693.560 37.750 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 710.770 386.480 711.090 386.540 ;
        RECT 715.370 386.480 715.690 386.540 ;
        RECT 710.770 386.340 715.690 386.480 ;
        RECT 710.770 386.280 711.090 386.340 ;
        RECT 715.370 386.280 715.690 386.340 ;
      LAYER via ;
        RECT 710.800 386.280 711.060 386.540 ;
        RECT 715.400 386.280 715.660 386.540 ;
      LAYER met2 ;
        RECT 716.670 400.250 716.950 404.000 ;
        RECT 715.460 400.110 716.950 400.250 ;
        RECT 715.460 386.570 715.600 400.110 ;
        RECT 716.670 400.000 716.950 400.110 ;
        RECT 710.800 386.250 711.060 386.570 ;
        RECT 715.400 386.250 715.660 386.570 ;
        RECT 710.860 38.605 711.000 386.250 ;
        RECT 710.790 38.235 711.070 38.605 ;
        RECT 1710.830 38.235 1711.110 38.605 ;
        RECT 1710.900 2.400 1711.040 38.235 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
      LAYER via2 ;
        RECT 710.790 38.280 711.070 38.560 ;
        RECT 1710.830 38.280 1711.110 38.560 ;
      LAYER met3 ;
        RECT 710.765 38.570 711.095 38.585 ;
        RECT 1710.805 38.570 1711.135 38.585 ;
        RECT 710.765 38.270 1711.135 38.570 ;
        RECT 710.765 38.255 711.095 38.270 ;
        RECT 1710.805 38.255 1711.135 38.270 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.590 386.480 718.910 386.540 ;
        RECT 720.430 386.480 720.750 386.540 ;
        RECT 718.590 386.340 720.750 386.480 ;
        RECT 718.590 386.280 718.910 386.340 ;
        RECT 720.430 386.280 720.750 386.340 ;
        RECT 718.590 110.060 718.910 110.120 ;
        RECT 1725.070 110.060 1725.390 110.120 ;
        RECT 718.590 109.920 1725.390 110.060 ;
        RECT 718.590 109.860 718.910 109.920 ;
        RECT 1725.070 109.860 1725.390 109.920 ;
      LAYER via ;
        RECT 718.620 386.280 718.880 386.540 ;
        RECT 720.460 386.280 720.720 386.540 ;
        RECT 718.620 109.860 718.880 110.120 ;
        RECT 1725.100 109.860 1725.360 110.120 ;
      LAYER met2 ;
        RECT 721.730 400.250 722.010 404.000 ;
        RECT 720.520 400.110 722.010 400.250 ;
        RECT 720.520 386.570 720.660 400.110 ;
        RECT 721.730 400.000 722.010 400.110 ;
        RECT 718.620 386.250 718.880 386.570 ;
        RECT 720.460 386.250 720.720 386.570 ;
        RECT 718.680 110.150 718.820 386.250 ;
        RECT 718.620 109.830 718.880 110.150 ;
        RECT 1725.100 109.830 1725.360 110.150 ;
        RECT 1725.160 82.870 1725.300 109.830 ;
        RECT 1725.160 82.730 1726.680 82.870 ;
        RECT 1726.540 1.770 1726.680 82.730 ;
        RECT 1728.630 1.770 1729.190 2.400 ;
        RECT 1726.540 1.630 1729.190 1.770 ;
        RECT 1728.630 -4.800 1729.190 1.630 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.030 386.480 725.350 386.540 ;
        RECT 725.950 386.480 726.270 386.540 ;
        RECT 725.030 386.340 726.270 386.480 ;
        RECT 725.030 386.280 725.350 386.340 ;
        RECT 725.950 386.280 726.270 386.340 ;
        RECT 725.030 109.720 725.350 109.780 ;
        RECT 1745.770 109.720 1746.090 109.780 ;
        RECT 725.030 109.580 1746.090 109.720 ;
        RECT 725.030 109.520 725.350 109.580 ;
        RECT 1745.770 109.520 1746.090 109.580 ;
      LAYER via ;
        RECT 725.060 386.280 725.320 386.540 ;
        RECT 725.980 386.280 726.240 386.540 ;
        RECT 725.060 109.520 725.320 109.780 ;
        RECT 1745.800 109.520 1746.060 109.780 ;
      LAYER met2 ;
        RECT 727.250 400.250 727.530 404.000 ;
        RECT 726.040 400.110 727.530 400.250 ;
        RECT 726.040 386.570 726.180 400.110 ;
        RECT 727.250 400.000 727.530 400.110 ;
        RECT 725.060 386.250 725.320 386.570 ;
        RECT 725.980 386.250 726.240 386.570 ;
        RECT 725.120 109.810 725.260 386.250 ;
        RECT 725.060 109.490 725.320 109.810 ;
        RECT 1745.800 109.490 1746.060 109.810 ;
        RECT 1745.860 14.690 1746.000 109.490 ;
        RECT 1745.860 14.550 1746.460 14.690 ;
        RECT 1746.320 2.400 1746.460 14.550 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.930 116.520 732.250 116.580 ;
        RECT 1759.570 116.520 1759.890 116.580 ;
        RECT 731.930 116.380 1759.890 116.520 ;
        RECT 731.930 116.320 732.250 116.380 ;
        RECT 1759.570 116.320 1759.890 116.380 ;
      LAYER via ;
        RECT 731.960 116.320 732.220 116.580 ;
        RECT 1759.600 116.320 1759.860 116.580 ;
      LAYER met2 ;
        RECT 732.770 400.250 733.050 404.000 ;
        RECT 732.020 400.110 733.050 400.250 ;
        RECT 732.020 116.610 732.160 400.110 ;
        RECT 732.770 400.000 733.050 400.110 ;
        RECT 731.960 116.290 732.220 116.610 ;
        RECT 1759.600 116.290 1759.860 116.610 ;
        RECT 1759.660 82.870 1759.800 116.290 ;
        RECT 1759.660 82.730 1764.400 82.870 ;
        RECT 1764.260 2.400 1764.400 82.730 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.390 386.140 732.710 386.200 ;
        RECT 736.530 386.140 736.850 386.200 ;
        RECT 732.390 386.000 736.850 386.140 ;
        RECT 732.390 385.940 732.710 386.000 ;
        RECT 736.530 385.940 736.850 386.000 ;
        RECT 732.390 116.180 732.710 116.240 ;
        RECT 1780.270 116.180 1780.590 116.240 ;
        RECT 732.390 116.040 1780.590 116.180 ;
        RECT 732.390 115.980 732.710 116.040 ;
        RECT 1780.270 115.980 1780.590 116.040 ;
      LAYER via ;
        RECT 732.420 385.940 732.680 386.200 ;
        RECT 736.560 385.940 736.820 386.200 ;
        RECT 732.420 115.980 732.680 116.240 ;
        RECT 1780.300 115.980 1780.560 116.240 ;
      LAYER met2 ;
        RECT 737.830 400.250 738.110 404.000 ;
        RECT 736.620 400.110 738.110 400.250 ;
        RECT 736.620 386.230 736.760 400.110 ;
        RECT 737.830 400.000 738.110 400.110 ;
        RECT 732.420 385.910 732.680 386.230 ;
        RECT 736.560 385.910 736.820 386.230 ;
        RECT 732.480 116.270 732.620 385.910 ;
        RECT 732.420 115.950 732.680 116.270 ;
        RECT 1780.300 115.950 1780.560 116.270 ;
        RECT 1780.360 82.870 1780.500 115.950 ;
        RECT 1780.360 82.730 1781.880 82.870 ;
        RECT 1781.740 2.400 1781.880 82.730 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.830 386.480 739.150 386.540 ;
        RECT 742.050 386.480 742.370 386.540 ;
        RECT 738.830 386.340 742.370 386.480 ;
        RECT 738.830 386.280 739.150 386.340 ;
        RECT 742.050 386.280 742.370 386.340 ;
        RECT 738.830 115.840 739.150 115.900 ;
        RECT 1794.070 115.840 1794.390 115.900 ;
        RECT 738.830 115.700 1794.390 115.840 ;
        RECT 738.830 115.640 739.150 115.700 ;
        RECT 1794.070 115.640 1794.390 115.700 ;
      LAYER via ;
        RECT 738.860 386.280 739.120 386.540 ;
        RECT 742.080 386.280 742.340 386.540 ;
        RECT 738.860 115.640 739.120 115.900 ;
        RECT 1794.100 115.640 1794.360 115.900 ;
      LAYER met2 ;
        RECT 743.350 400.250 743.630 404.000 ;
        RECT 742.140 400.110 743.630 400.250 ;
        RECT 742.140 386.570 742.280 400.110 ;
        RECT 743.350 400.000 743.630 400.110 ;
        RECT 738.860 386.250 739.120 386.570 ;
        RECT 742.080 386.250 742.340 386.570 ;
        RECT 738.920 115.930 739.060 386.250 ;
        RECT 738.860 115.610 739.120 115.930 ;
        RECT 1794.100 115.610 1794.360 115.930 ;
        RECT 1794.160 82.870 1794.300 115.610 ;
        RECT 1794.160 82.730 1797.520 82.870 ;
        RECT 1797.380 1.770 1797.520 82.730 ;
        RECT 1799.470 1.770 1800.030 2.400 ;
        RECT 1797.380 1.630 1800.030 1.770 ;
        RECT 1799.470 -4.800 1800.030 1.630 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.270 386.140 745.590 386.200 ;
        RECT 747.570 386.140 747.890 386.200 ;
        RECT 745.270 386.000 747.890 386.140 ;
        RECT 745.270 385.940 745.590 386.000 ;
        RECT 747.570 385.940 747.890 386.000 ;
        RECT 745.270 43.080 745.590 43.140 ;
        RECT 1817.530 43.080 1817.850 43.140 ;
        RECT 745.270 42.940 1817.850 43.080 ;
        RECT 745.270 42.880 745.590 42.940 ;
        RECT 1817.530 42.880 1817.850 42.940 ;
      LAYER via ;
        RECT 745.300 385.940 745.560 386.200 ;
        RECT 747.600 385.940 747.860 386.200 ;
        RECT 745.300 42.880 745.560 43.140 ;
        RECT 1817.560 42.880 1817.820 43.140 ;
      LAYER met2 ;
        RECT 748.870 400.250 749.150 404.000 ;
        RECT 747.660 400.110 749.150 400.250 ;
        RECT 747.660 386.230 747.800 400.110 ;
        RECT 748.870 400.000 749.150 400.110 ;
        RECT 745.300 385.910 745.560 386.230 ;
        RECT 747.600 385.910 747.860 386.230 ;
        RECT 745.360 43.170 745.500 385.910 ;
        RECT 745.300 42.850 745.560 43.170 ;
        RECT 1817.560 42.850 1817.820 43.170 ;
        RECT 1817.620 2.400 1817.760 42.850 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.170 43.420 752.490 43.480 ;
        RECT 1835.010 43.420 1835.330 43.480 ;
        RECT 752.170 43.280 1835.330 43.420 ;
        RECT 752.170 43.220 752.490 43.280 ;
        RECT 1835.010 43.220 1835.330 43.280 ;
      LAYER via ;
        RECT 752.200 43.220 752.460 43.480 ;
        RECT 1835.040 43.220 1835.300 43.480 ;
      LAYER met2 ;
        RECT 753.930 400.250 754.210 404.000 ;
        RECT 752.720 400.110 754.210 400.250 ;
        RECT 752.720 386.480 752.860 400.110 ;
        RECT 753.930 400.000 754.210 400.110 ;
        RECT 752.260 386.340 752.860 386.480 ;
        RECT 752.260 43.510 752.400 386.340 ;
        RECT 752.200 43.190 752.460 43.510 ;
        RECT 1835.040 43.190 1835.300 43.510 ;
        RECT 1835.100 2.400 1835.240 43.190 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.070 48.180 759.390 48.240 ;
        RECT 765.050 48.180 765.370 48.240 ;
        RECT 759.070 48.040 765.370 48.180 ;
        RECT 759.070 47.980 759.390 48.040 ;
        RECT 765.050 47.980 765.370 48.040 ;
        RECT 765.050 43.760 765.370 43.820 ;
        RECT 1852.950 43.760 1853.270 43.820 ;
        RECT 765.050 43.620 1853.270 43.760 ;
        RECT 765.050 43.560 765.370 43.620 ;
        RECT 1852.950 43.560 1853.270 43.620 ;
      LAYER via ;
        RECT 759.100 47.980 759.360 48.240 ;
        RECT 765.080 47.980 765.340 48.240 ;
        RECT 765.080 43.560 765.340 43.820 ;
        RECT 1852.980 43.560 1853.240 43.820 ;
      LAYER met2 ;
        RECT 759.450 400.250 759.730 404.000 ;
        RECT 759.160 400.110 759.730 400.250 ;
        RECT 759.160 48.270 759.300 400.110 ;
        RECT 759.450 400.000 759.730 400.110 ;
        RECT 759.100 47.950 759.360 48.270 ;
        RECT 765.080 47.950 765.340 48.270 ;
        RECT 765.140 43.850 765.280 47.950 ;
        RECT 765.080 43.530 765.340 43.850 ;
        RECT 1852.980 43.530 1853.240 43.850 ;
        RECT 1853.040 2.400 1853.180 43.530 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.890 27.100 422.210 27.160 ;
        RECT 735.610 27.100 735.930 27.160 ;
        RECT 421.890 26.960 735.930 27.100 ;
        RECT 421.890 26.900 422.210 26.960 ;
        RECT 735.610 26.900 735.930 26.960 ;
      LAYER via ;
        RECT 421.920 26.900 422.180 27.160 ;
        RECT 735.640 26.900 735.900 27.160 ;
      LAYER met2 ;
        RECT 421.810 400.180 422.090 404.000 ;
        RECT 421.810 400.000 422.120 400.180 ;
        RECT 421.980 27.190 422.120 400.000 ;
        RECT 421.920 26.870 422.180 27.190 ;
        RECT 735.640 26.870 735.900 27.190 ;
        RECT 735.700 2.400 735.840 26.870 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.530 386.480 759.850 386.540 ;
        RECT 763.670 386.480 763.990 386.540 ;
        RECT 759.530 386.340 763.990 386.480 ;
        RECT 759.530 386.280 759.850 386.340 ;
        RECT 763.670 386.280 763.990 386.340 ;
        RECT 759.530 44.100 759.850 44.160 ;
        RECT 1870.430 44.100 1870.750 44.160 ;
        RECT 759.530 43.960 1870.750 44.100 ;
        RECT 759.530 43.900 759.850 43.960 ;
        RECT 1870.430 43.900 1870.750 43.960 ;
      LAYER via ;
        RECT 759.560 386.280 759.820 386.540 ;
        RECT 763.700 386.280 763.960 386.540 ;
        RECT 759.560 43.900 759.820 44.160 ;
        RECT 1870.460 43.900 1870.720 44.160 ;
      LAYER met2 ;
        RECT 764.970 400.250 765.250 404.000 ;
        RECT 763.760 400.110 765.250 400.250 ;
        RECT 763.760 386.570 763.900 400.110 ;
        RECT 764.970 400.000 765.250 400.110 ;
        RECT 759.560 386.250 759.820 386.570 ;
        RECT 763.700 386.250 763.960 386.570 ;
        RECT 759.620 44.190 759.760 386.250 ;
        RECT 759.560 43.870 759.820 44.190 ;
        RECT 1870.460 43.870 1870.720 44.190 ;
        RECT 1870.520 2.400 1870.660 43.870 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.970 386.480 766.290 386.540 ;
        RECT 768.730 386.480 769.050 386.540 ;
        RECT 765.970 386.340 769.050 386.480 ;
        RECT 765.970 386.280 766.290 386.340 ;
        RECT 768.730 386.280 769.050 386.340 ;
        RECT 765.970 44.440 766.290 44.500 ;
        RECT 1888.370 44.440 1888.690 44.500 ;
        RECT 765.970 44.300 1888.690 44.440 ;
        RECT 765.970 44.240 766.290 44.300 ;
        RECT 1888.370 44.240 1888.690 44.300 ;
      LAYER via ;
        RECT 766.000 386.280 766.260 386.540 ;
        RECT 768.760 386.280 769.020 386.540 ;
        RECT 766.000 44.240 766.260 44.500 ;
        RECT 1888.400 44.240 1888.660 44.500 ;
      LAYER met2 ;
        RECT 770.030 400.250 770.310 404.000 ;
        RECT 768.820 400.110 770.310 400.250 ;
        RECT 768.820 386.570 768.960 400.110 ;
        RECT 770.030 400.000 770.310 400.110 ;
        RECT 766.000 386.250 766.260 386.570 ;
        RECT 768.760 386.250 769.020 386.570 ;
        RECT 766.060 44.530 766.200 386.250 ;
        RECT 766.000 44.210 766.260 44.530 ;
        RECT 1888.400 44.210 1888.660 44.530 ;
        RECT 1888.460 2.400 1888.600 44.210 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 772.870 48.180 773.190 48.240 ;
        RECT 1905.850 48.180 1906.170 48.240 ;
        RECT 772.870 48.040 1906.170 48.180 ;
        RECT 772.870 47.980 773.190 48.040 ;
        RECT 1905.850 47.980 1906.170 48.040 ;
      LAYER via ;
        RECT 772.900 47.980 773.160 48.240 ;
        RECT 1905.880 47.980 1906.140 48.240 ;
      LAYER met2 ;
        RECT 775.550 400.250 775.830 404.000 ;
        RECT 774.340 400.110 775.830 400.250 ;
        RECT 774.340 386.470 774.480 400.110 ;
        RECT 775.550 400.000 775.830 400.110 ;
        RECT 772.960 386.330 774.480 386.470 ;
        RECT 772.960 48.270 773.100 386.330 ;
        RECT 772.900 47.950 773.160 48.270 ;
        RECT 1905.880 47.950 1906.140 48.270 ;
        RECT 1905.940 2.400 1906.080 47.950 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.230 47.840 780.550 47.900 ;
        RECT 1923.790 47.840 1924.110 47.900 ;
        RECT 780.230 47.700 1924.110 47.840 ;
        RECT 780.230 47.640 780.550 47.700 ;
        RECT 1923.790 47.640 1924.110 47.700 ;
      LAYER via ;
        RECT 780.260 47.640 780.520 47.900 ;
        RECT 1923.820 47.640 1924.080 47.900 ;
      LAYER met2 ;
        RECT 780.610 400.250 780.890 404.000 ;
        RECT 780.320 400.110 780.890 400.250 ;
        RECT 780.320 47.930 780.460 400.110 ;
        RECT 780.610 400.000 780.890 400.110 ;
        RECT 780.260 47.610 780.520 47.930 ;
        RECT 1923.820 47.610 1924.080 47.930 ;
        RECT 1923.880 2.400 1924.020 47.610 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 779.770 386.480 780.090 386.540 ;
        RECT 784.830 386.480 785.150 386.540 ;
        RECT 779.770 386.340 785.150 386.480 ;
        RECT 779.770 386.280 780.090 386.340 ;
        RECT 784.830 386.280 785.150 386.340 ;
        RECT 779.770 47.500 780.090 47.560 ;
        RECT 1941.270 47.500 1941.590 47.560 ;
        RECT 779.770 47.360 1941.590 47.500 ;
        RECT 779.770 47.300 780.090 47.360 ;
        RECT 1941.270 47.300 1941.590 47.360 ;
      LAYER via ;
        RECT 779.800 386.280 780.060 386.540 ;
        RECT 784.860 386.280 785.120 386.540 ;
        RECT 779.800 47.300 780.060 47.560 ;
        RECT 1941.300 47.300 1941.560 47.560 ;
      LAYER met2 ;
        RECT 786.130 400.250 786.410 404.000 ;
        RECT 784.920 400.110 786.410 400.250 ;
        RECT 784.920 386.570 785.060 400.110 ;
        RECT 786.130 400.000 786.410 400.110 ;
        RECT 779.800 386.250 780.060 386.570 ;
        RECT 784.860 386.250 785.120 386.570 ;
        RECT 779.860 47.590 780.000 386.250 ;
        RECT 779.800 47.270 780.060 47.590 ;
        RECT 1941.300 47.270 1941.560 47.590 ;
        RECT 1941.360 2.400 1941.500 47.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 786.670 386.480 786.990 386.540 ;
        RECT 790.350 386.480 790.670 386.540 ;
        RECT 786.670 386.340 790.670 386.480 ;
        RECT 786.670 386.280 786.990 386.340 ;
        RECT 790.350 386.280 790.670 386.340 ;
        RECT 786.670 47.160 786.990 47.220 ;
        RECT 1959.210 47.160 1959.530 47.220 ;
        RECT 786.670 47.020 1959.530 47.160 ;
        RECT 786.670 46.960 786.990 47.020 ;
        RECT 1959.210 46.960 1959.530 47.020 ;
      LAYER via ;
        RECT 786.700 386.280 786.960 386.540 ;
        RECT 790.380 386.280 790.640 386.540 ;
        RECT 786.700 46.960 786.960 47.220 ;
        RECT 1959.240 46.960 1959.500 47.220 ;
      LAYER met2 ;
        RECT 791.650 400.250 791.930 404.000 ;
        RECT 790.440 400.110 791.930 400.250 ;
        RECT 790.440 386.570 790.580 400.110 ;
        RECT 791.650 400.000 791.930 400.110 ;
        RECT 786.700 386.250 786.960 386.570 ;
        RECT 790.380 386.250 790.640 386.570 ;
        RECT 786.760 47.250 786.900 386.250 ;
        RECT 786.700 46.930 786.960 47.250 ;
        RECT 1959.240 46.930 1959.500 47.250 ;
        RECT 1959.300 2.400 1959.440 46.930 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 793.570 386.480 793.890 386.540 ;
        RECT 795.870 386.480 796.190 386.540 ;
        RECT 793.570 386.340 796.190 386.480 ;
        RECT 793.570 386.280 793.890 386.340 ;
        RECT 795.870 386.280 796.190 386.340 ;
        RECT 793.570 46.820 793.890 46.880 ;
        RECT 1976.690 46.820 1977.010 46.880 ;
        RECT 793.570 46.680 1977.010 46.820 ;
        RECT 793.570 46.620 793.890 46.680 ;
        RECT 1976.690 46.620 1977.010 46.680 ;
      LAYER via ;
        RECT 793.600 386.280 793.860 386.540 ;
        RECT 795.900 386.280 796.160 386.540 ;
        RECT 793.600 46.620 793.860 46.880 ;
        RECT 1976.720 46.620 1976.980 46.880 ;
      LAYER met2 ;
        RECT 796.710 400.250 796.990 404.000 ;
        RECT 795.960 400.110 796.990 400.250 ;
        RECT 795.960 386.570 796.100 400.110 ;
        RECT 796.710 400.000 796.990 400.110 ;
        RECT 793.600 386.250 793.860 386.570 ;
        RECT 795.900 386.250 796.160 386.570 ;
        RECT 793.660 46.910 793.800 386.250 ;
        RECT 793.600 46.590 793.860 46.910 ;
        RECT 1976.720 46.590 1976.980 46.910 ;
        RECT 1976.780 2.400 1976.920 46.590 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.470 46.480 800.790 46.540 ;
        RECT 1994.630 46.480 1994.950 46.540 ;
        RECT 800.470 46.340 1994.950 46.480 ;
        RECT 800.470 46.280 800.790 46.340 ;
        RECT 1994.630 46.280 1994.950 46.340 ;
      LAYER via ;
        RECT 800.500 46.280 800.760 46.540 ;
        RECT 1994.660 46.280 1994.920 46.540 ;
      LAYER met2 ;
        RECT 802.230 400.250 802.510 404.000 ;
        RECT 801.020 400.110 802.510 400.250 ;
        RECT 801.020 385.970 801.160 400.110 ;
        RECT 802.230 400.000 802.510 400.110 ;
        RECT 800.560 385.830 801.160 385.970 ;
        RECT 800.560 46.570 800.700 385.830 ;
        RECT 800.500 46.250 800.760 46.570 ;
        RECT 1994.660 46.250 1994.920 46.570 ;
        RECT 1994.720 2.400 1994.860 46.250 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.830 46.140 808.150 46.200 ;
        RECT 2012.570 46.140 2012.890 46.200 ;
        RECT 807.830 46.000 2012.890 46.140 ;
        RECT 807.830 45.940 808.150 46.000 ;
        RECT 2012.570 45.940 2012.890 46.000 ;
      LAYER via ;
        RECT 807.860 45.940 808.120 46.200 ;
        RECT 2012.600 45.940 2012.860 46.200 ;
      LAYER met2 ;
        RECT 807.750 400.180 808.030 404.000 ;
        RECT 807.750 400.000 808.060 400.180 ;
        RECT 807.920 46.230 808.060 400.000 ;
        RECT 807.860 45.910 808.120 46.230 ;
        RECT 2012.600 45.910 2012.860 46.230 ;
        RECT 2012.660 2.400 2012.800 45.910 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.370 386.480 807.690 386.540 ;
        RECT 811.510 386.480 811.830 386.540 ;
        RECT 807.370 386.340 811.830 386.480 ;
        RECT 807.370 386.280 807.690 386.340 ;
        RECT 811.510 386.280 811.830 386.340 ;
        RECT 807.370 45.800 807.690 45.860 ;
        RECT 2030.050 45.800 2030.370 45.860 ;
        RECT 807.370 45.660 2030.370 45.800 ;
        RECT 807.370 45.600 807.690 45.660 ;
        RECT 2030.050 45.600 2030.370 45.660 ;
      LAYER via ;
        RECT 807.400 386.280 807.660 386.540 ;
        RECT 811.540 386.280 811.800 386.540 ;
        RECT 807.400 45.600 807.660 45.860 ;
        RECT 2030.080 45.600 2030.340 45.860 ;
      LAYER met2 ;
        RECT 812.810 400.250 813.090 404.000 ;
        RECT 811.600 400.110 813.090 400.250 ;
        RECT 811.600 386.570 811.740 400.110 ;
        RECT 812.810 400.000 813.090 400.110 ;
        RECT 807.400 386.250 807.660 386.570 ;
        RECT 811.540 386.250 811.800 386.570 ;
        RECT 807.460 45.890 807.600 386.250 ;
        RECT 807.400 45.570 807.660 45.890 ;
        RECT 2030.080 45.570 2030.340 45.890 ;
        RECT 2030.140 2.400 2030.280 45.570 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.430 386.140 421.750 386.200 ;
        RECT 426.030 386.140 426.350 386.200 ;
        RECT 421.430 386.000 426.350 386.140 ;
        RECT 421.430 385.940 421.750 386.000 ;
        RECT 426.030 385.940 426.350 386.000 ;
        RECT 421.430 26.760 421.750 26.820 ;
        RECT 753.090 26.760 753.410 26.820 ;
        RECT 421.430 26.620 753.410 26.760 ;
        RECT 421.430 26.560 421.750 26.620 ;
        RECT 753.090 26.560 753.410 26.620 ;
      LAYER via ;
        RECT 421.460 385.940 421.720 386.200 ;
        RECT 426.060 385.940 426.320 386.200 ;
        RECT 421.460 26.560 421.720 26.820 ;
        RECT 753.120 26.560 753.380 26.820 ;
      LAYER met2 ;
        RECT 427.330 400.250 427.610 404.000 ;
        RECT 426.120 400.110 427.610 400.250 ;
        RECT 426.120 386.230 426.260 400.110 ;
        RECT 427.330 400.000 427.610 400.110 ;
        RECT 421.460 385.910 421.720 386.230 ;
        RECT 426.060 385.910 426.320 386.230 ;
        RECT 421.520 26.850 421.660 385.910 ;
        RECT 421.460 26.530 421.720 26.850 ;
        RECT 753.120 26.530 753.380 26.850 ;
        RECT 753.180 2.400 753.320 26.530 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.270 386.480 814.590 386.540 ;
        RECT 817.030 386.480 817.350 386.540 ;
        RECT 814.270 386.340 817.350 386.480 ;
        RECT 814.270 386.280 814.590 386.340 ;
        RECT 817.030 386.280 817.350 386.340 ;
        RECT 814.270 45.460 814.590 45.520 ;
        RECT 2047.990 45.460 2048.310 45.520 ;
        RECT 814.270 45.320 2048.310 45.460 ;
        RECT 814.270 45.260 814.590 45.320 ;
        RECT 2047.990 45.260 2048.310 45.320 ;
      LAYER via ;
        RECT 814.300 386.280 814.560 386.540 ;
        RECT 817.060 386.280 817.320 386.540 ;
        RECT 814.300 45.260 814.560 45.520 ;
        RECT 2048.020 45.260 2048.280 45.520 ;
      LAYER met2 ;
        RECT 818.330 400.250 818.610 404.000 ;
        RECT 817.120 400.110 818.610 400.250 ;
        RECT 817.120 386.570 817.260 400.110 ;
        RECT 818.330 400.000 818.610 400.110 ;
        RECT 814.300 386.250 814.560 386.570 ;
        RECT 817.060 386.250 817.320 386.570 ;
        RECT 814.360 45.550 814.500 386.250 ;
        RECT 814.300 45.230 814.560 45.550 ;
        RECT 2048.020 45.230 2048.280 45.550 ;
        RECT 2048.080 2.400 2048.220 45.230 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.170 386.480 821.490 386.540 ;
        RECT 822.550 386.480 822.870 386.540 ;
        RECT 821.170 386.340 822.870 386.480 ;
        RECT 821.170 386.280 821.490 386.340 ;
        RECT 822.550 386.280 822.870 386.340 ;
        RECT 821.170 45.120 821.490 45.180 ;
        RECT 2065.470 45.120 2065.790 45.180 ;
        RECT 821.170 44.980 2065.790 45.120 ;
        RECT 821.170 44.920 821.490 44.980 ;
        RECT 2065.470 44.920 2065.790 44.980 ;
      LAYER via ;
        RECT 821.200 386.280 821.460 386.540 ;
        RECT 822.580 386.280 822.840 386.540 ;
        RECT 821.200 44.920 821.460 45.180 ;
        RECT 2065.500 44.920 2065.760 45.180 ;
      LAYER met2 ;
        RECT 823.850 400.250 824.130 404.000 ;
        RECT 822.640 400.110 824.130 400.250 ;
        RECT 822.640 386.570 822.780 400.110 ;
        RECT 823.850 400.000 824.130 400.110 ;
        RECT 821.200 386.250 821.460 386.570 ;
        RECT 822.580 386.250 822.840 386.570 ;
        RECT 821.260 45.210 821.400 386.250 ;
        RECT 821.200 44.890 821.460 45.210 ;
        RECT 2065.500 44.890 2065.760 45.210 ;
        RECT 2065.560 2.400 2065.700 44.890 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.530 44.780 828.850 44.840 ;
        RECT 2083.410 44.780 2083.730 44.840 ;
        RECT 828.530 44.640 2083.730 44.780 ;
        RECT 828.530 44.580 828.850 44.640 ;
        RECT 2083.410 44.580 2083.730 44.640 ;
      LAYER via ;
        RECT 828.560 44.580 828.820 44.840 ;
        RECT 2083.440 44.580 2083.700 44.840 ;
      LAYER met2 ;
        RECT 828.910 400.250 829.190 404.000 ;
        RECT 828.620 400.110 829.190 400.250 ;
        RECT 828.620 44.870 828.760 400.110 ;
        RECT 828.910 400.000 829.190 400.110 ;
        RECT 828.560 44.550 828.820 44.870 ;
        RECT 2083.440 44.550 2083.700 44.870 ;
        RECT 2083.500 2.400 2083.640 44.550 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.070 386.480 828.390 386.540 ;
        RECT 833.130 386.480 833.450 386.540 ;
        RECT 828.070 386.340 833.450 386.480 ;
        RECT 828.070 386.280 828.390 386.340 ;
        RECT 833.130 386.280 833.450 386.340 ;
      LAYER via ;
        RECT 828.100 386.280 828.360 386.540 ;
        RECT 833.160 386.280 833.420 386.540 ;
      LAYER met2 ;
        RECT 834.430 400.250 834.710 404.000 ;
        RECT 833.220 400.110 834.710 400.250 ;
        RECT 833.220 386.570 833.360 400.110 ;
        RECT 834.430 400.000 834.710 400.110 ;
        RECT 828.100 386.250 828.360 386.570 ;
        RECT 833.160 386.250 833.420 386.570 ;
        RECT 828.160 44.725 828.300 386.250 ;
        RECT 828.090 44.355 828.370 44.725 ;
        RECT 2100.910 44.355 2101.190 44.725 ;
        RECT 2100.980 2.400 2101.120 44.355 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
      LAYER via2 ;
        RECT 828.090 44.400 828.370 44.680 ;
        RECT 2100.910 44.400 2101.190 44.680 ;
      LAYER met3 ;
        RECT 828.065 44.690 828.395 44.705 ;
        RECT 2100.885 44.690 2101.215 44.705 ;
        RECT 828.065 44.390 2101.215 44.690 ;
        RECT 828.065 44.375 828.395 44.390 ;
        RECT 2100.885 44.375 2101.215 44.390 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.890 109.380 836.210 109.440 ;
        RECT 2118.370 109.380 2118.690 109.440 ;
        RECT 835.890 109.240 2118.690 109.380 ;
        RECT 835.890 109.180 836.210 109.240 ;
        RECT 2118.370 109.180 2118.690 109.240 ;
      LAYER via ;
        RECT 835.920 109.180 836.180 109.440 ;
        RECT 2118.400 109.180 2118.660 109.440 ;
      LAYER met2 ;
        RECT 839.950 400.250 840.230 404.000 ;
        RECT 838.740 400.110 840.230 400.250 ;
        RECT 838.740 324.370 838.880 400.110 ;
        RECT 839.950 400.000 840.230 400.110 ;
        RECT 835.980 324.230 838.880 324.370 ;
        RECT 835.980 109.470 836.120 324.230 ;
        RECT 835.920 109.150 836.180 109.470 ;
        RECT 2118.400 109.150 2118.660 109.470 ;
        RECT 2118.460 15.370 2118.600 109.150 ;
        RECT 2118.460 15.230 2119.060 15.370 ;
        RECT 2118.920 2.400 2119.060 15.230 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.790 115.500 843.110 115.560 ;
        RECT 2132.170 115.500 2132.490 115.560 ;
        RECT 842.790 115.360 2132.490 115.500 ;
        RECT 842.790 115.300 843.110 115.360 ;
        RECT 2132.170 115.300 2132.490 115.360 ;
      LAYER via ;
        RECT 842.820 115.300 843.080 115.560 ;
        RECT 2132.200 115.300 2132.460 115.560 ;
      LAYER met2 ;
        RECT 845.010 400.250 845.290 404.000 ;
        RECT 843.800 400.110 845.290 400.250 ;
        RECT 843.800 324.370 843.940 400.110 ;
        RECT 845.010 400.000 845.290 400.110 ;
        RECT 842.880 324.230 843.940 324.370 ;
        RECT 842.880 115.590 843.020 324.230 ;
        RECT 842.820 115.270 843.080 115.590 ;
        RECT 2132.200 115.270 2132.460 115.590 ;
        RECT 2132.260 82.870 2132.400 115.270 ;
        RECT 2132.260 82.730 2134.240 82.870 ;
        RECT 2134.100 1.770 2134.240 82.730 ;
        RECT 2136.190 1.770 2136.750 2.400 ;
        RECT 2134.100 1.630 2136.750 1.770 ;
        RECT 2136.190 -4.800 2136.750 1.630 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 850.150 115.160 850.470 115.220 ;
        RECT 2152.870 115.160 2153.190 115.220 ;
        RECT 850.150 115.020 2153.190 115.160 ;
        RECT 850.150 114.960 850.470 115.020 ;
        RECT 2152.870 114.960 2153.190 115.020 ;
      LAYER via ;
        RECT 850.180 114.960 850.440 115.220 ;
        RECT 2152.900 114.960 2153.160 115.220 ;
      LAYER met2 ;
        RECT 850.530 400.250 850.810 404.000 ;
        RECT 850.240 400.110 850.810 400.250 ;
        RECT 850.240 115.250 850.380 400.110 ;
        RECT 850.530 400.000 850.810 400.110 ;
        RECT 850.180 114.930 850.440 115.250 ;
        RECT 2152.900 114.930 2153.160 115.250 ;
        RECT 2152.960 82.870 2153.100 114.930 ;
        RECT 2152.960 82.730 2154.480 82.870 ;
        RECT 2154.340 2.400 2154.480 82.730 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.590 114.820 856.910 114.880 ;
        RECT 2166.670 114.820 2166.990 114.880 ;
        RECT 856.590 114.680 2166.990 114.820 ;
        RECT 856.590 114.620 856.910 114.680 ;
        RECT 2166.670 114.620 2166.990 114.680 ;
      LAYER via ;
        RECT 856.620 114.620 856.880 114.880 ;
        RECT 2166.700 114.620 2166.960 114.880 ;
      LAYER met2 ;
        RECT 856.050 400.250 856.330 404.000 ;
        RECT 856.050 400.110 856.820 400.250 ;
        RECT 856.050 400.000 856.330 400.110 ;
        RECT 856.680 114.910 856.820 400.110 ;
        RECT 856.620 114.590 856.880 114.910 ;
        RECT 2166.700 114.590 2166.960 114.910 ;
        RECT 2166.760 82.870 2166.900 114.590 ;
        RECT 2166.760 82.730 2170.120 82.870 ;
        RECT 2169.980 1.770 2170.120 82.730 ;
        RECT 2172.070 1.770 2172.630 2.400 ;
        RECT 2169.980 1.630 2172.630 1.770 ;
        RECT 2172.070 -4.800 2172.630 1.630 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 857.050 114.480 857.370 114.540 ;
        RECT 2187.370 114.480 2187.690 114.540 ;
        RECT 857.050 114.340 2187.690 114.480 ;
        RECT 857.050 114.280 857.370 114.340 ;
        RECT 2187.370 114.280 2187.690 114.340 ;
      LAYER via ;
        RECT 857.080 114.280 857.340 114.540 ;
        RECT 2187.400 114.280 2187.660 114.540 ;
      LAYER met2 ;
        RECT 861.110 400.250 861.390 404.000 ;
        RECT 859.900 400.110 861.390 400.250 ;
        RECT 859.900 324.370 860.040 400.110 ;
        RECT 861.110 400.000 861.390 400.110 ;
        RECT 857.140 324.230 860.040 324.370 ;
        RECT 857.140 114.570 857.280 324.230 ;
        RECT 857.080 114.250 857.340 114.570 ;
        RECT 2187.400 114.250 2187.660 114.570 ;
        RECT 2187.460 1.770 2187.600 114.250 ;
        RECT 2189.550 1.770 2190.110 2.400 ;
        RECT 2187.460 1.630 2190.110 1.770 ;
        RECT 2189.550 -4.800 2190.110 1.630 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.030 376.620 863.350 376.680 ;
        RECT 865.330 376.620 865.650 376.680 ;
        RECT 863.030 376.480 865.650 376.620 ;
        RECT 863.030 376.420 863.350 376.480 ;
        RECT 865.330 376.420 865.650 376.480 ;
        RECT 863.030 50.220 863.350 50.280 ;
        RECT 2201.630 50.220 2201.950 50.280 ;
        RECT 863.030 50.080 2201.950 50.220 ;
        RECT 863.030 50.020 863.350 50.080 ;
        RECT 2201.630 50.020 2201.950 50.080 ;
        RECT 2201.630 16.900 2201.950 16.960 ;
        RECT 2207.610 16.900 2207.930 16.960 ;
        RECT 2201.630 16.760 2207.930 16.900 ;
        RECT 2201.630 16.700 2201.950 16.760 ;
        RECT 2207.610 16.700 2207.930 16.760 ;
      LAYER via ;
        RECT 863.060 376.420 863.320 376.680 ;
        RECT 865.360 376.420 865.620 376.680 ;
        RECT 863.060 50.020 863.320 50.280 ;
        RECT 2201.660 50.020 2201.920 50.280 ;
        RECT 2201.660 16.700 2201.920 16.960 ;
        RECT 2207.640 16.700 2207.900 16.960 ;
      LAYER met2 ;
        RECT 866.630 400.250 866.910 404.000 ;
        RECT 865.420 400.110 866.910 400.250 ;
        RECT 865.420 376.710 865.560 400.110 ;
        RECT 866.630 400.000 866.910 400.110 ;
        RECT 863.060 376.390 863.320 376.710 ;
        RECT 865.360 376.390 865.620 376.710 ;
        RECT 863.120 50.310 863.260 376.390 ;
        RECT 863.060 49.990 863.320 50.310 ;
        RECT 2201.660 49.990 2201.920 50.310 ;
        RECT 2201.720 16.990 2201.860 49.990 ;
        RECT 2201.660 16.670 2201.920 16.990 ;
        RECT 2207.640 16.670 2207.900 16.990 ;
        RECT 2207.700 2.400 2207.840 16.670 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.330 385.800 428.650 385.860 ;
        RECT 431.090 385.800 431.410 385.860 ;
        RECT 428.330 385.660 431.410 385.800 ;
        RECT 428.330 385.600 428.650 385.660 ;
        RECT 431.090 385.600 431.410 385.660 ;
        RECT 428.330 29.140 428.650 29.200 ;
        RECT 611.870 29.140 612.190 29.200 ;
        RECT 428.330 29.000 612.190 29.140 ;
        RECT 428.330 28.940 428.650 29.000 ;
        RECT 611.870 28.940 612.190 29.000 ;
        RECT 611.870 16.900 612.190 16.960 ;
        RECT 771.030 16.900 771.350 16.960 ;
        RECT 611.870 16.760 771.350 16.900 ;
        RECT 611.870 16.700 612.190 16.760 ;
        RECT 771.030 16.700 771.350 16.760 ;
      LAYER via ;
        RECT 428.360 385.600 428.620 385.860 ;
        RECT 431.120 385.600 431.380 385.860 ;
        RECT 428.360 28.940 428.620 29.200 ;
        RECT 611.900 28.940 612.160 29.200 ;
        RECT 611.900 16.700 612.160 16.960 ;
        RECT 771.060 16.700 771.320 16.960 ;
      LAYER met2 ;
        RECT 432.390 400.250 432.670 404.000 ;
        RECT 431.180 400.110 432.670 400.250 ;
        RECT 431.180 385.890 431.320 400.110 ;
        RECT 432.390 400.000 432.670 400.110 ;
        RECT 428.360 385.570 428.620 385.890 ;
        RECT 431.120 385.570 431.380 385.890 ;
        RECT 428.420 29.230 428.560 385.570 ;
        RECT 428.360 28.910 428.620 29.230 ;
        RECT 611.900 28.910 612.160 29.230 ;
        RECT 611.960 16.990 612.100 28.910 ;
        RECT 611.900 16.670 612.160 16.990 ;
        RECT 771.060 16.670 771.320 16.990 ;
        RECT 771.120 2.400 771.260 16.670 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 870.390 50.560 870.710 50.620 ;
        RECT 2225.090 50.560 2225.410 50.620 ;
        RECT 870.390 50.420 2225.410 50.560 ;
        RECT 870.390 50.360 870.710 50.420 ;
        RECT 2225.090 50.360 2225.410 50.420 ;
      LAYER via ;
        RECT 870.420 50.360 870.680 50.620 ;
        RECT 2225.120 50.360 2225.380 50.620 ;
      LAYER met2 ;
        RECT 871.690 400.250 871.970 404.000 ;
        RECT 870.940 400.110 871.970 400.250 ;
        RECT 870.940 351.970 871.080 400.110 ;
        RECT 871.690 400.000 871.970 400.110 ;
        RECT 870.480 351.830 871.080 351.970 ;
        RECT 870.480 50.650 870.620 351.830 ;
        RECT 870.420 50.330 870.680 50.650 ;
        RECT 2225.120 50.330 2225.380 50.650 ;
        RECT 2225.180 2.400 2225.320 50.330 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.830 50.900 877.150 50.960 ;
        RECT 2243.030 50.900 2243.350 50.960 ;
        RECT 876.830 50.760 2243.350 50.900 ;
        RECT 876.830 50.700 877.150 50.760 ;
        RECT 2243.030 50.700 2243.350 50.760 ;
      LAYER via ;
        RECT 876.860 50.700 877.120 50.960 ;
        RECT 2243.060 50.700 2243.320 50.960 ;
      LAYER met2 ;
        RECT 877.210 400.250 877.490 404.000 ;
        RECT 876.920 400.110 877.490 400.250 ;
        RECT 876.920 50.990 877.060 400.110 ;
        RECT 877.210 400.000 877.490 400.110 ;
        RECT 876.860 50.670 877.120 50.990 ;
        RECT 2243.060 50.670 2243.320 50.990 ;
        RECT 2243.120 2.400 2243.260 50.670 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 877.290 376.280 877.610 376.340 ;
        RECT 881.430 376.280 881.750 376.340 ;
        RECT 877.290 376.140 881.750 376.280 ;
        RECT 877.290 376.080 877.610 376.140 ;
        RECT 881.430 376.080 881.750 376.140 ;
        RECT 877.290 51.240 877.610 51.300 ;
        RECT 2258.210 51.240 2258.530 51.300 ;
        RECT 877.290 51.100 2258.530 51.240 ;
        RECT 877.290 51.040 877.610 51.100 ;
        RECT 2258.210 51.040 2258.530 51.100 ;
      LAYER via ;
        RECT 877.320 376.080 877.580 376.340 ;
        RECT 881.460 376.080 881.720 376.340 ;
        RECT 877.320 51.040 877.580 51.300 ;
        RECT 2258.240 51.040 2258.500 51.300 ;
      LAYER met2 ;
        RECT 882.730 400.250 883.010 404.000 ;
        RECT 881.520 400.110 883.010 400.250 ;
        RECT 881.520 376.370 881.660 400.110 ;
        RECT 882.730 400.000 883.010 400.110 ;
        RECT 877.320 376.050 877.580 376.370 ;
        RECT 881.460 376.050 881.720 376.370 ;
        RECT 877.380 51.330 877.520 376.050 ;
        RECT 877.320 51.010 877.580 51.330 ;
        RECT 2258.240 51.010 2258.500 51.330 ;
        RECT 2258.300 1.770 2258.440 51.010 ;
        RECT 2260.390 1.770 2260.950 2.400 ;
        RECT 2258.300 1.630 2260.950 1.770 ;
        RECT 2260.390 -4.800 2260.950 1.630 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.730 376.280 884.050 376.340 ;
        RECT 886.950 376.280 887.270 376.340 ;
        RECT 883.730 376.140 887.270 376.280 ;
        RECT 883.730 376.080 884.050 376.140 ;
        RECT 886.950 376.080 887.270 376.140 ;
        RECT 883.730 54.980 884.050 55.040 ;
        RECT 2278.450 54.980 2278.770 55.040 ;
        RECT 883.730 54.840 2278.770 54.980 ;
        RECT 883.730 54.780 884.050 54.840 ;
        RECT 2278.450 54.780 2278.770 54.840 ;
      LAYER via ;
        RECT 883.760 376.080 884.020 376.340 ;
        RECT 886.980 376.080 887.240 376.340 ;
        RECT 883.760 54.780 884.020 55.040 ;
        RECT 2278.480 54.780 2278.740 55.040 ;
      LAYER met2 ;
        RECT 887.790 400.250 888.070 404.000 ;
        RECT 887.040 400.110 888.070 400.250 ;
        RECT 887.040 376.370 887.180 400.110 ;
        RECT 887.790 400.000 888.070 400.110 ;
        RECT 883.760 376.050 884.020 376.370 ;
        RECT 886.980 376.050 887.240 376.370 ;
        RECT 883.820 55.070 883.960 376.050 ;
        RECT 883.760 54.750 884.020 55.070 ;
        RECT 2278.480 54.750 2278.740 55.070 ;
        RECT 2278.540 2.400 2278.680 54.750 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.630 54.640 890.950 54.700 ;
        RECT 2295.930 54.640 2296.250 54.700 ;
        RECT 890.630 54.500 2296.250 54.640 ;
        RECT 890.630 54.440 890.950 54.500 ;
        RECT 2295.930 54.440 2296.250 54.500 ;
      LAYER via ;
        RECT 890.660 54.440 890.920 54.700 ;
        RECT 2295.960 54.440 2296.220 54.700 ;
      LAYER met2 ;
        RECT 893.310 400.250 893.590 404.000 ;
        RECT 892.100 400.110 893.590 400.250 ;
        RECT 892.100 351.970 892.240 400.110 ;
        RECT 893.310 400.000 893.590 400.110 ;
        RECT 890.720 351.830 892.240 351.970 ;
        RECT 890.720 54.730 890.860 351.830 ;
        RECT 890.660 54.410 890.920 54.730 ;
        RECT 2295.960 54.410 2296.220 54.730 ;
        RECT 2296.020 2.400 2296.160 54.410 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.990 54.300 898.310 54.360 ;
        RECT 2311.570 54.300 2311.890 54.360 ;
        RECT 897.990 54.160 2311.890 54.300 ;
        RECT 897.990 54.100 898.310 54.160 ;
        RECT 2311.570 54.100 2311.890 54.160 ;
      LAYER via ;
        RECT 898.020 54.100 898.280 54.360 ;
        RECT 2311.600 54.100 2311.860 54.360 ;
      LAYER met2 ;
        RECT 898.830 400.250 899.110 404.000 ;
        RECT 898.080 400.110 899.110 400.250 ;
        RECT 898.080 54.390 898.220 400.110 ;
        RECT 898.830 400.000 899.110 400.110 ;
        RECT 898.020 54.070 898.280 54.390 ;
        RECT 2311.600 54.070 2311.860 54.390 ;
        RECT 2311.660 1.770 2311.800 54.070 ;
        RECT 2313.750 1.770 2314.310 2.400 ;
        RECT 2311.660 1.630 2314.310 1.770 ;
        RECT 2313.750 -4.800 2314.310 1.630 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.890 53.960 905.210 54.020 ;
        RECT 2329.050 53.960 2329.370 54.020 ;
        RECT 904.890 53.820 2329.370 53.960 ;
        RECT 904.890 53.760 905.210 53.820 ;
        RECT 2329.050 53.760 2329.370 53.820 ;
      LAYER via ;
        RECT 904.920 53.760 905.180 54.020 ;
        RECT 2329.080 53.760 2329.340 54.020 ;
      LAYER met2 ;
        RECT 903.890 400.250 904.170 404.000 ;
        RECT 903.890 400.110 905.120 400.250 ;
        RECT 903.890 400.000 904.170 400.110 ;
        RECT 904.980 54.050 905.120 400.110 ;
        RECT 904.920 53.730 905.180 54.050 ;
        RECT 2329.080 53.730 2329.340 54.050 ;
        RECT 2329.140 1.770 2329.280 53.730 ;
        RECT 2331.230 1.770 2331.790 2.400 ;
        RECT 2329.140 1.630 2331.790 1.770 ;
        RECT 2331.230 -4.800 2331.790 1.630 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.430 376.280 904.750 376.340 ;
        RECT 908.110 376.280 908.430 376.340 ;
        RECT 904.430 376.140 908.430 376.280 ;
        RECT 904.430 376.080 904.750 376.140 ;
        RECT 908.110 376.080 908.430 376.140 ;
        RECT 904.430 53.620 904.750 53.680 ;
        RECT 2349.290 53.620 2349.610 53.680 ;
        RECT 904.430 53.480 2349.610 53.620 ;
        RECT 904.430 53.420 904.750 53.480 ;
        RECT 2349.290 53.420 2349.610 53.480 ;
      LAYER via ;
        RECT 904.460 376.080 904.720 376.340 ;
        RECT 908.140 376.080 908.400 376.340 ;
        RECT 904.460 53.420 904.720 53.680 ;
        RECT 2349.320 53.420 2349.580 53.680 ;
      LAYER met2 ;
        RECT 909.410 400.250 909.690 404.000 ;
        RECT 908.200 400.110 909.690 400.250 ;
        RECT 908.200 376.370 908.340 400.110 ;
        RECT 909.410 400.000 909.690 400.110 ;
        RECT 904.460 376.050 904.720 376.370 ;
        RECT 908.140 376.050 908.400 376.370 ;
        RECT 904.520 53.710 904.660 376.050 ;
        RECT 904.460 53.390 904.720 53.710 ;
        RECT 2349.320 53.390 2349.580 53.710 ;
        RECT 2349.380 2.400 2349.520 53.390 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.330 375.940 911.650 376.000 ;
        RECT 913.630 375.940 913.950 376.000 ;
        RECT 911.330 375.800 913.950 375.940 ;
        RECT 911.330 375.740 911.650 375.800 ;
        RECT 913.630 375.740 913.950 375.800 ;
        RECT 911.330 53.280 911.650 53.340 ;
        RECT 2367.230 53.280 2367.550 53.340 ;
        RECT 911.330 53.140 2367.550 53.280 ;
        RECT 911.330 53.080 911.650 53.140 ;
        RECT 2367.230 53.080 2367.550 53.140 ;
      LAYER via ;
        RECT 911.360 375.740 911.620 376.000 ;
        RECT 913.660 375.740 913.920 376.000 ;
        RECT 911.360 53.080 911.620 53.340 ;
        RECT 2367.260 53.080 2367.520 53.340 ;
      LAYER met2 ;
        RECT 914.930 400.250 915.210 404.000 ;
        RECT 913.720 400.110 915.210 400.250 ;
        RECT 913.720 376.030 913.860 400.110 ;
        RECT 914.930 400.000 915.210 400.110 ;
        RECT 911.360 375.710 911.620 376.030 ;
        RECT 913.660 375.710 913.920 376.030 ;
        RECT 911.420 53.370 911.560 375.710 ;
        RECT 911.360 53.050 911.620 53.370 ;
        RECT 2367.260 53.050 2367.520 53.370 ;
        RECT 2367.320 2.400 2367.460 53.050 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.690 52.940 919.010 53.000 ;
        RECT 2382.410 52.940 2382.730 53.000 ;
        RECT 918.690 52.800 2382.730 52.940 ;
        RECT 918.690 52.740 919.010 52.800 ;
        RECT 2382.410 52.740 2382.730 52.800 ;
      LAYER via ;
        RECT 918.720 52.740 918.980 53.000 ;
        RECT 2382.440 52.740 2382.700 53.000 ;
      LAYER met2 ;
        RECT 919.990 400.250 920.270 404.000 ;
        RECT 918.780 400.110 920.270 400.250 ;
        RECT 918.780 53.030 918.920 400.110 ;
        RECT 919.990 400.000 920.270 400.110 ;
        RECT 918.720 52.710 918.980 53.030 ;
        RECT 2382.440 52.710 2382.700 53.030 ;
        RECT 2382.500 1.770 2382.640 52.710 ;
        RECT 2384.590 1.770 2385.150 2.400 ;
        RECT 2382.500 1.630 2385.150 1.770 ;
        RECT 2384.590 -4.800 2385.150 1.630 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.230 31.520 435.550 31.580 ;
        RECT 788.970 31.520 789.290 31.580 ;
        RECT 435.230 31.380 789.290 31.520 ;
        RECT 435.230 31.320 435.550 31.380 ;
        RECT 788.970 31.320 789.290 31.380 ;
      LAYER via ;
        RECT 435.260 31.320 435.520 31.580 ;
        RECT 789.000 31.320 789.260 31.580 ;
      LAYER met2 ;
        RECT 437.910 400.250 438.190 404.000 ;
        RECT 436.700 400.110 438.190 400.250 ;
        RECT 436.700 386.480 436.840 400.110 ;
        RECT 437.910 400.000 438.190 400.110 ;
        RECT 435.320 386.340 436.840 386.480 ;
        RECT 435.320 31.610 435.460 386.340 ;
        RECT 435.260 31.290 435.520 31.610 ;
        RECT 789.000 31.290 789.260 31.610 ;
        RECT 789.060 2.400 789.200 31.290 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.930 29.480 387.250 29.540 ;
        RECT 634.870 29.480 635.190 29.540 ;
        RECT 386.930 29.340 635.190 29.480 ;
        RECT 386.930 29.280 387.250 29.340 ;
        RECT 634.870 29.280 635.190 29.340 ;
      LAYER via ;
        RECT 386.960 29.280 387.220 29.540 ;
        RECT 634.900 29.280 635.160 29.540 ;
      LAYER met2 ;
        RECT 391.450 400.250 391.730 404.000 ;
        RECT 390.240 400.110 391.730 400.250 ;
        RECT 390.240 399.570 390.380 400.110 ;
        RECT 391.450 400.000 391.730 400.110 ;
        RECT 389.320 399.430 390.380 399.570 ;
        RECT 389.320 351.970 389.460 399.430 ;
        RECT 387.020 351.830 389.460 351.970 ;
        RECT 387.020 29.570 387.160 351.830 ;
        RECT 386.960 29.250 387.220 29.570 ;
        RECT 634.900 29.250 635.160 29.570 ;
        RECT 634.960 2.400 635.100 29.250 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 924.670 399.740 924.990 399.800 ;
        RECT 926.050 399.740 926.370 399.800 ;
        RECT 924.670 399.600 926.370 399.740 ;
        RECT 924.670 399.540 924.990 399.600 ;
        RECT 926.050 399.540 926.370 399.600 ;
        RECT 924.670 52.600 924.990 52.660 ;
        RECT 2408.630 52.600 2408.950 52.660 ;
        RECT 924.670 52.460 2408.950 52.600 ;
        RECT 924.670 52.400 924.990 52.460 ;
        RECT 2408.630 52.400 2408.950 52.460 ;
      LAYER via ;
        RECT 924.700 399.540 924.960 399.800 ;
        RECT 926.080 399.540 926.340 399.800 ;
        RECT 924.700 52.400 924.960 52.660 ;
        RECT 2408.660 52.400 2408.920 52.660 ;
      LAYER met2 ;
        RECT 927.350 400.250 927.630 404.000 ;
        RECT 926.140 400.110 927.630 400.250 ;
        RECT 926.140 399.830 926.280 400.110 ;
        RECT 927.350 400.000 927.630 400.110 ;
        RECT 924.700 399.510 924.960 399.830 ;
        RECT 926.080 399.510 926.340 399.830 ;
        RECT 924.760 52.690 924.900 399.510 ;
        RECT 924.700 52.370 924.960 52.690 ;
        RECT 2408.660 52.370 2408.920 52.690 ;
        RECT 2408.720 2.400 2408.860 52.370 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 52.260 931.890 52.320 ;
        RECT 2423.810 52.260 2424.130 52.320 ;
        RECT 931.570 52.120 2424.130 52.260 ;
        RECT 931.570 52.060 931.890 52.120 ;
        RECT 2423.810 52.060 2424.130 52.120 ;
      LAYER via ;
        RECT 931.600 52.060 931.860 52.320 ;
        RECT 2423.840 52.060 2424.100 52.320 ;
      LAYER met2 ;
        RECT 932.870 400.250 933.150 404.000 ;
        RECT 931.660 400.110 933.150 400.250 ;
        RECT 931.660 52.350 931.800 400.110 ;
        RECT 932.870 400.000 933.150 400.110 ;
        RECT 931.600 52.030 931.860 52.350 ;
        RECT 2423.840 52.030 2424.100 52.350 ;
        RECT 2423.900 1.770 2424.040 52.030 ;
        RECT 2425.990 1.770 2426.550 2.400 ;
        RECT 2423.900 1.630 2426.550 1.770 ;
        RECT 2425.990 -4.800 2426.550 1.630 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.030 376.280 932.350 376.340 ;
        RECT 936.630 376.280 936.950 376.340 ;
        RECT 932.030 376.140 936.950 376.280 ;
        RECT 932.030 376.080 932.350 376.140 ;
        RECT 936.630 376.080 936.950 376.140 ;
        RECT 932.030 51.920 932.350 51.980 ;
        RECT 2444.050 51.920 2444.370 51.980 ;
        RECT 932.030 51.780 2444.370 51.920 ;
        RECT 932.030 51.720 932.350 51.780 ;
        RECT 2444.050 51.720 2444.370 51.780 ;
      LAYER via ;
        RECT 932.060 376.080 932.320 376.340 ;
        RECT 936.660 376.080 936.920 376.340 ;
        RECT 932.060 51.720 932.320 51.980 ;
        RECT 2444.080 51.720 2444.340 51.980 ;
      LAYER met2 ;
        RECT 937.930 400.250 938.210 404.000 ;
        RECT 936.720 400.110 938.210 400.250 ;
        RECT 936.720 376.370 936.860 400.110 ;
        RECT 937.930 400.000 938.210 400.110 ;
        RECT 932.060 376.050 932.320 376.370 ;
        RECT 936.660 376.050 936.920 376.370 ;
        RECT 932.120 52.010 932.260 376.050 ;
        RECT 932.060 51.690 932.320 52.010 ;
        RECT 2444.080 51.690 2444.340 52.010 ;
        RECT 2444.140 2.400 2444.280 51.690 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.470 376.280 938.790 376.340 ;
        RECT 942.150 376.280 942.470 376.340 ;
        RECT 938.470 376.140 942.470 376.280 ;
        RECT 938.470 376.080 938.790 376.140 ;
        RECT 942.150 376.080 942.470 376.140 ;
        RECT 938.470 51.580 938.790 51.640 ;
        RECT 2461.530 51.580 2461.850 51.640 ;
        RECT 938.470 51.440 2461.850 51.580 ;
        RECT 938.470 51.380 938.790 51.440 ;
        RECT 2461.530 51.380 2461.850 51.440 ;
      LAYER via ;
        RECT 938.500 376.080 938.760 376.340 ;
        RECT 942.180 376.080 942.440 376.340 ;
        RECT 938.500 51.380 938.760 51.640 ;
        RECT 2461.560 51.380 2461.820 51.640 ;
      LAYER met2 ;
        RECT 943.450 400.250 943.730 404.000 ;
        RECT 942.240 400.110 943.730 400.250 ;
        RECT 942.240 376.370 942.380 400.110 ;
        RECT 943.450 400.000 943.730 400.110 ;
        RECT 938.500 376.050 938.760 376.370 ;
        RECT 942.180 376.050 942.440 376.370 ;
        RECT 938.560 51.670 938.700 376.050 ;
        RECT 938.500 51.350 938.760 51.670 ;
        RECT 2461.560 51.350 2461.820 51.670 ;
        RECT 2461.620 2.400 2461.760 51.350 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.370 375.940 945.690 376.000 ;
        RECT 947.670 375.940 947.990 376.000 ;
        RECT 945.370 375.800 947.990 375.940 ;
        RECT 945.370 375.740 945.690 375.800 ;
        RECT 947.670 375.740 947.990 375.800 ;
      LAYER via ;
        RECT 945.400 375.740 945.660 376.000 ;
        RECT 947.700 375.740 947.960 376.000 ;
      LAYER met2 ;
        RECT 948.510 400.250 948.790 404.000 ;
        RECT 947.760 400.110 948.790 400.250 ;
        RECT 947.760 376.030 947.900 400.110 ;
        RECT 948.510 400.000 948.790 400.110 ;
        RECT 945.400 375.710 945.660 376.030 ;
        RECT 947.700 375.710 947.960 376.030 ;
        RECT 945.460 52.205 945.600 375.710 ;
        RECT 945.390 51.835 945.670 52.205 ;
        RECT 2477.190 51.835 2477.470 52.205 ;
        RECT 2477.260 1.770 2477.400 51.835 ;
        RECT 2479.350 1.770 2479.910 2.400 ;
        RECT 2477.260 1.630 2479.910 1.770 ;
        RECT 2479.350 -4.800 2479.910 1.630 ;
      LAYER via2 ;
        RECT 945.390 51.880 945.670 52.160 ;
        RECT 2477.190 51.880 2477.470 52.160 ;
      LAYER met3 ;
        RECT 945.365 52.170 945.695 52.185 ;
        RECT 2477.165 52.170 2477.495 52.185 ;
        RECT 945.365 51.870 2477.495 52.170 ;
        RECT 945.365 51.855 945.695 51.870 ;
        RECT 2477.165 51.855 2477.495 51.870 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.030 400.250 954.310 404.000 ;
        RECT 953.280 400.110 954.310 400.250 ;
        RECT 953.280 51.525 953.420 400.110 ;
        RECT 954.030 400.000 954.310 400.110 ;
        RECT 953.210 51.155 953.490 51.525 ;
        RECT 2494.670 51.155 2494.950 51.525 ;
        RECT 2494.740 1.770 2494.880 51.155 ;
        RECT 2496.830 1.770 2497.390 2.400 ;
        RECT 2494.740 1.630 2497.390 1.770 ;
        RECT 2496.830 -4.800 2497.390 1.630 ;
      LAYER via2 ;
        RECT 953.210 51.200 953.490 51.480 ;
        RECT 2494.670 51.200 2494.950 51.480 ;
      LAYER met3 ;
        RECT 953.185 51.490 953.515 51.505 ;
        RECT 2494.645 51.490 2494.975 51.505 ;
        RECT 953.185 51.190 2494.975 51.490 ;
        RECT 953.185 51.175 953.515 51.190 ;
        RECT 2494.645 51.175 2494.975 51.190 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.630 392.940 959.950 393.000 ;
        RECT 961.010 392.940 961.330 393.000 ;
        RECT 959.630 392.800 961.330 392.940 ;
        RECT 959.630 392.740 959.950 392.800 ;
        RECT 961.010 392.740 961.330 392.800 ;
        RECT 960.090 114.140 960.410 114.200 ;
        RECT 2511.670 114.140 2511.990 114.200 ;
        RECT 960.090 114.000 2511.990 114.140 ;
        RECT 960.090 113.940 960.410 114.000 ;
        RECT 2511.670 113.940 2511.990 114.000 ;
      LAYER via ;
        RECT 959.660 392.740 959.920 393.000 ;
        RECT 961.040 392.740 961.300 393.000 ;
        RECT 960.120 113.940 960.380 114.200 ;
        RECT 2511.700 113.940 2511.960 114.200 ;
      LAYER met2 ;
        RECT 959.550 400.180 959.830 404.000 ;
        RECT 959.550 400.000 959.860 400.180 ;
        RECT 959.720 393.030 959.860 400.000 ;
        RECT 959.660 392.710 959.920 393.030 ;
        RECT 961.040 392.710 961.300 393.030 ;
        RECT 961.100 386.470 961.240 392.710 ;
        RECT 960.180 386.330 961.240 386.470 ;
        RECT 960.180 114.230 960.320 386.330 ;
        RECT 960.120 113.910 960.380 114.230 ;
        RECT 2511.700 113.910 2511.960 114.230 ;
        RECT 2511.760 82.870 2511.900 113.910 ;
        RECT 2511.760 82.730 2515.120 82.870 ;
        RECT 2514.980 2.400 2515.120 82.730 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.550 113.800 960.870 113.860 ;
        RECT 2532.370 113.800 2532.690 113.860 ;
        RECT 960.550 113.660 2532.690 113.800 ;
        RECT 960.550 113.600 960.870 113.660 ;
        RECT 2532.370 113.600 2532.690 113.660 ;
      LAYER via ;
        RECT 960.580 113.600 960.840 113.860 ;
        RECT 2532.400 113.600 2532.660 113.860 ;
      LAYER met2 ;
        RECT 964.610 400.250 964.890 404.000 ;
        RECT 963.860 400.110 964.890 400.250 ;
        RECT 963.860 324.370 964.000 400.110 ;
        RECT 964.610 400.000 964.890 400.110 ;
        RECT 960.640 324.230 964.000 324.370 ;
        RECT 960.640 113.890 960.780 324.230 ;
        RECT 960.580 113.570 960.840 113.890 ;
        RECT 2532.400 113.570 2532.660 113.890 ;
        RECT 2532.460 2.400 2532.600 113.570 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.130 400.250 970.410 404.000 ;
        RECT 968.920 400.110 970.410 400.250 ;
        RECT 968.920 324.370 969.060 400.110 ;
        RECT 970.130 400.000 970.410 400.110 ;
        RECT 967.540 324.230 969.060 324.370 ;
        RECT 967.540 114.085 967.680 324.230 ;
        RECT 967.470 113.715 967.750 114.085 ;
        RECT 2546.190 113.715 2546.470 114.085 ;
        RECT 2546.260 82.870 2546.400 113.715 ;
        RECT 2546.260 82.730 2548.240 82.870 ;
        RECT 2548.100 1.770 2548.240 82.730 ;
        RECT 2550.190 1.770 2550.750 2.400 ;
        RECT 2548.100 1.630 2550.750 1.770 ;
        RECT 2550.190 -4.800 2550.750 1.630 ;
      LAYER via2 ;
        RECT 967.470 113.760 967.750 114.040 ;
        RECT 2546.190 113.760 2546.470 114.040 ;
      LAYER met3 ;
        RECT 967.445 114.050 967.775 114.065 ;
        RECT 2546.165 114.050 2546.495 114.065 ;
        RECT 967.445 113.750 2546.495 114.050 ;
        RECT 967.445 113.735 967.775 113.750 ;
        RECT 2546.165 113.735 2546.495 113.750 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.650 400.250 975.930 404.000 ;
        RECT 974.440 400.110 975.930 400.250 ;
        RECT 974.440 113.405 974.580 400.110 ;
        RECT 975.650 400.000 975.930 400.110 ;
        RECT 974.370 113.035 974.650 113.405 ;
        RECT 2566.890 113.035 2567.170 113.405 ;
        RECT 2566.960 1.770 2567.100 113.035 ;
        RECT 2567.670 1.770 2568.230 2.400 ;
        RECT 2566.960 1.630 2568.230 1.770 ;
        RECT 2567.670 -4.800 2568.230 1.630 ;
      LAYER via2 ;
        RECT 974.370 113.080 974.650 113.360 ;
        RECT 2566.890 113.080 2567.170 113.360 ;
      LAYER met3 ;
        RECT 974.345 113.370 974.675 113.385 ;
        RECT 2566.865 113.370 2567.195 113.385 ;
        RECT 974.345 113.070 2567.195 113.370 ;
        RECT 974.345 113.055 974.675 113.070 ;
        RECT 2566.865 113.055 2567.195 113.070 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 387.840 441.990 387.900 ;
        RECT 443.970 387.840 444.290 387.900 ;
        RECT 441.670 387.700 444.290 387.840 ;
        RECT 441.670 387.640 441.990 387.700 ;
        RECT 443.970 387.640 444.290 387.700 ;
        RECT 442.130 31.180 442.450 31.240 ;
        RECT 812.430 31.180 812.750 31.240 ;
        RECT 442.130 31.040 812.750 31.180 ;
        RECT 442.130 30.980 442.450 31.040 ;
        RECT 812.430 30.980 812.750 31.040 ;
      LAYER via ;
        RECT 441.700 387.640 441.960 387.900 ;
        RECT 444.000 387.640 444.260 387.900 ;
        RECT 442.160 30.980 442.420 31.240 ;
        RECT 812.460 30.980 812.720 31.240 ;
      LAYER met2 ;
        RECT 444.810 400.250 445.090 404.000 ;
        RECT 444.060 400.110 445.090 400.250 ;
        RECT 444.060 387.930 444.200 400.110 ;
        RECT 444.810 400.000 445.090 400.110 ;
        RECT 441.700 387.610 441.960 387.930 ;
        RECT 444.000 387.610 444.260 387.930 ;
        RECT 441.760 372.670 441.900 387.610 ;
        RECT 441.760 372.530 442.360 372.670 ;
        RECT 442.220 31.270 442.360 372.530 ;
        RECT 442.160 30.950 442.420 31.270 ;
        RECT 812.460 30.950 812.720 31.270 ;
        RECT 812.520 2.400 812.660 30.950 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.330 57.360 980.650 57.420 ;
        RECT 2585.730 57.360 2586.050 57.420 ;
        RECT 980.330 57.220 2586.050 57.360 ;
        RECT 980.330 57.160 980.650 57.220 ;
        RECT 2585.730 57.160 2586.050 57.220 ;
      LAYER via ;
        RECT 980.360 57.160 980.620 57.420 ;
        RECT 2585.760 57.160 2586.020 57.420 ;
      LAYER met2 ;
        RECT 980.710 400.250 980.990 404.000 ;
        RECT 980.420 400.110 980.990 400.250 ;
        RECT 980.420 57.450 980.560 400.110 ;
        RECT 980.710 400.000 980.990 400.110 ;
        RECT 980.360 57.130 980.620 57.450 ;
        RECT 2585.760 57.130 2586.020 57.450 ;
        RECT 2585.820 2.400 2585.960 57.130 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.790 386.480 981.110 386.540 ;
        RECT 984.930 386.480 985.250 386.540 ;
        RECT 980.790 386.340 985.250 386.480 ;
        RECT 980.790 386.280 981.110 386.340 ;
        RECT 984.930 386.280 985.250 386.340 ;
        RECT 980.790 57.700 981.110 57.760 ;
        RECT 2601.370 57.700 2601.690 57.760 ;
        RECT 980.790 57.560 2601.690 57.700 ;
        RECT 980.790 57.500 981.110 57.560 ;
        RECT 2601.370 57.500 2601.690 57.560 ;
      LAYER via ;
        RECT 980.820 386.280 981.080 386.540 ;
        RECT 984.960 386.280 985.220 386.540 ;
        RECT 980.820 57.500 981.080 57.760 ;
        RECT 2601.400 57.500 2601.660 57.760 ;
      LAYER met2 ;
        RECT 986.230 400.250 986.510 404.000 ;
        RECT 985.020 400.110 986.510 400.250 ;
        RECT 985.020 386.570 985.160 400.110 ;
        RECT 986.230 400.000 986.510 400.110 ;
        RECT 980.820 386.250 981.080 386.570 ;
        RECT 984.960 386.250 985.220 386.570 ;
        RECT 980.880 57.790 981.020 386.250 ;
        RECT 980.820 57.470 981.080 57.790 ;
        RECT 2601.400 57.470 2601.660 57.790 ;
        RECT 2601.460 1.770 2601.600 57.470 ;
        RECT 2603.550 1.770 2604.110 2.400 ;
        RECT 2601.460 1.630 2604.110 1.770 ;
        RECT 2603.550 -4.800 2604.110 1.630 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.230 386.140 987.550 386.200 ;
        RECT 990.450 386.140 990.770 386.200 ;
        RECT 987.230 386.000 990.770 386.140 ;
        RECT 987.230 385.940 987.550 386.000 ;
        RECT 990.450 385.940 990.770 386.000 ;
        RECT 987.230 58.040 987.550 58.100 ;
        RECT 2618.850 58.040 2619.170 58.100 ;
        RECT 987.230 57.900 2619.170 58.040 ;
        RECT 987.230 57.840 987.550 57.900 ;
        RECT 2618.850 57.840 2619.170 57.900 ;
      LAYER via ;
        RECT 987.260 385.940 987.520 386.200 ;
        RECT 990.480 385.940 990.740 386.200 ;
        RECT 987.260 57.840 987.520 58.100 ;
        RECT 2618.880 57.840 2619.140 58.100 ;
      LAYER met2 ;
        RECT 991.750 400.250 992.030 404.000 ;
        RECT 990.540 400.110 992.030 400.250 ;
        RECT 990.540 386.230 990.680 400.110 ;
        RECT 991.750 400.000 992.030 400.110 ;
        RECT 987.260 385.910 987.520 386.230 ;
        RECT 990.480 385.910 990.740 386.230 ;
        RECT 987.320 58.130 987.460 385.910 ;
        RECT 987.260 57.810 987.520 58.130 ;
        RECT 2618.880 57.810 2619.140 58.130 ;
        RECT 2618.940 1.770 2619.080 57.810 ;
        RECT 2621.030 1.770 2621.590 2.400 ;
        RECT 2618.940 1.630 2621.590 1.770 ;
        RECT 2621.030 -4.800 2621.590 1.630 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.130 58.380 994.450 58.440 ;
        RECT 2639.090 58.380 2639.410 58.440 ;
        RECT 994.130 58.240 2639.410 58.380 ;
        RECT 994.130 58.180 994.450 58.240 ;
        RECT 2639.090 58.180 2639.410 58.240 ;
      LAYER via ;
        RECT 994.160 58.180 994.420 58.440 ;
        RECT 2639.120 58.180 2639.380 58.440 ;
      LAYER met2 ;
        RECT 996.810 400.250 997.090 404.000 ;
        RECT 995.600 400.110 997.090 400.250 ;
        RECT 995.600 385.970 995.740 400.110 ;
        RECT 996.810 400.000 997.090 400.110 ;
        RECT 994.220 385.830 995.740 385.970 ;
        RECT 994.220 58.470 994.360 385.830 ;
        RECT 994.160 58.150 994.420 58.470 ;
        RECT 2639.120 58.150 2639.380 58.470 ;
        RECT 2639.180 2.400 2639.320 58.150 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.490 62.120 1001.810 62.180 ;
        RECT 2657.030 62.120 2657.350 62.180 ;
        RECT 1001.490 61.980 2657.350 62.120 ;
        RECT 1001.490 61.920 1001.810 61.980 ;
        RECT 2657.030 61.920 2657.350 61.980 ;
      LAYER via ;
        RECT 1001.520 61.920 1001.780 62.180 ;
        RECT 2657.060 61.920 2657.320 62.180 ;
      LAYER met2 ;
        RECT 1002.330 400.250 1002.610 404.000 ;
        RECT 1001.580 400.110 1002.610 400.250 ;
        RECT 1001.580 62.210 1001.720 400.110 ;
        RECT 1002.330 400.000 1002.610 400.110 ;
        RECT 1001.520 61.890 1001.780 62.210 ;
        RECT 2657.060 61.890 2657.320 62.210 ;
        RECT 2657.120 16.730 2657.260 61.890 ;
        RECT 2656.660 16.590 2657.260 16.730 ;
        RECT 2656.660 2.400 2656.800 16.590 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1008.390 61.780 1008.710 61.840 ;
        RECT 2672.210 61.780 2672.530 61.840 ;
        RECT 1008.390 61.640 2672.530 61.780 ;
        RECT 1008.390 61.580 1008.710 61.640 ;
        RECT 2672.210 61.580 2672.530 61.640 ;
      LAYER via ;
        RECT 1008.420 61.580 1008.680 61.840 ;
        RECT 2672.240 61.580 2672.500 61.840 ;
      LAYER met2 ;
        RECT 1007.850 400.250 1008.130 404.000 ;
        RECT 1007.850 400.110 1008.620 400.250 ;
        RECT 1007.850 400.000 1008.130 400.110 ;
        RECT 1008.480 61.870 1008.620 400.110 ;
        RECT 1008.420 61.550 1008.680 61.870 ;
        RECT 2672.240 61.550 2672.500 61.870 ;
        RECT 2672.300 1.770 2672.440 61.550 ;
        RECT 2674.390 1.770 2674.950 2.400 ;
        RECT 2672.300 1.630 2674.950 1.770 ;
        RECT 2674.390 -4.800 2674.950 1.630 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.930 386.140 1008.250 386.200 ;
        RECT 1011.610 386.140 1011.930 386.200 ;
        RECT 1007.930 386.000 1011.930 386.140 ;
        RECT 1007.930 385.940 1008.250 386.000 ;
        RECT 1011.610 385.940 1011.930 386.000 ;
        RECT 1007.930 61.440 1008.250 61.500 ;
        RECT 2691.070 61.440 2691.390 61.500 ;
        RECT 1007.930 61.300 2691.390 61.440 ;
        RECT 1007.930 61.240 1008.250 61.300 ;
        RECT 2691.070 61.240 2691.390 61.300 ;
      LAYER via ;
        RECT 1007.960 385.940 1008.220 386.200 ;
        RECT 1011.640 385.940 1011.900 386.200 ;
        RECT 1007.960 61.240 1008.220 61.500 ;
        RECT 2691.100 61.240 2691.360 61.500 ;
      LAYER met2 ;
        RECT 1012.910 400.250 1013.190 404.000 ;
        RECT 1011.700 400.110 1013.190 400.250 ;
        RECT 1011.700 386.230 1011.840 400.110 ;
        RECT 1012.910 400.000 1013.190 400.110 ;
        RECT 1007.960 385.910 1008.220 386.230 ;
        RECT 1011.640 385.910 1011.900 386.230 ;
        RECT 1008.020 61.530 1008.160 385.910 ;
        RECT 1007.960 61.210 1008.220 61.530 ;
        RECT 2691.100 61.210 2691.360 61.530 ;
        RECT 2691.160 1.770 2691.300 61.210 ;
        RECT 2691.870 1.770 2692.430 2.400 ;
        RECT 2691.160 1.630 2692.430 1.770 ;
        RECT 2691.870 -4.800 2692.430 1.630 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.830 386.140 1015.150 386.200 ;
        RECT 1017.130 386.140 1017.450 386.200 ;
        RECT 1014.830 386.000 1017.450 386.140 ;
        RECT 1014.830 385.940 1015.150 386.000 ;
        RECT 1017.130 385.940 1017.450 386.000 ;
        RECT 1014.830 61.100 1015.150 61.160 ;
        RECT 2709.930 61.100 2710.250 61.160 ;
        RECT 1014.830 60.960 2710.250 61.100 ;
        RECT 1014.830 60.900 1015.150 60.960 ;
        RECT 2709.930 60.900 2710.250 60.960 ;
      LAYER via ;
        RECT 1014.860 385.940 1015.120 386.200 ;
        RECT 1017.160 385.940 1017.420 386.200 ;
        RECT 1014.860 60.900 1015.120 61.160 ;
        RECT 2709.960 60.900 2710.220 61.160 ;
      LAYER met2 ;
        RECT 1018.430 400.250 1018.710 404.000 ;
        RECT 1017.220 400.110 1018.710 400.250 ;
        RECT 1017.220 386.230 1017.360 400.110 ;
        RECT 1018.430 400.000 1018.710 400.110 ;
        RECT 1014.860 385.910 1015.120 386.230 ;
        RECT 1017.160 385.910 1017.420 386.230 ;
        RECT 1014.920 61.190 1015.060 385.910 ;
        RECT 1014.860 60.870 1015.120 61.190 ;
        RECT 2709.960 60.870 2710.220 61.190 ;
        RECT 2710.020 2.400 2710.160 60.870 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.190 60.760 1022.510 60.820 ;
        RECT 2727.410 60.760 2727.730 60.820 ;
        RECT 1022.190 60.620 2727.730 60.760 ;
        RECT 1022.190 60.560 1022.510 60.620 ;
        RECT 2727.410 60.560 2727.730 60.620 ;
      LAYER via ;
        RECT 1022.220 60.560 1022.480 60.820 ;
        RECT 2727.440 60.560 2727.700 60.820 ;
      LAYER met2 ;
        RECT 1023.950 400.250 1024.230 404.000 ;
        RECT 1022.740 400.110 1024.230 400.250 ;
        RECT 1022.740 386.650 1022.880 400.110 ;
        RECT 1023.950 400.000 1024.230 400.110 ;
        RECT 1022.280 386.510 1022.880 386.650 ;
        RECT 1022.280 60.850 1022.420 386.510 ;
        RECT 1022.220 60.530 1022.480 60.850 ;
        RECT 2727.440 60.530 2727.700 60.850 ;
        RECT 2727.500 2.400 2727.640 60.530 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1029.090 60.420 1029.410 60.480 ;
        RECT 2743.050 60.420 2743.370 60.480 ;
        RECT 1029.090 60.280 2743.370 60.420 ;
        RECT 1029.090 60.220 1029.410 60.280 ;
        RECT 2743.050 60.220 2743.370 60.280 ;
      LAYER via ;
        RECT 1029.120 60.220 1029.380 60.480 ;
        RECT 2743.080 60.220 2743.340 60.480 ;
      LAYER met2 ;
        RECT 1029.010 400.180 1029.290 404.000 ;
        RECT 1029.010 400.000 1029.320 400.180 ;
        RECT 1029.180 60.510 1029.320 400.000 ;
        RECT 1029.120 60.190 1029.380 60.510 ;
        RECT 2743.080 60.190 2743.340 60.510 ;
        RECT 2743.140 1.770 2743.280 60.190 ;
        RECT 2745.230 1.770 2745.790 2.400 ;
        RECT 2743.140 1.630 2745.790 1.770 ;
        RECT 2745.230 -4.800 2745.790 1.630 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 30.840 448.890 30.900 ;
        RECT 830.370 30.840 830.690 30.900 ;
        RECT 448.570 30.700 830.690 30.840 ;
        RECT 448.570 30.640 448.890 30.700 ;
        RECT 830.370 30.640 830.690 30.700 ;
      LAYER via ;
        RECT 448.600 30.640 448.860 30.900 ;
        RECT 830.400 30.640 830.660 30.900 ;
      LAYER met2 ;
        RECT 450.330 400.250 450.610 404.000 ;
        RECT 449.120 400.110 450.610 400.250 ;
        RECT 449.120 386.480 449.260 400.110 ;
        RECT 450.330 400.000 450.610 400.110 ;
        RECT 448.660 386.340 449.260 386.480 ;
        RECT 448.660 30.930 448.800 386.340 ;
        RECT 448.600 30.610 448.860 30.930 ;
        RECT 830.400 30.610 830.660 30.930 ;
        RECT 830.460 2.400 830.600 30.610 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.630 375.940 1028.950 376.000 ;
        RECT 1033.230 375.940 1033.550 376.000 ;
        RECT 1028.630 375.800 1033.550 375.940 ;
        RECT 1028.630 375.740 1028.950 375.800 ;
        RECT 1033.230 375.740 1033.550 375.800 ;
        RECT 1028.630 60.080 1028.950 60.140 ;
        RECT 2763.290 60.080 2763.610 60.140 ;
        RECT 1028.630 59.940 2763.610 60.080 ;
        RECT 1028.630 59.880 1028.950 59.940 ;
        RECT 2763.290 59.880 2763.610 59.940 ;
      LAYER via ;
        RECT 1028.660 375.740 1028.920 376.000 ;
        RECT 1033.260 375.740 1033.520 376.000 ;
        RECT 1028.660 59.880 1028.920 60.140 ;
        RECT 2763.320 59.880 2763.580 60.140 ;
      LAYER met2 ;
        RECT 1034.530 400.250 1034.810 404.000 ;
        RECT 1033.320 400.110 1034.810 400.250 ;
        RECT 1033.320 376.030 1033.460 400.110 ;
        RECT 1034.530 400.000 1034.810 400.110 ;
        RECT 1028.660 375.710 1028.920 376.030 ;
        RECT 1033.260 375.710 1033.520 376.030 ;
        RECT 1028.720 60.170 1028.860 375.710 ;
        RECT 1028.660 59.850 1028.920 60.170 ;
        RECT 2763.320 59.850 2763.580 60.170 ;
        RECT 2763.380 2.400 2763.520 59.850 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.530 376.280 1035.850 376.340 ;
        RECT 1038.750 376.280 1039.070 376.340 ;
        RECT 1035.530 376.140 1039.070 376.280 ;
        RECT 1035.530 376.080 1035.850 376.140 ;
        RECT 1038.750 376.080 1039.070 376.140 ;
        RECT 1035.530 59.740 1035.850 59.800 ;
        RECT 2781.230 59.740 2781.550 59.800 ;
        RECT 1035.530 59.600 2781.550 59.740 ;
        RECT 1035.530 59.540 1035.850 59.600 ;
        RECT 2781.230 59.540 2781.550 59.600 ;
      LAYER via ;
        RECT 1035.560 376.080 1035.820 376.340 ;
        RECT 1038.780 376.080 1039.040 376.340 ;
        RECT 1035.560 59.540 1035.820 59.800 ;
        RECT 2781.260 59.540 2781.520 59.800 ;
      LAYER met2 ;
        RECT 1039.590 400.250 1039.870 404.000 ;
        RECT 1038.840 400.110 1039.870 400.250 ;
        RECT 1038.840 376.370 1038.980 400.110 ;
        RECT 1039.590 400.000 1039.870 400.110 ;
        RECT 1035.560 376.050 1035.820 376.370 ;
        RECT 1038.780 376.050 1039.040 376.370 ;
        RECT 1035.620 59.830 1035.760 376.050 ;
        RECT 1035.560 59.510 1035.820 59.830 ;
        RECT 2781.260 59.510 2781.520 59.830 ;
        RECT 2781.320 16.730 2781.460 59.510 ;
        RECT 2780.860 16.590 2781.460 16.730 ;
        RECT 2780.860 2.400 2781.000 16.590 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.970 375.940 1042.290 376.000 ;
        RECT 1043.810 375.940 1044.130 376.000 ;
        RECT 1041.970 375.800 1044.130 375.940 ;
        RECT 1041.970 375.740 1042.290 375.800 ;
        RECT 1043.810 375.740 1044.130 375.800 ;
        RECT 1041.970 59.400 1042.290 59.460 ;
        RECT 2796.410 59.400 2796.730 59.460 ;
        RECT 1041.970 59.260 2796.730 59.400 ;
        RECT 1041.970 59.200 1042.290 59.260 ;
        RECT 2796.410 59.200 2796.730 59.260 ;
      LAYER via ;
        RECT 1042.000 375.740 1042.260 376.000 ;
        RECT 1043.840 375.740 1044.100 376.000 ;
        RECT 1042.000 59.200 1042.260 59.460 ;
        RECT 2796.440 59.200 2796.700 59.460 ;
      LAYER met2 ;
        RECT 1045.110 400.250 1045.390 404.000 ;
        RECT 1043.900 400.110 1045.390 400.250 ;
        RECT 1043.900 376.030 1044.040 400.110 ;
        RECT 1045.110 400.000 1045.390 400.110 ;
        RECT 1042.000 375.710 1042.260 376.030 ;
        RECT 1043.840 375.710 1044.100 376.030 ;
        RECT 1042.060 59.490 1042.200 375.710 ;
        RECT 1042.000 59.170 1042.260 59.490 ;
        RECT 2796.440 59.170 2796.700 59.490 ;
        RECT 2796.500 1.770 2796.640 59.170 ;
        RECT 2798.590 1.770 2799.150 2.400 ;
        RECT 2796.500 1.630 2799.150 1.770 ;
        RECT 2798.590 -4.800 2799.150 1.630 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1048.870 375.940 1049.190 376.000 ;
        RECT 1050.250 375.940 1050.570 376.000 ;
        RECT 1048.870 375.800 1050.570 375.940 ;
        RECT 1048.870 375.740 1049.190 375.800 ;
        RECT 1050.250 375.740 1050.570 375.800 ;
        RECT 1048.870 59.060 1049.190 59.120 ;
        RECT 2815.270 59.060 2815.590 59.120 ;
        RECT 1048.870 58.920 2815.590 59.060 ;
        RECT 1048.870 58.860 1049.190 58.920 ;
        RECT 2815.270 58.860 2815.590 58.920 ;
      LAYER via ;
        RECT 1048.900 375.740 1049.160 376.000 ;
        RECT 1050.280 375.740 1050.540 376.000 ;
        RECT 1048.900 58.860 1049.160 59.120 ;
        RECT 2815.300 58.860 2815.560 59.120 ;
      LAYER met2 ;
        RECT 1050.630 400.250 1050.910 404.000 ;
        RECT 1050.340 400.110 1050.910 400.250 ;
        RECT 1050.340 376.030 1050.480 400.110 ;
        RECT 1050.630 400.000 1050.910 400.110 ;
        RECT 1048.900 375.710 1049.160 376.030 ;
        RECT 1050.280 375.710 1050.540 376.030 ;
        RECT 1048.960 59.150 1049.100 375.710 ;
        RECT 1048.900 58.830 1049.160 59.150 ;
        RECT 2815.300 58.830 2815.560 59.150 ;
        RECT 2815.360 1.770 2815.500 58.830 ;
        RECT 2816.070 1.770 2816.630 2.400 ;
        RECT 2815.360 1.630 2816.630 1.770 ;
        RECT 2816.070 -4.800 2816.630 1.630 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.690 400.250 1055.970 404.000 ;
        RECT 1055.690 400.110 1056.460 400.250 ;
        RECT 1055.690 400.000 1055.970 400.110 ;
        RECT 1056.320 59.005 1056.460 400.110 ;
        RECT 1056.250 58.635 1056.530 59.005 ;
        RECT 2834.150 58.635 2834.430 59.005 ;
        RECT 2834.220 2.400 2834.360 58.635 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
      LAYER via2 ;
        RECT 1056.250 58.680 1056.530 58.960 ;
        RECT 2834.150 58.680 2834.430 58.960 ;
      LAYER met3 ;
        RECT 1056.225 58.970 1056.555 58.985 ;
        RECT 2834.125 58.970 2834.455 58.985 ;
        RECT 1056.225 58.670 2834.455 58.970 ;
        RECT 1056.225 58.655 1056.555 58.670 ;
        RECT 2834.125 58.655 2834.455 58.670 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.210 400.250 1061.490 404.000 ;
        RECT 1060.000 400.110 1061.490 400.250 ;
        RECT 1060.000 324.370 1060.140 400.110 ;
        RECT 1061.210 400.000 1061.490 400.110 ;
        RECT 1057.240 324.230 1060.140 324.370 ;
        RECT 1057.240 58.325 1057.380 324.230 ;
        RECT 1057.170 57.955 1057.450 58.325 ;
        RECT 2851.630 57.955 2851.910 58.325 ;
        RECT 2851.700 2.400 2851.840 57.955 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
      LAYER via2 ;
        RECT 1057.170 58.000 1057.450 58.280 ;
        RECT 2851.630 58.000 2851.910 58.280 ;
      LAYER met3 ;
        RECT 1057.145 58.290 1057.475 58.305 ;
        RECT 2851.605 58.290 2851.935 58.305 ;
        RECT 1057.145 57.990 2851.935 58.290 ;
        RECT 1057.145 57.975 1057.475 57.990 ;
        RECT 2851.605 57.975 2851.935 57.990 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.130 375.940 1063.450 376.000 ;
        RECT 1065.430 375.940 1065.750 376.000 ;
        RECT 1063.130 375.800 1065.750 375.940 ;
        RECT 1063.130 375.740 1063.450 375.800 ;
        RECT 1065.430 375.740 1065.750 375.800 ;
        RECT 1063.130 58.720 1063.450 58.780 ;
        RECT 2867.250 58.720 2867.570 58.780 ;
        RECT 1063.130 58.580 2867.570 58.720 ;
        RECT 1063.130 58.520 1063.450 58.580 ;
        RECT 2867.250 58.520 2867.570 58.580 ;
      LAYER via ;
        RECT 1063.160 375.740 1063.420 376.000 ;
        RECT 1065.460 375.740 1065.720 376.000 ;
        RECT 1063.160 58.520 1063.420 58.780 ;
        RECT 2867.280 58.520 2867.540 58.780 ;
      LAYER met2 ;
        RECT 1066.730 400.250 1067.010 404.000 ;
        RECT 1065.520 400.110 1067.010 400.250 ;
        RECT 1065.520 376.030 1065.660 400.110 ;
        RECT 1066.730 400.000 1067.010 400.110 ;
        RECT 1063.160 375.710 1063.420 376.030 ;
        RECT 1065.460 375.710 1065.720 376.030 ;
        RECT 1063.220 58.810 1063.360 375.710 ;
        RECT 1063.160 58.490 1063.420 58.810 ;
        RECT 2867.280 58.490 2867.540 58.810 ;
        RECT 2867.340 1.770 2867.480 58.490 ;
        RECT 2869.430 1.770 2869.990 2.400 ;
        RECT 2867.340 1.630 2869.990 1.770 ;
        RECT 2869.430 -4.800 2869.990 1.630 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.030 30.840 1070.350 30.900 ;
        RECT 2887.030 30.840 2887.350 30.900 ;
        RECT 1070.030 30.700 2887.350 30.840 ;
        RECT 1070.030 30.640 1070.350 30.700 ;
        RECT 2887.030 30.640 2887.350 30.700 ;
      LAYER via ;
        RECT 1070.060 30.640 1070.320 30.900 ;
        RECT 2887.060 30.640 2887.320 30.900 ;
      LAYER met2 ;
        RECT 1071.790 400.250 1072.070 404.000 ;
        RECT 1070.580 400.110 1072.070 400.250 ;
        RECT 1070.580 398.210 1070.720 400.110 ;
        RECT 1071.790 400.000 1072.070 400.110 ;
        RECT 1070.120 398.070 1070.720 398.210 ;
        RECT 1070.120 30.930 1070.260 398.070 ;
        RECT 1070.060 30.610 1070.320 30.930 ;
        RECT 2887.060 30.610 2887.320 30.930 ;
        RECT 2887.120 2.400 2887.260 30.610 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 40.020 455.790 40.080 ;
        RECT 621.070 40.020 621.390 40.080 ;
        RECT 455.470 39.880 621.390 40.020 ;
        RECT 455.470 39.820 455.790 39.880 ;
        RECT 621.070 39.820 621.390 39.880 ;
        RECT 621.070 19.620 621.390 19.680 ;
        RECT 847.850 19.620 848.170 19.680 ;
        RECT 621.070 19.480 848.170 19.620 ;
        RECT 621.070 19.420 621.390 19.480 ;
        RECT 847.850 19.420 848.170 19.480 ;
      LAYER via ;
        RECT 455.500 39.820 455.760 40.080 ;
        RECT 621.100 39.820 621.360 40.080 ;
        RECT 621.100 19.420 621.360 19.680 ;
        RECT 847.880 19.420 848.140 19.680 ;
      LAYER met2 ;
        RECT 455.850 400.250 456.130 404.000 ;
        RECT 455.560 400.110 456.130 400.250 ;
        RECT 455.560 40.110 455.700 400.110 ;
        RECT 455.850 400.000 456.130 400.110 ;
        RECT 455.500 39.790 455.760 40.110 ;
        RECT 621.100 39.790 621.360 40.110 ;
        RECT 621.160 19.710 621.300 39.790 ;
        RECT 621.100 19.390 621.360 19.710 ;
        RECT 847.880 19.390 848.140 19.710 ;
        RECT 847.940 2.400 848.080 19.390 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 385.800 456.710 385.860 ;
        RECT 460.070 385.800 460.390 385.860 ;
        RECT 456.390 385.660 460.390 385.800 ;
        RECT 456.390 385.600 456.710 385.660 ;
        RECT 460.070 385.600 460.390 385.660 ;
        RECT 456.390 53.280 456.710 53.340 ;
        RECT 863.490 53.280 863.810 53.340 ;
        RECT 456.390 53.140 863.810 53.280 ;
        RECT 456.390 53.080 456.710 53.140 ;
        RECT 863.490 53.080 863.810 53.140 ;
      LAYER via ;
        RECT 456.420 385.600 456.680 385.860 ;
        RECT 460.100 385.600 460.360 385.860 ;
        RECT 456.420 53.080 456.680 53.340 ;
        RECT 863.520 53.080 863.780 53.340 ;
      LAYER met2 ;
        RECT 460.910 400.250 461.190 404.000 ;
        RECT 460.160 400.110 461.190 400.250 ;
        RECT 460.160 385.890 460.300 400.110 ;
        RECT 460.910 400.000 461.190 400.110 ;
        RECT 456.420 385.570 456.680 385.890 ;
        RECT 460.100 385.570 460.360 385.890 ;
        RECT 456.480 53.370 456.620 385.570 ;
        RECT 456.420 53.050 456.680 53.370 ;
        RECT 863.520 53.050 863.780 53.370 ;
        RECT 863.580 1.770 863.720 53.050 ;
        RECT 865.670 1.770 866.230 2.400 ;
        RECT 863.580 1.630 866.230 1.770 ;
        RECT 865.670 -4.800 866.230 1.630 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 387.160 462.690 387.220 ;
        RECT 465.130 387.160 465.450 387.220 ;
        RECT 462.370 387.020 465.450 387.160 ;
        RECT 462.370 386.960 462.690 387.020 ;
        RECT 465.130 386.960 465.450 387.020 ;
        RECT 462.370 52.260 462.690 52.320 ;
        RECT 884.190 52.260 884.510 52.320 ;
        RECT 462.370 52.120 884.510 52.260 ;
        RECT 462.370 52.060 462.690 52.120 ;
        RECT 884.190 52.060 884.510 52.120 ;
      LAYER via ;
        RECT 462.400 386.960 462.660 387.220 ;
        RECT 465.160 386.960 465.420 387.220 ;
        RECT 462.400 52.060 462.660 52.320 ;
        RECT 884.220 52.060 884.480 52.320 ;
      LAYER met2 ;
        RECT 466.430 400.250 466.710 404.000 ;
        RECT 465.220 400.110 466.710 400.250 ;
        RECT 465.220 387.250 465.360 400.110 ;
        RECT 466.430 400.000 466.710 400.110 ;
        RECT 462.400 386.930 462.660 387.250 ;
        RECT 465.160 386.930 465.420 387.250 ;
        RECT 462.460 52.350 462.600 386.930 ;
        RECT 462.400 52.030 462.660 52.350 ;
        RECT 884.220 52.030 884.480 52.350 ;
        RECT 884.280 17.410 884.420 52.030 ;
        RECT 883.360 17.270 884.420 17.410 ;
        RECT 883.360 2.400 883.500 17.270 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.650 51.920 470.970 51.980 ;
        RECT 901.210 51.920 901.530 51.980 ;
        RECT 470.650 51.780 901.530 51.920 ;
        RECT 470.650 51.720 470.970 51.780 ;
        RECT 901.210 51.720 901.530 51.780 ;
      LAYER via ;
        RECT 470.680 51.720 470.940 51.980 ;
        RECT 901.240 51.720 901.500 51.980 ;
      LAYER met2 ;
        RECT 471.950 400.250 472.230 404.000 ;
        RECT 470.740 400.110 472.230 400.250 ;
        RECT 470.740 52.010 470.880 400.110 ;
        RECT 471.950 400.000 472.230 400.110 ;
        RECT 470.680 51.690 470.940 52.010 ;
        RECT 901.240 51.690 901.500 52.010 ;
        RECT 901.300 2.400 901.440 51.690 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 477.090 392.940 477.410 393.000 ;
        RECT 638.090 392.940 638.410 393.000 ;
        RECT 477.090 392.800 638.410 392.940 ;
        RECT 477.090 392.740 477.410 392.800 ;
        RECT 638.090 392.740 638.410 392.800 ;
        RECT 638.090 23.020 638.410 23.080 ;
        RECT 918.690 23.020 919.010 23.080 ;
        RECT 638.090 22.880 919.010 23.020 ;
        RECT 638.090 22.820 638.410 22.880 ;
        RECT 918.690 22.820 919.010 22.880 ;
      LAYER via ;
        RECT 477.120 392.740 477.380 393.000 ;
        RECT 638.120 392.740 638.380 393.000 ;
        RECT 638.120 22.820 638.380 23.080 ;
        RECT 918.720 22.820 918.980 23.080 ;
      LAYER met2 ;
        RECT 477.010 400.180 477.290 404.000 ;
        RECT 477.010 400.000 477.320 400.180 ;
        RECT 477.180 393.030 477.320 400.000 ;
        RECT 477.120 392.710 477.380 393.030 ;
        RECT 638.120 392.710 638.380 393.030 ;
        RECT 638.180 23.110 638.320 392.710 ;
        RECT 638.120 22.790 638.380 23.110 ;
        RECT 918.720 22.790 918.980 23.110 ;
        RECT 918.780 2.400 918.920 22.790 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 482.610 392.260 482.930 392.320 ;
        RECT 658.790 392.260 659.110 392.320 ;
        RECT 482.610 392.120 659.110 392.260 ;
        RECT 482.610 392.060 482.930 392.120 ;
        RECT 658.790 392.060 659.110 392.120 ;
        RECT 658.790 22.340 659.110 22.400 ;
        RECT 936.630 22.340 936.950 22.400 ;
        RECT 658.790 22.200 936.950 22.340 ;
        RECT 658.790 22.140 659.110 22.200 ;
        RECT 936.630 22.140 936.950 22.200 ;
      LAYER via ;
        RECT 482.640 392.060 482.900 392.320 ;
        RECT 658.820 392.060 659.080 392.320 ;
        RECT 658.820 22.140 659.080 22.400 ;
        RECT 936.660 22.140 936.920 22.400 ;
      LAYER met2 ;
        RECT 482.530 400.180 482.810 404.000 ;
        RECT 482.530 400.000 482.840 400.180 ;
        RECT 482.700 392.350 482.840 400.000 ;
        RECT 482.640 392.030 482.900 392.350 ;
        RECT 658.820 392.030 659.080 392.350 ;
        RECT 658.880 22.430 659.020 392.030 ;
        RECT 658.820 22.110 659.080 22.430 ;
        RECT 936.660 22.110 936.920 22.430 ;
        RECT 936.720 2.400 936.860 22.110 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 488.130 391.920 488.450 391.980 ;
        RECT 665.690 391.920 666.010 391.980 ;
        RECT 488.130 391.780 666.010 391.920 ;
        RECT 488.130 391.720 488.450 391.780 ;
        RECT 665.690 391.720 666.010 391.780 ;
        RECT 665.690 23.360 666.010 23.420 ;
        RECT 954.110 23.360 954.430 23.420 ;
        RECT 665.690 23.220 954.430 23.360 ;
        RECT 665.690 23.160 666.010 23.220 ;
        RECT 954.110 23.160 954.430 23.220 ;
      LAYER via ;
        RECT 488.160 391.720 488.420 391.980 ;
        RECT 665.720 391.720 665.980 391.980 ;
        RECT 665.720 23.160 665.980 23.420 ;
        RECT 954.140 23.160 954.400 23.420 ;
      LAYER met2 ;
        RECT 488.050 400.180 488.330 404.000 ;
        RECT 488.050 400.000 488.360 400.180 ;
        RECT 488.220 392.010 488.360 400.000 ;
        RECT 488.160 391.690 488.420 392.010 ;
        RECT 665.720 391.690 665.980 392.010 ;
        RECT 665.780 23.450 665.920 391.690 ;
        RECT 665.720 23.130 665.980 23.450 ;
        RECT 954.140 23.130 954.400 23.450 ;
        RECT 954.200 2.400 954.340 23.130 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.730 391.580 493.050 391.640 ;
        RECT 693.290 391.580 693.610 391.640 ;
        RECT 492.730 391.440 693.610 391.580 ;
        RECT 492.730 391.380 493.050 391.440 ;
        RECT 693.290 391.380 693.610 391.440 ;
        RECT 693.290 21.320 693.610 21.380 ;
        RECT 972.050 21.320 972.370 21.380 ;
        RECT 693.290 21.180 972.370 21.320 ;
        RECT 693.290 21.120 693.610 21.180 ;
        RECT 972.050 21.120 972.370 21.180 ;
      LAYER via ;
        RECT 492.760 391.380 493.020 391.640 ;
        RECT 693.320 391.380 693.580 391.640 ;
        RECT 693.320 21.120 693.580 21.380 ;
        RECT 972.080 21.120 972.340 21.380 ;
      LAYER met2 ;
        RECT 493.110 400.250 493.390 404.000 ;
        RECT 492.820 400.110 493.390 400.250 ;
        RECT 492.820 391.670 492.960 400.110 ;
        RECT 493.110 400.000 493.390 400.110 ;
        RECT 492.760 391.350 493.020 391.670 ;
        RECT 693.320 391.350 693.580 391.670 ;
        RECT 693.380 21.410 693.520 391.350 ;
        RECT 693.320 21.090 693.580 21.410 ;
        RECT 972.080 21.090 972.340 21.410 ;
        RECT 972.140 2.400 972.280 21.090 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.750 393.620 395.070 393.680 ;
        RECT 397.050 393.620 397.370 393.680 ;
        RECT 394.750 393.480 397.370 393.620 ;
        RECT 394.750 393.420 395.070 393.480 ;
        RECT 397.050 393.420 397.370 393.480 ;
        RECT 394.750 39.000 395.070 39.060 ;
        RECT 652.810 39.000 653.130 39.060 ;
        RECT 394.750 38.860 653.130 39.000 ;
        RECT 394.750 38.800 395.070 38.860 ;
        RECT 652.810 38.800 653.130 38.860 ;
      LAYER via ;
        RECT 394.780 393.420 395.040 393.680 ;
        RECT 397.080 393.420 397.340 393.680 ;
        RECT 394.780 38.800 395.040 39.060 ;
        RECT 652.840 38.800 653.100 39.060 ;
      LAYER met2 ;
        RECT 396.970 400.180 397.250 404.000 ;
        RECT 396.970 400.000 397.280 400.180 ;
        RECT 397.140 393.710 397.280 400.000 ;
        RECT 394.780 393.390 395.040 393.710 ;
        RECT 397.080 393.390 397.340 393.710 ;
        RECT 394.840 39.090 394.980 393.390 ;
        RECT 394.780 38.770 395.040 39.090 ;
        RECT 652.840 38.770 653.100 39.090 ;
        RECT 652.900 2.400 653.040 38.770 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.790 59.740 498.110 59.800 ;
        RECT 989.530 59.740 989.850 59.800 ;
        RECT 497.790 59.600 989.850 59.740 ;
        RECT 497.790 59.540 498.110 59.600 ;
        RECT 989.530 59.540 989.850 59.600 ;
      LAYER via ;
        RECT 497.820 59.540 498.080 59.800 ;
        RECT 989.560 59.540 989.820 59.800 ;
      LAYER met2 ;
        RECT 498.630 400.250 498.910 404.000 ;
        RECT 497.880 400.110 498.910 400.250 ;
        RECT 497.880 59.830 498.020 400.110 ;
        RECT 498.630 400.000 498.910 400.110 ;
        RECT 497.820 59.510 498.080 59.830 ;
        RECT 989.560 59.510 989.820 59.830 ;
        RECT 989.620 2.400 989.760 59.510 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 391.240 504.550 391.300 ;
        RECT 713.990 391.240 714.310 391.300 ;
        RECT 504.230 391.100 714.310 391.240 ;
        RECT 504.230 391.040 504.550 391.100 ;
        RECT 713.990 391.040 714.310 391.100 ;
        RECT 713.990 22.000 714.310 22.060 ;
        RECT 1007.470 22.000 1007.790 22.060 ;
        RECT 713.990 21.860 1007.790 22.000 ;
        RECT 713.990 21.800 714.310 21.860 ;
        RECT 1007.470 21.800 1007.790 21.860 ;
      LAYER via ;
        RECT 504.260 391.040 504.520 391.300 ;
        RECT 714.020 391.040 714.280 391.300 ;
        RECT 714.020 21.800 714.280 22.060 ;
        RECT 1007.500 21.800 1007.760 22.060 ;
      LAYER met2 ;
        RECT 504.150 400.180 504.430 404.000 ;
        RECT 504.150 400.000 504.460 400.180 ;
        RECT 504.320 391.330 504.460 400.000 ;
        RECT 504.260 391.010 504.520 391.330 ;
        RECT 714.020 391.010 714.280 391.330 ;
        RECT 714.080 22.090 714.220 391.010 ;
        RECT 714.020 21.770 714.280 22.090 ;
        RECT 1007.500 21.770 1007.760 22.090 ;
        RECT 1007.560 2.400 1007.700 21.770 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 509.290 390.900 509.610 390.960 ;
        RECT 727.330 390.900 727.650 390.960 ;
        RECT 509.290 390.760 727.650 390.900 ;
        RECT 509.290 390.700 509.610 390.760 ;
        RECT 727.330 390.700 727.650 390.760 ;
        RECT 727.790 21.660 728.110 21.720 ;
        RECT 1025.410 21.660 1025.730 21.720 ;
        RECT 727.790 21.520 1025.730 21.660 ;
        RECT 727.790 21.460 728.110 21.520 ;
        RECT 1025.410 21.460 1025.730 21.520 ;
      LAYER via ;
        RECT 509.320 390.700 509.580 390.960 ;
        RECT 727.360 390.700 727.620 390.960 ;
        RECT 727.820 21.460 728.080 21.720 ;
        RECT 1025.440 21.460 1025.700 21.720 ;
      LAYER met2 ;
        RECT 509.210 400.180 509.490 404.000 ;
        RECT 509.210 400.000 509.520 400.180 ;
        RECT 509.380 390.990 509.520 400.000 ;
        RECT 509.320 390.670 509.580 390.990 ;
        RECT 727.360 390.670 727.620 390.990 ;
        RECT 727.420 372.670 727.560 390.670 ;
        RECT 727.420 372.530 728.020 372.670 ;
        RECT 727.880 21.750 728.020 372.530 ;
        RECT 727.820 21.430 728.080 21.750 ;
        RECT 1025.440 21.430 1025.700 21.750 ;
        RECT 1025.500 2.400 1025.640 21.430 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 386.820 511.450 386.880 ;
        RECT 513.430 386.820 513.750 386.880 ;
        RECT 511.130 386.680 513.750 386.820 ;
        RECT 511.130 386.620 511.450 386.680 ;
        RECT 513.430 386.620 513.750 386.680 ;
        RECT 511.130 49.880 511.450 49.940 ;
        RECT 1042.890 49.880 1043.210 49.940 ;
        RECT 511.130 49.740 1043.210 49.880 ;
        RECT 511.130 49.680 511.450 49.740 ;
        RECT 1042.890 49.680 1043.210 49.740 ;
      LAYER via ;
        RECT 511.160 386.620 511.420 386.880 ;
        RECT 513.460 386.620 513.720 386.880 ;
        RECT 511.160 49.680 511.420 49.940 ;
        RECT 1042.920 49.680 1043.180 49.940 ;
      LAYER met2 ;
        RECT 514.730 400.250 515.010 404.000 ;
        RECT 513.520 400.110 515.010 400.250 ;
        RECT 513.520 386.910 513.660 400.110 ;
        RECT 514.730 400.000 515.010 400.110 ;
        RECT 511.160 386.590 511.420 386.910 ;
        RECT 513.460 386.590 513.720 386.910 ;
        RECT 511.220 49.970 511.360 386.590 ;
        RECT 511.160 49.650 511.420 49.970 ;
        RECT 1042.920 49.650 1043.180 49.970 ;
        RECT 1042.980 2.400 1043.120 49.650 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 520.330 390.220 520.650 390.280 ;
        RECT 782.990 390.220 783.310 390.280 ;
        RECT 520.330 390.080 783.310 390.220 ;
        RECT 520.330 390.020 520.650 390.080 ;
        RECT 782.990 390.020 783.310 390.080 ;
        RECT 782.990 28.800 783.310 28.860 ;
        RECT 1060.830 28.800 1061.150 28.860 ;
        RECT 782.990 28.660 1061.150 28.800 ;
        RECT 782.990 28.600 783.310 28.660 ;
        RECT 1060.830 28.600 1061.150 28.660 ;
      LAYER via ;
        RECT 520.360 390.020 520.620 390.280 ;
        RECT 783.020 390.020 783.280 390.280 ;
        RECT 783.020 28.600 783.280 28.860 ;
        RECT 1060.860 28.600 1061.120 28.860 ;
      LAYER met2 ;
        RECT 520.250 400.180 520.530 404.000 ;
        RECT 520.250 400.000 520.560 400.180 ;
        RECT 520.420 390.310 520.560 400.000 ;
        RECT 520.360 389.990 520.620 390.310 ;
        RECT 783.020 389.990 783.280 390.310 ;
        RECT 783.080 28.890 783.220 389.990 ;
        RECT 783.020 28.570 783.280 28.890 ;
        RECT 1060.860 28.570 1061.120 28.890 ;
        RECT 1060.920 2.400 1061.060 28.570 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 57.020 524.790 57.080 ;
        RECT 1076.930 57.020 1077.250 57.080 ;
        RECT 524.470 56.880 1077.250 57.020 ;
        RECT 524.470 56.820 524.790 56.880 ;
        RECT 1076.930 56.820 1077.250 56.880 ;
      LAYER via ;
        RECT 524.500 56.820 524.760 57.080 ;
        RECT 1076.960 56.820 1077.220 57.080 ;
      LAYER met2 ;
        RECT 525.310 400.250 525.590 404.000 ;
        RECT 524.560 400.110 525.590 400.250 ;
        RECT 524.560 57.110 524.700 400.110 ;
        RECT 525.310 400.000 525.590 400.110 ;
        RECT 524.500 56.790 524.760 57.110 ;
        RECT 1076.960 56.790 1077.220 57.110 ;
        RECT 1077.020 1.770 1077.160 56.790 ;
        RECT 1078.190 1.770 1078.750 2.400 ;
        RECT 1077.020 1.630 1078.750 1.770 ;
        RECT 1078.190 -4.800 1078.750 1.630 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.390 385.800 525.710 385.860 ;
        RECT 529.530 385.800 529.850 385.860 ;
        RECT 525.390 385.660 529.850 385.800 ;
        RECT 525.390 385.600 525.710 385.660 ;
        RECT 529.530 385.600 529.850 385.660 ;
        RECT 525.390 112.100 525.710 112.160 ;
        RECT 1090.270 112.100 1090.590 112.160 ;
        RECT 525.390 111.960 1090.590 112.100 ;
        RECT 525.390 111.900 525.710 111.960 ;
        RECT 1090.270 111.900 1090.590 111.960 ;
        RECT 1090.270 15.200 1090.590 15.260 ;
        RECT 1096.250 15.200 1096.570 15.260 ;
        RECT 1090.270 15.060 1096.570 15.200 ;
        RECT 1090.270 15.000 1090.590 15.060 ;
        RECT 1096.250 15.000 1096.570 15.060 ;
      LAYER via ;
        RECT 525.420 385.600 525.680 385.860 ;
        RECT 529.560 385.600 529.820 385.860 ;
        RECT 525.420 111.900 525.680 112.160 ;
        RECT 1090.300 111.900 1090.560 112.160 ;
        RECT 1090.300 15.000 1090.560 15.260 ;
        RECT 1096.280 15.000 1096.540 15.260 ;
      LAYER met2 ;
        RECT 530.830 400.250 531.110 404.000 ;
        RECT 529.620 400.110 531.110 400.250 ;
        RECT 529.620 385.890 529.760 400.110 ;
        RECT 530.830 400.000 531.110 400.110 ;
        RECT 525.420 385.570 525.680 385.890 ;
        RECT 529.560 385.570 529.820 385.890 ;
        RECT 525.480 112.190 525.620 385.570 ;
        RECT 525.420 111.870 525.680 112.190 ;
        RECT 1090.300 111.870 1090.560 112.190 ;
        RECT 1090.360 15.290 1090.500 111.870 ;
        RECT 1090.300 14.970 1090.560 15.290 ;
        RECT 1096.280 14.970 1096.540 15.290 ;
        RECT 1096.340 2.400 1096.480 14.970 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.290 112.440 532.610 112.500 ;
        RECT 1110.970 112.440 1111.290 112.500 ;
        RECT 532.290 112.300 1111.290 112.440 ;
        RECT 532.290 112.240 532.610 112.300 ;
        RECT 1110.970 112.240 1111.290 112.300 ;
      LAYER via ;
        RECT 532.320 112.240 532.580 112.500 ;
        RECT 1111.000 112.240 1111.260 112.500 ;
      LAYER met2 ;
        RECT 535.890 400.250 536.170 404.000 ;
        RECT 535.140 400.110 536.170 400.250 ;
        RECT 535.140 386.480 535.280 400.110 ;
        RECT 535.890 400.000 536.170 400.110 ;
        RECT 532.380 386.340 535.280 386.480 ;
        RECT 532.380 112.530 532.520 386.340 ;
        RECT 532.320 112.210 532.580 112.530 ;
        RECT 1111.000 112.210 1111.260 112.530 ;
        RECT 1111.060 82.870 1111.200 112.210 ;
        RECT 1111.060 82.730 1113.960 82.870 ;
        RECT 1113.820 2.400 1113.960 82.730 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.190 112.780 539.510 112.840 ;
        RECT 1131.670 112.780 1131.990 112.840 ;
        RECT 539.190 112.640 1131.990 112.780 ;
        RECT 539.190 112.580 539.510 112.640 ;
        RECT 1131.670 112.580 1131.990 112.640 ;
      LAYER via ;
        RECT 539.220 112.580 539.480 112.840 ;
        RECT 1131.700 112.580 1131.960 112.840 ;
      LAYER met2 ;
        RECT 541.410 400.250 541.690 404.000 ;
        RECT 540.200 400.110 541.690 400.250 ;
        RECT 540.200 324.370 540.340 400.110 ;
        RECT 541.410 400.000 541.690 400.110 ;
        RECT 539.280 324.230 540.340 324.370 ;
        RECT 539.280 112.870 539.420 324.230 ;
        RECT 539.220 112.550 539.480 112.870 ;
        RECT 1131.700 112.550 1131.960 112.870 ;
        RECT 1131.760 2.400 1131.900 112.550 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.550 113.120 546.870 113.180 ;
        RECT 1145.470 113.120 1145.790 113.180 ;
        RECT 546.550 112.980 1145.790 113.120 ;
        RECT 546.550 112.920 546.870 112.980 ;
        RECT 1145.470 112.920 1145.790 112.980 ;
      LAYER via ;
        RECT 546.580 112.920 546.840 113.180 ;
        RECT 1145.500 112.920 1145.760 113.180 ;
      LAYER met2 ;
        RECT 546.930 400.250 547.210 404.000 ;
        RECT 546.640 400.110 547.210 400.250 ;
        RECT 546.640 113.210 546.780 400.110 ;
        RECT 546.930 400.000 547.210 400.110 ;
        RECT 546.580 112.890 546.840 113.210 ;
        RECT 1145.500 112.890 1145.760 113.210 ;
        RECT 1145.560 82.870 1145.700 112.890 ;
        RECT 1145.560 82.730 1147.080 82.870 ;
        RECT 1146.940 1.770 1147.080 82.730 ;
        RECT 1149.030 1.770 1149.590 2.400 ;
        RECT 1146.940 1.630 1149.590 1.770 ;
        RECT 1149.030 -4.800 1149.590 1.630 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 401.650 38.320 401.970 38.380 ;
        RECT 670.750 38.320 671.070 38.380 ;
        RECT 401.650 38.180 671.070 38.320 ;
        RECT 401.650 38.120 401.970 38.180 ;
        RECT 670.750 38.120 671.070 38.180 ;
      LAYER via ;
        RECT 401.680 38.120 401.940 38.380 ;
        RECT 670.780 38.120 671.040 38.380 ;
      LAYER met2 ;
        RECT 402.030 400.250 402.310 404.000 ;
        RECT 401.740 400.110 402.310 400.250 ;
        RECT 401.740 38.410 401.880 400.110 ;
        RECT 402.030 400.000 402.310 400.110 ;
        RECT 401.680 38.090 401.940 38.410 ;
        RECT 670.780 38.090 671.040 38.410 ;
        RECT 670.840 2.400 670.980 38.090 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.450 113.460 553.770 113.520 ;
        RECT 1166.170 113.460 1166.490 113.520 ;
        RECT 553.450 113.320 1166.490 113.460 ;
        RECT 553.450 113.260 553.770 113.320 ;
        RECT 1166.170 113.260 1166.490 113.320 ;
      LAYER via ;
        RECT 553.480 113.260 553.740 113.520 ;
        RECT 1166.200 113.260 1166.460 113.520 ;
      LAYER met2 ;
        RECT 551.990 400.250 552.270 404.000 ;
        RECT 551.990 400.110 552.760 400.250 ;
        RECT 551.990 400.000 552.270 400.110 ;
        RECT 552.620 399.570 552.760 400.110 ;
        RECT 552.620 399.430 553.680 399.570 ;
        RECT 553.540 113.550 553.680 399.430 ;
        RECT 553.480 113.230 553.740 113.550 ;
        RECT 1166.200 113.230 1166.460 113.550 ;
        RECT 1166.260 82.870 1166.400 113.230 ;
        RECT 1166.260 82.730 1167.320 82.870 ;
        RECT 1167.180 2.400 1167.320 82.730 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.530 376.280 552.850 376.340 ;
        RECT 556.210 376.280 556.530 376.340 ;
        RECT 552.530 376.140 556.530 376.280 ;
        RECT 552.530 376.080 552.850 376.140 ;
        RECT 556.210 376.080 556.530 376.140 ;
        RECT 552.530 63.820 552.850 63.880 ;
        RECT 1182.730 63.820 1183.050 63.880 ;
        RECT 552.530 63.680 1183.050 63.820 ;
        RECT 552.530 63.620 552.850 63.680 ;
        RECT 1182.730 63.620 1183.050 63.680 ;
      LAYER via ;
        RECT 552.560 376.080 552.820 376.340 ;
        RECT 556.240 376.080 556.500 376.340 ;
        RECT 552.560 63.620 552.820 63.880 ;
        RECT 1182.760 63.620 1183.020 63.880 ;
      LAYER met2 ;
        RECT 557.510 400.250 557.790 404.000 ;
        RECT 556.300 400.110 557.790 400.250 ;
        RECT 556.300 376.370 556.440 400.110 ;
        RECT 557.510 400.000 557.790 400.110 ;
        RECT 552.560 376.050 552.820 376.370 ;
        RECT 556.240 376.050 556.500 376.370 ;
        RECT 552.620 63.910 552.760 376.050 ;
        RECT 552.560 63.590 552.820 63.910 ;
        RECT 1182.760 63.590 1183.020 63.910 ;
        RECT 1182.820 1.770 1182.960 63.590 ;
        RECT 1184.910 1.770 1185.470 2.400 ;
        RECT 1182.820 1.630 1185.470 1.770 ;
        RECT 1184.910 -4.800 1185.470 1.630 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 377.300 559.750 377.360 ;
        RECT 561.730 377.300 562.050 377.360 ;
        RECT 559.430 377.160 562.050 377.300 ;
        RECT 559.430 377.100 559.750 377.160 ;
        RECT 561.730 377.100 562.050 377.160 ;
        RECT 559.430 64.160 559.750 64.220 ;
        RECT 1200.670 64.160 1200.990 64.220 ;
        RECT 559.430 64.020 1200.990 64.160 ;
        RECT 559.430 63.960 559.750 64.020 ;
        RECT 1200.670 63.960 1200.990 64.020 ;
      LAYER via ;
        RECT 559.460 377.100 559.720 377.360 ;
        RECT 561.760 377.100 562.020 377.360 ;
        RECT 559.460 63.960 559.720 64.220 ;
        RECT 1200.700 63.960 1200.960 64.220 ;
      LAYER met2 ;
        RECT 563.030 400.250 563.310 404.000 ;
        RECT 561.820 400.110 563.310 400.250 ;
        RECT 561.820 377.390 561.960 400.110 ;
        RECT 563.030 400.000 563.310 400.110 ;
        RECT 559.460 377.070 559.720 377.390 ;
        RECT 561.760 377.070 562.020 377.390 ;
        RECT 559.520 64.250 559.660 377.070 ;
        RECT 559.460 63.930 559.720 64.250 ;
        RECT 1200.700 63.930 1200.960 64.250 ;
        RECT 1200.760 1.770 1200.900 63.930 ;
        RECT 1202.390 1.770 1202.950 2.400 ;
        RECT 1200.760 1.630 1202.950 1.770 ;
        RECT 1202.390 -4.800 1202.950 1.630 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 64.500 567.110 64.560 ;
        RECT 1214.470 64.500 1214.790 64.560 ;
        RECT 566.790 64.360 1214.790 64.500 ;
        RECT 566.790 64.300 567.110 64.360 ;
        RECT 1214.470 64.300 1214.790 64.360 ;
        RECT 1214.470 15.200 1214.790 15.260 ;
        RECT 1220.450 15.200 1220.770 15.260 ;
        RECT 1214.470 15.060 1220.770 15.200 ;
        RECT 1214.470 15.000 1214.790 15.060 ;
        RECT 1220.450 15.000 1220.770 15.060 ;
      LAYER via ;
        RECT 566.820 64.300 567.080 64.560 ;
        RECT 1214.500 64.300 1214.760 64.560 ;
        RECT 1214.500 15.000 1214.760 15.260 ;
        RECT 1220.480 15.000 1220.740 15.260 ;
      LAYER met2 ;
        RECT 568.090 400.250 568.370 404.000 ;
        RECT 567.340 400.110 568.370 400.250 ;
        RECT 567.340 351.970 567.480 400.110 ;
        RECT 568.090 400.000 568.370 400.110 ;
        RECT 566.880 351.830 567.480 351.970 ;
        RECT 566.880 64.590 567.020 351.830 ;
        RECT 566.820 64.270 567.080 64.590 ;
        RECT 1214.500 64.270 1214.760 64.590 ;
        RECT 1214.560 15.290 1214.700 64.270 ;
        RECT 1214.500 14.970 1214.760 15.290 ;
        RECT 1220.480 14.970 1220.740 15.290 ;
        RECT 1220.540 2.400 1220.680 14.970 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.230 64.840 573.550 64.900 ;
        RECT 1237.930 64.840 1238.250 64.900 ;
        RECT 573.230 64.700 1238.250 64.840 ;
        RECT 573.230 64.640 573.550 64.700 ;
        RECT 1237.930 64.640 1238.250 64.700 ;
      LAYER via ;
        RECT 573.260 64.640 573.520 64.900 ;
        RECT 1237.960 64.640 1238.220 64.900 ;
      LAYER met2 ;
        RECT 573.610 400.250 573.890 404.000 ;
        RECT 573.320 400.110 573.890 400.250 ;
        RECT 573.320 64.930 573.460 400.110 ;
        RECT 573.610 400.000 573.890 400.110 ;
        RECT 573.260 64.610 573.520 64.930 ;
        RECT 1237.960 64.610 1238.220 64.930 ;
        RECT 1238.020 2.400 1238.160 64.610 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.690 376.280 574.010 376.340 ;
        RECT 577.830 376.280 578.150 376.340 ;
        RECT 573.690 376.140 578.150 376.280 ;
        RECT 573.690 376.080 574.010 376.140 ;
        RECT 577.830 376.080 578.150 376.140 ;
        RECT 573.690 65.180 574.010 65.240 ;
        RECT 1256.330 65.180 1256.650 65.240 ;
        RECT 573.690 65.040 1256.650 65.180 ;
        RECT 573.690 64.980 574.010 65.040 ;
        RECT 1256.330 64.980 1256.650 65.040 ;
      LAYER via ;
        RECT 573.720 376.080 573.980 376.340 ;
        RECT 577.860 376.080 578.120 376.340 ;
        RECT 573.720 64.980 573.980 65.240 ;
        RECT 1256.360 64.980 1256.620 65.240 ;
      LAYER met2 ;
        RECT 579.130 400.250 579.410 404.000 ;
        RECT 577.920 400.110 579.410 400.250 ;
        RECT 577.920 376.370 578.060 400.110 ;
        RECT 579.130 400.000 579.410 400.110 ;
        RECT 573.720 376.050 573.980 376.370 ;
        RECT 577.860 376.050 578.120 376.370 ;
        RECT 573.780 65.270 573.920 376.050 ;
        RECT 573.720 64.950 573.980 65.270 ;
        RECT 1256.360 64.950 1256.620 65.270 ;
        RECT 1256.420 17.410 1256.560 64.950 ;
        RECT 1255.960 17.270 1256.560 17.410 ;
        RECT 1255.960 2.400 1256.100 17.270 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.130 399.740 580.450 399.800 ;
        RECT 582.890 399.740 583.210 399.800 ;
        RECT 580.130 399.600 583.210 399.740 ;
        RECT 580.130 399.540 580.450 399.600 ;
        RECT 582.890 399.540 583.210 399.600 ;
        RECT 580.130 68.920 580.450 68.980 ;
        RECT 1271.050 68.920 1271.370 68.980 ;
        RECT 580.130 68.780 1271.370 68.920 ;
        RECT 580.130 68.720 580.450 68.780 ;
        RECT 1271.050 68.720 1271.370 68.780 ;
      LAYER via ;
        RECT 580.160 399.540 580.420 399.800 ;
        RECT 582.920 399.540 583.180 399.800 ;
        RECT 580.160 68.720 580.420 68.980 ;
        RECT 1271.080 68.720 1271.340 68.980 ;
      LAYER met2 ;
        RECT 584.190 400.250 584.470 404.000 ;
        RECT 582.980 400.110 584.470 400.250 ;
        RECT 582.980 399.830 583.120 400.110 ;
        RECT 584.190 400.000 584.470 400.110 ;
        RECT 580.160 399.510 580.420 399.830 ;
        RECT 582.920 399.510 583.180 399.830 ;
        RECT 580.220 69.010 580.360 399.510 ;
        RECT 580.160 68.690 580.420 69.010 ;
        RECT 1271.080 68.690 1271.340 69.010 ;
        RECT 1271.140 1.770 1271.280 68.690 ;
        RECT 1273.230 1.770 1273.790 2.400 ;
        RECT 1271.140 1.630 1273.790 1.770 ;
        RECT 1273.230 -4.800 1273.790 1.630 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.030 68.580 587.350 68.640 ;
        RECT 1291.290 68.580 1291.610 68.640 ;
        RECT 587.030 68.440 1291.610 68.580 ;
        RECT 587.030 68.380 587.350 68.440 ;
        RECT 1291.290 68.380 1291.610 68.440 ;
      LAYER via ;
        RECT 587.060 68.380 587.320 68.640 ;
        RECT 1291.320 68.380 1291.580 68.640 ;
      LAYER met2 ;
        RECT 589.710 400.250 589.990 404.000 ;
        RECT 588.500 400.110 589.990 400.250 ;
        RECT 588.500 399.570 588.640 400.110 ;
        RECT 589.710 400.000 589.990 400.110 ;
        RECT 587.120 399.430 588.640 399.570 ;
        RECT 587.120 68.670 587.260 399.430 ;
        RECT 587.060 68.350 587.320 68.670 ;
        RECT 1291.320 68.350 1291.580 68.670 ;
        RECT 1291.380 2.400 1291.520 68.350 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.930 68.240 594.250 68.300 ;
        RECT 1308.770 68.240 1309.090 68.300 ;
        RECT 593.930 68.100 1309.090 68.240 ;
        RECT 593.930 68.040 594.250 68.100 ;
        RECT 1308.770 68.040 1309.090 68.100 ;
      LAYER via ;
        RECT 593.960 68.040 594.220 68.300 ;
        RECT 1308.800 68.040 1309.060 68.300 ;
      LAYER met2 ;
        RECT 595.230 400.250 595.510 404.000 ;
        RECT 594.020 400.110 595.510 400.250 ;
        RECT 594.020 68.330 594.160 400.110 ;
        RECT 595.230 400.000 595.510 400.110 ;
        RECT 593.960 68.010 594.220 68.330 ;
        RECT 1308.800 68.010 1309.060 68.330 ;
        RECT 1308.860 2.400 1309.000 68.010 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 67.900 600.690 67.960 ;
        RECT 1324.870 67.900 1325.190 67.960 ;
        RECT 600.370 67.760 1325.190 67.900 ;
        RECT 600.370 67.700 600.690 67.760 ;
        RECT 1324.870 67.700 1325.190 67.760 ;
      LAYER via ;
        RECT 600.400 67.700 600.660 67.960 ;
        RECT 1324.900 67.700 1325.160 67.960 ;
      LAYER met2 ;
        RECT 600.290 400.180 600.570 404.000 ;
        RECT 600.290 400.000 600.600 400.180 ;
        RECT 600.460 67.990 600.600 400.000 ;
        RECT 600.400 67.670 600.660 67.990 ;
        RECT 1324.900 67.670 1325.160 67.990 ;
        RECT 1324.960 1.770 1325.100 67.670 ;
        RECT 1326.590 1.770 1327.150 2.400 ;
        RECT 1324.960 1.630 1327.150 1.770 ;
        RECT 1326.590 -4.800 1327.150 1.630 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 386.480 407.490 386.540 ;
        RECT 408.550 386.480 408.870 386.540 ;
        RECT 407.170 386.340 408.870 386.480 ;
        RECT 407.170 386.280 407.490 386.340 ;
        RECT 408.550 386.280 408.870 386.340 ;
        RECT 408.550 37.980 408.870 38.040 ;
        RECT 688.230 37.980 688.550 38.040 ;
        RECT 408.550 37.840 688.550 37.980 ;
        RECT 408.550 37.780 408.870 37.840 ;
        RECT 688.230 37.780 688.550 37.840 ;
      LAYER via ;
        RECT 407.200 386.280 407.460 386.540 ;
        RECT 408.580 386.280 408.840 386.540 ;
        RECT 408.580 37.780 408.840 38.040 ;
        RECT 688.260 37.780 688.520 38.040 ;
      LAYER met2 ;
        RECT 407.550 400.250 407.830 404.000 ;
        RECT 407.260 400.110 407.830 400.250 ;
        RECT 407.260 386.570 407.400 400.110 ;
        RECT 407.550 400.000 407.830 400.110 ;
        RECT 407.200 386.250 407.460 386.570 ;
        RECT 408.580 386.250 408.840 386.570 ;
        RECT 408.640 38.070 408.780 386.250 ;
        RECT 408.580 37.750 408.840 38.070 ;
        RECT 688.260 37.750 688.520 38.070 ;
        RECT 688.320 2.400 688.460 37.750 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.830 376.280 601.150 376.340 ;
        RECT 604.510 376.280 604.830 376.340 ;
        RECT 600.830 376.140 604.830 376.280 ;
        RECT 600.830 376.080 601.150 376.140 ;
        RECT 604.510 376.080 604.830 376.140 ;
        RECT 600.830 67.560 601.150 67.620 ;
        RECT 1341.890 67.560 1342.210 67.620 ;
        RECT 600.830 67.420 1342.210 67.560 ;
        RECT 600.830 67.360 601.150 67.420 ;
        RECT 1341.890 67.360 1342.210 67.420 ;
      LAYER via ;
        RECT 600.860 376.080 601.120 376.340 ;
        RECT 604.540 376.080 604.800 376.340 ;
        RECT 600.860 67.360 601.120 67.620 ;
        RECT 1341.920 67.360 1342.180 67.620 ;
      LAYER met2 ;
        RECT 605.810 400.250 606.090 404.000 ;
        RECT 604.600 400.110 606.090 400.250 ;
        RECT 604.600 376.370 604.740 400.110 ;
        RECT 605.810 400.000 606.090 400.110 ;
        RECT 600.860 376.050 601.120 376.370 ;
        RECT 604.540 376.050 604.800 376.370 ;
        RECT 600.920 67.650 601.060 376.050 ;
        RECT 600.860 67.330 601.120 67.650 ;
        RECT 1341.920 67.330 1342.180 67.650 ;
        RECT 1341.980 1.770 1342.120 67.330 ;
        RECT 1344.070 1.770 1344.630 2.400 ;
        RECT 1341.980 1.630 1344.630 1.770 ;
        RECT 1344.070 -4.800 1344.630 1.630 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.270 376.280 607.590 376.340 ;
        RECT 610.030 376.280 610.350 376.340 ;
        RECT 607.270 376.140 610.350 376.280 ;
        RECT 607.270 376.080 607.590 376.140 ;
        RECT 610.030 376.080 610.350 376.140 ;
        RECT 607.270 67.220 607.590 67.280 ;
        RECT 1362.130 67.220 1362.450 67.280 ;
        RECT 607.270 67.080 1362.450 67.220 ;
        RECT 607.270 67.020 607.590 67.080 ;
        RECT 1362.130 67.020 1362.450 67.080 ;
      LAYER via ;
        RECT 607.300 376.080 607.560 376.340 ;
        RECT 610.060 376.080 610.320 376.340 ;
        RECT 607.300 67.020 607.560 67.280 ;
        RECT 1362.160 67.020 1362.420 67.280 ;
      LAYER met2 ;
        RECT 611.330 400.250 611.610 404.000 ;
        RECT 610.120 400.110 611.610 400.250 ;
        RECT 610.120 376.370 610.260 400.110 ;
        RECT 611.330 400.000 611.610 400.110 ;
        RECT 607.300 376.050 607.560 376.370 ;
        RECT 610.060 376.050 610.320 376.370 ;
        RECT 607.360 67.310 607.500 376.050 ;
        RECT 607.300 66.990 607.560 67.310 ;
        RECT 1362.160 66.990 1362.420 67.310 ;
        RECT 1362.220 2.400 1362.360 66.990 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 379.680 614.490 379.740 ;
        RECT 616.470 379.680 616.790 379.740 ;
        RECT 614.170 379.540 616.790 379.680 ;
        RECT 614.170 379.480 614.490 379.540 ;
        RECT 616.470 379.480 616.790 379.540 ;
        RECT 614.170 66.880 614.490 66.940 ;
        RECT 1380.530 66.880 1380.850 66.940 ;
        RECT 614.170 66.740 1380.850 66.880 ;
        RECT 614.170 66.680 614.490 66.740 ;
        RECT 1380.530 66.680 1380.850 66.740 ;
      LAYER via ;
        RECT 614.200 379.480 614.460 379.740 ;
        RECT 616.500 379.480 616.760 379.740 ;
        RECT 614.200 66.680 614.460 66.940 ;
        RECT 1380.560 66.680 1380.820 66.940 ;
      LAYER met2 ;
        RECT 616.390 400.180 616.670 404.000 ;
        RECT 616.390 400.000 616.700 400.180 ;
        RECT 616.560 379.770 616.700 400.000 ;
        RECT 614.200 379.450 614.460 379.770 ;
        RECT 616.500 379.450 616.760 379.770 ;
        RECT 614.260 66.970 614.400 379.450 ;
        RECT 614.200 66.650 614.460 66.970 ;
        RECT 1380.560 66.650 1380.820 66.970 ;
        RECT 1380.620 17.410 1380.760 66.650 ;
        RECT 1380.160 17.270 1380.760 17.410 ;
        RECT 1380.160 2.400 1380.300 17.270 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 66.540 621.390 66.600 ;
        RECT 1395.250 66.540 1395.570 66.600 ;
        RECT 621.070 66.400 1395.570 66.540 ;
        RECT 621.070 66.340 621.390 66.400 ;
        RECT 1395.250 66.340 1395.570 66.400 ;
      LAYER via ;
        RECT 621.100 66.340 621.360 66.600 ;
        RECT 1395.280 66.340 1395.540 66.600 ;
      LAYER met2 ;
        RECT 621.910 400.250 622.190 404.000 ;
        RECT 621.160 400.110 622.190 400.250 ;
        RECT 621.160 66.630 621.300 400.110 ;
        RECT 621.910 400.000 622.190 400.110 ;
        RECT 621.100 66.310 621.360 66.630 ;
        RECT 1395.280 66.310 1395.540 66.630 ;
        RECT 1395.340 1.770 1395.480 66.310 ;
        RECT 1397.430 1.770 1397.990 2.400 ;
        RECT 1395.340 1.630 1397.990 1.770 ;
        RECT 1397.430 -4.800 1397.990 1.630 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.530 376.280 621.850 376.340 ;
        RECT 626.130 376.280 626.450 376.340 ;
        RECT 621.530 376.140 626.450 376.280 ;
        RECT 621.530 376.080 621.850 376.140 ;
        RECT 626.130 376.080 626.450 376.140 ;
        RECT 621.530 66.200 621.850 66.260 ;
        RECT 1415.490 66.200 1415.810 66.260 ;
        RECT 621.530 66.060 1415.810 66.200 ;
        RECT 621.530 66.000 621.850 66.060 ;
        RECT 1415.490 66.000 1415.810 66.060 ;
      LAYER via ;
        RECT 621.560 376.080 621.820 376.340 ;
        RECT 626.160 376.080 626.420 376.340 ;
        RECT 621.560 66.000 621.820 66.260 ;
        RECT 1415.520 66.000 1415.780 66.260 ;
      LAYER met2 ;
        RECT 627.430 400.250 627.710 404.000 ;
        RECT 626.220 400.110 627.710 400.250 ;
        RECT 626.220 376.370 626.360 400.110 ;
        RECT 627.430 400.000 627.710 400.110 ;
        RECT 621.560 376.050 621.820 376.370 ;
        RECT 626.160 376.050 626.420 376.370 ;
        RECT 621.620 66.290 621.760 376.050 ;
        RECT 621.560 65.970 621.820 66.290 ;
        RECT 1415.520 65.970 1415.780 66.290 ;
        RECT 1415.580 2.400 1415.720 65.970 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.430 375.940 628.750 376.000 ;
        RECT 631.190 375.940 631.510 376.000 ;
        RECT 628.430 375.800 631.510 375.940 ;
        RECT 628.430 375.740 628.750 375.800 ;
        RECT 631.190 375.740 631.510 375.800 ;
        RECT 628.430 65.860 628.750 65.920 ;
        RECT 1432.970 65.860 1433.290 65.920 ;
        RECT 628.430 65.720 1433.290 65.860 ;
        RECT 628.430 65.660 628.750 65.720 ;
        RECT 1432.970 65.660 1433.290 65.720 ;
      LAYER via ;
        RECT 628.460 375.740 628.720 376.000 ;
        RECT 631.220 375.740 631.480 376.000 ;
        RECT 628.460 65.660 628.720 65.920 ;
        RECT 1433.000 65.660 1433.260 65.920 ;
      LAYER met2 ;
        RECT 632.490 400.250 632.770 404.000 ;
        RECT 631.280 400.110 632.770 400.250 ;
        RECT 631.280 376.030 631.420 400.110 ;
        RECT 632.490 400.000 632.770 400.110 ;
        RECT 628.460 375.710 628.720 376.030 ;
        RECT 631.220 375.710 631.480 376.030 ;
        RECT 628.520 65.950 628.660 375.710 ;
        RECT 628.460 65.630 628.720 65.950 ;
        RECT 1433.000 65.630 1433.260 65.950 ;
        RECT 1433.060 2.400 1433.200 65.630 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.330 65.520 635.650 65.580 ;
        RECT 1449.070 65.520 1449.390 65.580 ;
        RECT 635.330 65.380 1449.390 65.520 ;
        RECT 635.330 65.320 635.650 65.380 ;
        RECT 1449.070 65.320 1449.390 65.380 ;
      LAYER via ;
        RECT 635.360 65.320 635.620 65.580 ;
        RECT 1449.100 65.320 1449.360 65.580 ;
      LAYER met2 ;
        RECT 638.010 400.250 638.290 404.000 ;
        RECT 636.800 400.110 638.290 400.250 ;
        RECT 636.800 399.570 636.940 400.110 ;
        RECT 638.010 400.000 638.290 400.110 ;
        RECT 635.420 399.430 636.940 399.570 ;
        RECT 635.420 65.610 635.560 399.430 ;
        RECT 635.360 65.290 635.620 65.610 ;
        RECT 1449.100 65.290 1449.360 65.610 ;
        RECT 1449.160 1.770 1449.300 65.290 ;
        RECT 1450.790 1.770 1451.350 2.400 ;
        RECT 1449.160 1.630 1451.350 1.770 ;
        RECT 1450.790 -4.800 1451.350 1.630 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.070 400.250 643.350 404.000 ;
        RECT 642.780 400.110 643.350 400.250 ;
        RECT 642.780 65.125 642.920 400.110 ;
        RECT 643.070 400.000 643.350 400.110 ;
        RECT 642.710 64.755 642.990 65.125 ;
        RECT 1466.110 64.755 1466.390 65.125 ;
        RECT 1466.180 1.770 1466.320 64.755 ;
        RECT 1468.270 1.770 1468.830 2.400 ;
        RECT 1466.180 1.630 1468.830 1.770 ;
        RECT 1468.270 -4.800 1468.830 1.630 ;
      LAYER via2 ;
        RECT 642.710 64.800 642.990 65.080 ;
        RECT 1466.110 64.800 1466.390 65.080 ;
      LAYER met3 ;
        RECT 642.685 65.090 643.015 65.105 ;
        RECT 1466.085 65.090 1466.415 65.105 ;
        RECT 642.685 64.790 1466.415 65.090 ;
        RECT 642.685 64.775 643.015 64.790 ;
        RECT 1466.085 64.775 1466.415 64.790 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 376.280 648.990 376.340 ;
        RECT 649.590 376.280 649.910 376.340 ;
        RECT 648.670 376.140 649.910 376.280 ;
        RECT 648.670 376.080 648.990 376.140 ;
        RECT 649.590 376.080 649.910 376.140 ;
        RECT 649.590 116.860 649.910 116.920 ;
        RECT 1483.570 116.860 1483.890 116.920 ;
        RECT 649.590 116.720 1483.890 116.860 ;
        RECT 649.590 116.660 649.910 116.720 ;
        RECT 1483.570 116.660 1483.890 116.720 ;
      LAYER via ;
        RECT 648.700 376.080 648.960 376.340 ;
        RECT 649.620 376.080 649.880 376.340 ;
        RECT 649.620 116.660 649.880 116.920 ;
        RECT 1483.600 116.660 1483.860 116.920 ;
      LAYER met2 ;
        RECT 648.590 400.180 648.870 404.000 ;
        RECT 648.590 400.000 648.900 400.180 ;
        RECT 648.760 376.370 648.900 400.000 ;
        RECT 648.700 376.050 648.960 376.370 ;
        RECT 649.620 376.050 649.880 376.370 ;
        RECT 649.680 116.950 649.820 376.050 ;
        RECT 649.620 116.630 649.880 116.950 ;
        RECT 1483.600 116.630 1483.860 116.950 ;
        RECT 1483.660 82.870 1483.800 116.630 ;
        RECT 1483.660 82.730 1486.560 82.870 ;
        RECT 1486.420 2.400 1486.560 82.730 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.050 119.240 650.370 119.300 ;
        RECT 1497.370 119.240 1497.690 119.300 ;
        RECT 650.050 119.100 1497.690 119.240 ;
        RECT 650.050 119.040 650.370 119.100 ;
        RECT 1497.370 119.040 1497.690 119.100 ;
        RECT 1497.370 15.200 1497.690 15.260 ;
        RECT 1503.810 15.200 1504.130 15.260 ;
        RECT 1497.370 15.060 1504.130 15.200 ;
        RECT 1497.370 15.000 1497.690 15.060 ;
        RECT 1503.810 15.000 1504.130 15.060 ;
      LAYER via ;
        RECT 650.080 119.040 650.340 119.300 ;
        RECT 1497.400 119.040 1497.660 119.300 ;
        RECT 1497.400 15.000 1497.660 15.260 ;
        RECT 1503.840 15.000 1504.100 15.260 ;
      LAYER met2 ;
        RECT 654.110 400.250 654.390 404.000 ;
        RECT 652.900 400.110 654.390 400.250 ;
        RECT 652.900 324.370 653.040 400.110 ;
        RECT 654.110 400.000 654.390 400.110 ;
        RECT 650.140 324.230 653.040 324.370 ;
        RECT 650.140 119.330 650.280 324.230 ;
        RECT 650.080 119.010 650.340 119.330 ;
        RECT 1497.400 119.010 1497.660 119.330 ;
        RECT 1497.460 15.290 1497.600 119.010 ;
        RECT 1497.400 14.970 1497.660 15.290 ;
        RECT 1503.840 14.970 1504.100 15.290 ;
        RECT 1503.900 2.400 1504.040 14.970 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.090 386.140 408.410 386.200 ;
        RECT 411.770 386.140 412.090 386.200 ;
        RECT 408.090 386.000 412.090 386.140 ;
        RECT 408.090 385.940 408.410 386.000 ;
        RECT 411.770 385.940 412.090 386.000 ;
        RECT 408.090 31.860 408.410 31.920 ;
        RECT 706.170 31.860 706.490 31.920 ;
        RECT 408.090 31.720 706.490 31.860 ;
        RECT 408.090 31.660 408.410 31.720 ;
        RECT 706.170 31.660 706.490 31.720 ;
      LAYER via ;
        RECT 408.120 385.940 408.380 386.200 ;
        RECT 411.800 385.940 412.060 386.200 ;
        RECT 408.120 31.660 408.380 31.920 ;
        RECT 706.200 31.660 706.460 31.920 ;
      LAYER met2 ;
        RECT 413.070 400.250 413.350 404.000 ;
        RECT 411.860 400.110 413.350 400.250 ;
        RECT 411.860 386.230 412.000 400.110 ;
        RECT 413.070 400.000 413.350 400.110 ;
        RECT 408.120 385.910 408.380 386.230 ;
        RECT 411.800 385.910 412.060 386.230 ;
        RECT 408.180 31.950 408.320 385.910 ;
        RECT 408.120 31.630 408.380 31.950 ;
        RECT 706.200 31.630 706.460 31.950 ;
        RECT 706.260 2.400 706.400 31.630 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.950 119.580 657.270 119.640 ;
        RECT 1518.070 119.580 1518.390 119.640 ;
        RECT 656.950 119.440 1518.390 119.580 ;
        RECT 656.950 119.380 657.270 119.440 ;
        RECT 1518.070 119.380 1518.390 119.440 ;
      LAYER via ;
        RECT 656.980 119.380 657.240 119.640 ;
        RECT 1518.100 119.380 1518.360 119.640 ;
      LAYER met2 ;
        RECT 659.170 400.250 659.450 404.000 ;
        RECT 658.420 400.110 659.450 400.250 ;
        RECT 658.420 324.370 658.560 400.110 ;
        RECT 659.170 400.000 659.450 400.110 ;
        RECT 657.040 324.230 658.560 324.370 ;
        RECT 657.040 119.670 657.180 324.230 ;
        RECT 656.980 119.350 657.240 119.670 ;
        RECT 1518.100 119.350 1518.360 119.670 ;
        RECT 1518.160 82.870 1518.300 119.350 ;
        RECT 1518.160 82.730 1519.680 82.870 ;
        RECT 1519.540 1.770 1519.680 82.730 ;
        RECT 1521.630 1.770 1522.190 2.400 ;
        RECT 1519.540 1.630 1522.190 1.770 ;
        RECT 1521.630 -4.800 1522.190 1.630 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.850 119.920 664.170 119.980 ;
        RECT 1538.770 119.920 1539.090 119.980 ;
        RECT 663.850 119.780 1539.090 119.920 ;
        RECT 663.850 119.720 664.170 119.780 ;
        RECT 1538.770 119.720 1539.090 119.780 ;
      LAYER via ;
        RECT 663.880 119.720 664.140 119.980 ;
        RECT 1538.800 119.720 1539.060 119.980 ;
      LAYER met2 ;
        RECT 664.690 400.250 664.970 404.000 ;
        RECT 664.400 400.110 664.970 400.250 ;
        RECT 664.400 351.970 664.540 400.110 ;
        RECT 664.690 400.000 664.970 400.110 ;
        RECT 663.940 351.830 664.540 351.970 ;
        RECT 663.940 120.010 664.080 351.830 ;
        RECT 663.880 119.690 664.140 120.010 ;
        RECT 1538.800 119.690 1539.060 120.010 ;
        RECT 1538.860 17.410 1539.000 119.690 ;
        RECT 1538.860 17.270 1539.920 17.410 ;
        RECT 1539.780 2.400 1539.920 17.270 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.750 120.260 671.070 120.320 ;
        RECT 1552.570 120.260 1552.890 120.320 ;
        RECT 670.750 120.120 1552.890 120.260 ;
        RECT 670.750 120.060 671.070 120.120 ;
        RECT 1552.570 120.060 1552.890 120.120 ;
      LAYER via ;
        RECT 670.780 120.060 671.040 120.320 ;
        RECT 1552.600 120.060 1552.860 120.320 ;
      LAYER met2 ;
        RECT 670.210 400.250 670.490 404.000 ;
        RECT 670.210 400.110 670.980 400.250 ;
        RECT 670.210 400.000 670.490 400.110 ;
        RECT 670.840 120.350 670.980 400.110 ;
        RECT 670.780 120.030 671.040 120.350 ;
        RECT 1552.600 120.030 1552.860 120.350 ;
        RECT 1552.660 82.870 1552.800 120.030 ;
        RECT 1552.660 82.730 1557.400 82.870 ;
        RECT 1557.260 2.400 1557.400 82.730 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.830 376.620 670.150 376.680 ;
        RECT 673.970 376.620 674.290 376.680 ;
        RECT 669.830 376.480 674.290 376.620 ;
        RECT 669.830 376.420 670.150 376.480 ;
        RECT 673.970 376.420 674.290 376.480 ;
        RECT 669.830 70.620 670.150 70.680 ;
        RECT 1573.270 70.620 1573.590 70.680 ;
        RECT 669.830 70.480 1573.590 70.620 ;
        RECT 669.830 70.420 670.150 70.480 ;
        RECT 1573.270 70.420 1573.590 70.480 ;
      LAYER via ;
        RECT 669.860 376.420 670.120 376.680 ;
        RECT 674.000 376.420 674.260 376.680 ;
        RECT 669.860 70.420 670.120 70.680 ;
        RECT 1573.300 70.420 1573.560 70.680 ;
      LAYER met2 ;
        RECT 675.270 400.250 675.550 404.000 ;
        RECT 674.060 400.110 675.550 400.250 ;
        RECT 674.060 376.710 674.200 400.110 ;
        RECT 675.270 400.000 675.550 400.110 ;
        RECT 669.860 376.390 670.120 376.710 ;
        RECT 674.000 376.390 674.260 376.710 ;
        RECT 669.920 70.710 670.060 376.390 ;
        RECT 669.860 70.390 670.120 70.710 ;
        RECT 1573.300 70.390 1573.560 70.710 ;
        RECT 1573.360 1.770 1573.500 70.390 ;
        RECT 1574.990 1.770 1575.550 2.400 ;
        RECT 1573.360 1.630 1575.550 1.770 ;
        RECT 1574.990 -4.800 1575.550 1.630 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.730 375.940 677.050 376.000 ;
        RECT 679.490 375.940 679.810 376.000 ;
        RECT 676.730 375.800 679.810 375.940 ;
        RECT 676.730 375.740 677.050 375.800 ;
        RECT 679.490 375.740 679.810 375.800 ;
        RECT 676.730 70.960 677.050 71.020 ;
        RECT 1590.290 70.960 1590.610 71.020 ;
        RECT 676.730 70.820 1590.610 70.960 ;
        RECT 676.730 70.760 677.050 70.820 ;
        RECT 1590.290 70.760 1590.610 70.820 ;
      LAYER via ;
        RECT 676.760 375.740 677.020 376.000 ;
        RECT 679.520 375.740 679.780 376.000 ;
        RECT 676.760 70.760 677.020 71.020 ;
        RECT 1590.320 70.760 1590.580 71.020 ;
      LAYER met2 ;
        RECT 680.790 400.250 681.070 404.000 ;
        RECT 679.580 400.110 681.070 400.250 ;
        RECT 679.580 376.030 679.720 400.110 ;
        RECT 680.790 400.000 681.070 400.110 ;
        RECT 676.760 375.710 677.020 376.030 ;
        RECT 679.520 375.710 679.780 376.030 ;
        RECT 676.820 71.050 676.960 375.710 ;
        RECT 676.760 70.730 677.020 71.050 ;
        RECT 1590.320 70.730 1590.580 71.050 ;
        RECT 1590.380 1.770 1590.520 70.730 ;
        RECT 1592.470 1.770 1593.030 2.400 ;
        RECT 1590.380 1.630 1593.030 1.770 ;
        RECT 1592.470 -4.800 1593.030 1.630 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.090 71.300 684.410 71.360 ;
        RECT 1610.530 71.300 1610.850 71.360 ;
        RECT 684.090 71.160 1610.850 71.300 ;
        RECT 684.090 71.100 684.410 71.160 ;
        RECT 1610.530 71.100 1610.850 71.160 ;
      LAYER via ;
        RECT 684.120 71.100 684.380 71.360 ;
        RECT 1610.560 71.100 1610.820 71.360 ;
      LAYER met2 ;
        RECT 686.310 400.250 686.590 404.000 ;
        RECT 685.100 400.110 686.590 400.250 ;
        RECT 685.100 351.970 685.240 400.110 ;
        RECT 686.310 400.000 686.590 400.110 ;
        RECT 684.180 351.830 685.240 351.970 ;
        RECT 684.180 71.390 684.320 351.830 ;
        RECT 684.120 71.070 684.380 71.390 ;
        RECT 1610.560 71.070 1610.820 71.390 ;
        RECT 1610.620 2.400 1610.760 71.070 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.530 71.640 690.850 71.700 ;
        RECT 1621.570 71.640 1621.890 71.700 ;
        RECT 690.530 71.500 1621.890 71.640 ;
        RECT 690.530 71.440 690.850 71.500 ;
        RECT 1621.570 71.440 1621.890 71.500 ;
        RECT 1621.570 15.200 1621.890 15.260 ;
        RECT 1628.010 15.200 1628.330 15.260 ;
        RECT 1621.570 15.060 1628.330 15.200 ;
        RECT 1621.570 15.000 1621.890 15.060 ;
        RECT 1628.010 15.000 1628.330 15.060 ;
      LAYER via ;
        RECT 690.560 71.440 690.820 71.700 ;
        RECT 1621.600 71.440 1621.860 71.700 ;
        RECT 1621.600 15.000 1621.860 15.260 ;
        RECT 1628.040 15.000 1628.300 15.260 ;
      LAYER met2 ;
        RECT 691.370 400.250 691.650 404.000 ;
        RECT 690.620 400.110 691.650 400.250 ;
        RECT 690.620 71.730 690.760 400.110 ;
        RECT 691.370 400.000 691.650 400.110 ;
        RECT 690.560 71.410 690.820 71.730 ;
        RECT 1621.600 71.410 1621.860 71.730 ;
        RECT 1621.660 15.290 1621.800 71.410 ;
        RECT 1621.600 14.970 1621.860 15.290 ;
        RECT 1628.040 14.970 1628.300 15.290 ;
        RECT 1628.100 2.400 1628.240 14.970 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.890 71.980 698.210 72.040 ;
        RECT 1643.650 71.980 1643.970 72.040 ;
        RECT 697.890 71.840 1643.970 71.980 ;
        RECT 697.890 71.780 698.210 71.840 ;
        RECT 1643.650 71.780 1643.970 71.840 ;
      LAYER via ;
        RECT 697.920 71.780 698.180 72.040 ;
        RECT 1643.680 71.780 1643.940 72.040 ;
      LAYER met2 ;
        RECT 696.890 400.250 697.170 404.000 ;
        RECT 696.890 400.110 698.120 400.250 ;
        RECT 696.890 400.000 697.170 400.110 ;
        RECT 697.980 72.070 698.120 400.110 ;
        RECT 697.920 71.750 698.180 72.070 ;
        RECT 1643.680 71.750 1643.940 72.070 ;
        RECT 1643.740 1.770 1643.880 71.750 ;
        RECT 1645.830 1.770 1646.390 2.400 ;
        RECT 1643.740 1.630 1646.390 1.770 ;
        RECT 1645.830 -4.800 1646.390 1.630 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.430 386.480 697.750 386.540 ;
        RECT 701.110 386.480 701.430 386.540 ;
        RECT 697.430 386.340 701.430 386.480 ;
        RECT 697.430 386.280 697.750 386.340 ;
        RECT 701.110 386.280 701.430 386.340 ;
        RECT 697.430 75.720 697.750 75.780 ;
        RECT 1663.430 75.720 1663.750 75.780 ;
        RECT 697.430 75.580 1663.750 75.720 ;
        RECT 697.430 75.520 697.750 75.580 ;
        RECT 1663.430 75.520 1663.750 75.580 ;
      LAYER via ;
        RECT 697.460 386.280 697.720 386.540 ;
        RECT 701.140 386.280 701.400 386.540 ;
        RECT 697.460 75.520 697.720 75.780 ;
        RECT 1663.460 75.520 1663.720 75.780 ;
      LAYER met2 ;
        RECT 702.410 400.250 702.690 404.000 ;
        RECT 701.200 400.110 702.690 400.250 ;
        RECT 701.200 386.570 701.340 400.110 ;
        RECT 702.410 400.000 702.690 400.110 ;
        RECT 697.460 386.250 697.720 386.570 ;
        RECT 701.140 386.250 701.400 386.570 ;
        RECT 697.520 75.810 697.660 386.250 ;
        RECT 697.460 75.490 697.720 75.810 ;
        RECT 1663.460 75.490 1663.720 75.810 ;
        RECT 1663.520 2.400 1663.660 75.490 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.330 75.380 704.650 75.440 ;
        RECT 1681.370 75.380 1681.690 75.440 ;
        RECT 704.330 75.240 1681.690 75.380 ;
        RECT 704.330 75.180 704.650 75.240 ;
        RECT 1681.370 75.180 1681.690 75.240 ;
      LAYER via ;
        RECT 704.360 75.180 704.620 75.440 ;
        RECT 1681.400 75.180 1681.660 75.440 ;
      LAYER met2 ;
        RECT 707.470 400.250 707.750 404.000 ;
        RECT 706.260 400.110 707.750 400.250 ;
        RECT 706.260 385.970 706.400 400.110 ;
        RECT 707.470 400.000 707.750 400.110 ;
        RECT 704.420 385.830 706.400 385.970 ;
        RECT 704.420 75.470 704.560 385.830 ;
        RECT 704.360 75.150 704.620 75.470 ;
        RECT 1681.400 75.150 1681.660 75.470 ;
        RECT 1681.460 2.400 1681.600 75.150 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 415.450 46.140 415.770 46.200 ;
        RECT 723.650 46.140 723.970 46.200 ;
        RECT 415.450 46.000 723.970 46.140 ;
        RECT 415.450 45.940 415.770 46.000 ;
        RECT 723.650 45.940 723.970 46.000 ;
      LAYER via ;
        RECT 415.480 45.940 415.740 46.200 ;
        RECT 723.680 45.940 723.940 46.200 ;
      LAYER met2 ;
        RECT 418.130 400.250 418.410 404.000 ;
        RECT 416.920 400.110 418.410 400.250 ;
        RECT 416.920 324.370 417.060 400.110 ;
        RECT 418.130 400.000 418.410 400.110 ;
        RECT 415.540 324.230 417.060 324.370 ;
        RECT 415.540 46.230 415.680 324.230 ;
        RECT 415.480 45.910 415.740 46.230 ;
        RECT 723.680 45.910 723.940 46.230 ;
        RECT 723.740 2.400 723.880 45.910 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.690 75.040 712.010 75.100 ;
        RECT 1697.470 75.040 1697.790 75.100 ;
        RECT 711.690 74.900 1697.790 75.040 ;
        RECT 711.690 74.840 712.010 74.900 ;
        RECT 1697.470 74.840 1697.790 74.900 ;
      LAYER via ;
        RECT 711.720 74.840 711.980 75.100 ;
        RECT 1697.500 74.840 1697.760 75.100 ;
      LAYER met2 ;
        RECT 712.990 400.250 713.270 404.000 ;
        RECT 711.780 400.110 713.270 400.250 ;
        RECT 711.780 75.130 711.920 400.110 ;
        RECT 712.990 400.000 713.270 400.110 ;
        RECT 711.720 74.810 711.980 75.130 ;
        RECT 1697.500 74.810 1697.760 75.130 ;
        RECT 1697.560 1.770 1697.700 74.810 ;
        RECT 1699.190 1.770 1699.750 2.400 ;
        RECT 1697.560 1.630 1699.750 1.770 ;
        RECT 1699.190 -4.800 1699.750 1.630 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.130 74.700 718.450 74.760 ;
        RECT 1714.490 74.700 1714.810 74.760 ;
        RECT 718.130 74.560 1714.810 74.700 ;
        RECT 718.130 74.500 718.450 74.560 ;
        RECT 1714.490 74.500 1714.810 74.560 ;
      LAYER via ;
        RECT 718.160 74.500 718.420 74.760 ;
        RECT 1714.520 74.500 1714.780 74.760 ;
      LAYER met2 ;
        RECT 718.510 400.250 718.790 404.000 ;
        RECT 718.220 400.110 718.790 400.250 ;
        RECT 718.220 74.790 718.360 400.110 ;
        RECT 718.510 400.000 718.790 400.110 ;
        RECT 718.160 74.470 718.420 74.790 ;
        RECT 1714.520 74.470 1714.780 74.790 ;
        RECT 1714.580 1.770 1714.720 74.470 ;
        RECT 1716.670 1.770 1717.230 2.400 ;
        RECT 1714.580 1.630 1717.230 1.770 ;
        RECT 1716.670 -4.800 1717.230 1.630 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 717.670 386.140 717.990 386.200 ;
        RECT 722.270 386.140 722.590 386.200 ;
        RECT 717.670 386.000 722.590 386.140 ;
        RECT 717.670 385.940 717.990 386.000 ;
        RECT 722.270 385.940 722.590 386.000 ;
        RECT 717.670 74.360 717.990 74.420 ;
        RECT 1734.730 74.360 1735.050 74.420 ;
        RECT 717.670 74.220 1735.050 74.360 ;
        RECT 717.670 74.160 717.990 74.220 ;
        RECT 1734.730 74.160 1735.050 74.220 ;
      LAYER via ;
        RECT 717.700 385.940 717.960 386.200 ;
        RECT 722.300 385.940 722.560 386.200 ;
        RECT 717.700 74.160 717.960 74.420 ;
        RECT 1734.760 74.160 1735.020 74.420 ;
      LAYER met2 ;
        RECT 723.570 400.250 723.850 404.000 ;
        RECT 722.360 400.110 723.850 400.250 ;
        RECT 722.360 386.230 722.500 400.110 ;
        RECT 723.570 400.000 723.850 400.110 ;
        RECT 717.700 385.910 717.960 386.230 ;
        RECT 722.300 385.910 722.560 386.230 ;
        RECT 717.760 74.450 717.900 385.910 ;
        RECT 717.700 74.130 717.960 74.450 ;
        RECT 1734.760 74.130 1735.020 74.450 ;
        RECT 1734.820 2.400 1734.960 74.130 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 724.570 386.820 724.890 386.880 ;
        RECT 727.790 386.820 728.110 386.880 ;
        RECT 724.570 386.680 728.110 386.820 ;
        RECT 724.570 386.620 724.890 386.680 ;
        RECT 727.790 386.620 728.110 386.680 ;
        RECT 724.570 74.020 724.890 74.080 ;
        RECT 1746.230 74.020 1746.550 74.080 ;
        RECT 724.570 73.880 1746.550 74.020 ;
        RECT 724.570 73.820 724.890 73.880 ;
        RECT 1746.230 73.820 1746.550 73.880 ;
        RECT 1746.230 15.200 1746.550 15.260 ;
        RECT 1752.210 15.200 1752.530 15.260 ;
        RECT 1746.230 15.060 1752.530 15.200 ;
        RECT 1746.230 15.000 1746.550 15.060 ;
        RECT 1752.210 15.000 1752.530 15.060 ;
      LAYER via ;
        RECT 724.600 386.620 724.860 386.880 ;
        RECT 727.820 386.620 728.080 386.880 ;
        RECT 724.600 73.820 724.860 74.080 ;
        RECT 1746.260 73.820 1746.520 74.080 ;
        RECT 1746.260 15.000 1746.520 15.260 ;
        RECT 1752.240 15.000 1752.500 15.260 ;
      LAYER met2 ;
        RECT 729.090 400.250 729.370 404.000 ;
        RECT 727.880 400.110 729.370 400.250 ;
        RECT 727.880 386.910 728.020 400.110 ;
        RECT 729.090 400.000 729.370 400.110 ;
        RECT 724.600 386.590 724.860 386.910 ;
        RECT 727.820 386.590 728.080 386.910 ;
        RECT 724.660 74.110 724.800 386.590 ;
        RECT 724.600 73.790 724.860 74.110 ;
        RECT 1746.260 73.790 1746.520 74.110 ;
        RECT 1746.320 15.290 1746.460 73.790 ;
        RECT 1746.260 14.970 1746.520 15.290 ;
        RECT 1752.240 14.970 1752.500 15.290 ;
        RECT 1752.300 2.400 1752.440 14.970 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.470 386.480 731.790 386.540 ;
        RECT 733.310 386.480 733.630 386.540 ;
        RECT 731.470 386.340 733.630 386.480 ;
        RECT 731.470 386.280 731.790 386.340 ;
        RECT 733.310 386.280 733.630 386.340 ;
        RECT 731.470 73.680 731.790 73.740 ;
        RECT 1767.850 73.680 1768.170 73.740 ;
        RECT 731.470 73.540 1768.170 73.680 ;
        RECT 731.470 73.480 731.790 73.540 ;
        RECT 1767.850 73.480 1768.170 73.540 ;
      LAYER via ;
        RECT 731.500 386.280 731.760 386.540 ;
        RECT 733.340 386.280 733.600 386.540 ;
        RECT 731.500 73.480 731.760 73.740 ;
        RECT 1767.880 73.480 1768.140 73.740 ;
      LAYER met2 ;
        RECT 734.150 400.250 734.430 404.000 ;
        RECT 733.400 400.110 734.430 400.250 ;
        RECT 733.400 386.570 733.540 400.110 ;
        RECT 734.150 400.000 734.430 400.110 ;
        RECT 731.500 386.250 731.760 386.570 ;
        RECT 733.340 386.250 733.600 386.570 ;
        RECT 731.560 73.770 731.700 386.250 ;
        RECT 731.500 73.450 731.760 73.770 ;
        RECT 1767.880 73.450 1768.140 73.770 ;
        RECT 1767.940 1.770 1768.080 73.450 ;
        RECT 1770.030 1.770 1770.590 2.400 ;
        RECT 1767.940 1.630 1770.590 1.770 ;
        RECT 1770.030 -4.800 1770.590 1.630 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.370 73.340 738.690 73.400 ;
        RECT 1787.630 73.340 1787.950 73.400 ;
        RECT 738.370 73.200 1787.950 73.340 ;
        RECT 738.370 73.140 738.690 73.200 ;
        RECT 1787.630 73.140 1787.950 73.200 ;
      LAYER via ;
        RECT 738.400 73.140 738.660 73.400 ;
        RECT 1787.660 73.140 1787.920 73.400 ;
      LAYER met2 ;
        RECT 739.670 400.250 739.950 404.000 ;
        RECT 738.460 400.110 739.950 400.250 ;
        RECT 738.460 73.430 738.600 400.110 ;
        RECT 739.670 400.000 739.950 400.110 ;
        RECT 738.400 73.110 738.660 73.430 ;
        RECT 1787.660 73.110 1787.920 73.430 ;
        RECT 1787.720 2.400 1787.860 73.110 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 746.190 73.000 746.510 73.060 ;
        RECT 1805.570 73.000 1805.890 73.060 ;
        RECT 746.190 72.860 1805.890 73.000 ;
        RECT 746.190 72.800 746.510 72.860 ;
        RECT 1805.570 72.800 1805.890 72.860 ;
      LAYER via ;
        RECT 746.220 72.800 746.480 73.060 ;
        RECT 1805.600 72.800 1805.860 73.060 ;
      LAYER met2 ;
        RECT 745.190 400.250 745.470 404.000 ;
        RECT 745.190 400.110 746.420 400.250 ;
        RECT 745.190 400.000 745.470 400.110 ;
        RECT 746.280 73.090 746.420 400.110 ;
        RECT 746.220 72.770 746.480 73.090 ;
        RECT 1805.600 72.770 1805.860 73.090 ;
        RECT 1805.660 2.400 1805.800 72.770 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.730 386.480 746.050 386.540 ;
        RECT 749.410 386.480 749.730 386.540 ;
        RECT 745.730 386.340 749.730 386.480 ;
        RECT 745.730 386.280 746.050 386.340 ;
        RECT 749.410 386.280 749.730 386.340 ;
        RECT 745.730 72.660 746.050 72.720 ;
        RECT 1823.050 72.660 1823.370 72.720 ;
        RECT 745.730 72.520 1823.370 72.660 ;
        RECT 745.730 72.460 746.050 72.520 ;
        RECT 1823.050 72.460 1823.370 72.520 ;
      LAYER via ;
        RECT 745.760 386.280 746.020 386.540 ;
        RECT 749.440 386.280 749.700 386.540 ;
        RECT 745.760 72.460 746.020 72.720 ;
        RECT 1823.080 72.460 1823.340 72.720 ;
      LAYER met2 ;
        RECT 750.250 400.250 750.530 404.000 ;
        RECT 749.500 400.110 750.530 400.250 ;
        RECT 749.500 386.570 749.640 400.110 ;
        RECT 750.250 400.000 750.530 400.110 ;
        RECT 745.760 386.250 746.020 386.570 ;
        RECT 749.440 386.250 749.700 386.570 ;
        RECT 745.820 72.750 745.960 386.250 ;
        RECT 745.760 72.430 746.020 72.750 ;
        RECT 1823.080 72.430 1823.340 72.750 ;
        RECT 1823.140 2.400 1823.280 72.430 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.630 72.320 752.950 72.380 ;
        RECT 1838.690 72.320 1839.010 72.380 ;
        RECT 752.630 72.180 1839.010 72.320 ;
        RECT 752.630 72.120 752.950 72.180 ;
        RECT 1838.690 72.120 1839.010 72.180 ;
      LAYER via ;
        RECT 752.660 72.120 752.920 72.380 ;
        RECT 1838.720 72.120 1838.980 72.380 ;
      LAYER met2 ;
        RECT 755.770 400.250 756.050 404.000 ;
        RECT 754.560 400.110 756.050 400.250 ;
        RECT 754.560 385.970 754.700 400.110 ;
        RECT 755.770 400.000 756.050 400.110 ;
        RECT 752.720 385.830 754.700 385.970 ;
        RECT 752.720 72.410 752.860 385.830 ;
        RECT 752.660 72.090 752.920 72.410 ;
        RECT 1838.720 72.090 1838.980 72.410 ;
        RECT 1838.780 1.770 1838.920 72.090 ;
        RECT 1840.870 1.770 1841.430 2.400 ;
        RECT 1838.780 1.630 1841.430 1.770 ;
        RECT 1840.870 -4.800 1841.430 1.630 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.290 400.250 761.570 404.000 ;
        RECT 760.080 400.110 761.570 400.250 ;
        RECT 760.080 72.605 760.220 400.110 ;
        RECT 761.290 400.000 761.570 400.110 ;
        RECT 760.010 72.235 760.290 72.605 ;
        RECT 1856.190 72.235 1856.470 72.605 ;
        RECT 1856.260 1.770 1856.400 72.235 ;
        RECT 1858.350 1.770 1858.910 2.400 ;
        RECT 1856.260 1.630 1858.910 1.770 ;
        RECT 1858.350 -4.800 1858.910 1.630 ;
      LAYER via2 ;
        RECT 760.010 72.280 760.290 72.560 ;
        RECT 1856.190 72.280 1856.470 72.560 ;
      LAYER met3 ;
        RECT 759.985 72.570 760.315 72.585 ;
        RECT 1856.165 72.570 1856.495 72.585 ;
        RECT 759.985 72.270 1856.495 72.570 ;
        RECT 759.985 72.255 760.315 72.270 ;
        RECT 1856.165 72.255 1856.495 72.270 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 422.350 45.800 422.670 45.860 ;
        RECT 741.590 45.800 741.910 45.860 ;
        RECT 422.350 45.660 741.910 45.800 ;
        RECT 422.350 45.600 422.670 45.660 ;
        RECT 741.590 45.600 741.910 45.660 ;
      LAYER via ;
        RECT 422.380 45.600 422.640 45.860 ;
        RECT 741.620 45.600 741.880 45.860 ;
      LAYER met2 ;
        RECT 423.650 400.250 423.930 404.000 ;
        RECT 422.440 400.110 423.930 400.250 ;
        RECT 422.440 45.890 422.580 400.110 ;
        RECT 423.650 400.000 423.930 400.110 ;
        RECT 422.380 45.570 422.640 45.890 ;
        RECT 741.620 45.570 741.880 45.890 ;
        RECT 741.680 2.400 741.820 45.570 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.890 124.000 767.210 124.060 ;
        RECT 1869.970 124.000 1870.290 124.060 ;
        RECT 766.890 123.860 1870.290 124.000 ;
        RECT 766.890 123.800 767.210 123.860 ;
        RECT 1869.970 123.800 1870.290 123.860 ;
        RECT 1869.970 15.200 1870.290 15.260 ;
        RECT 1876.410 15.200 1876.730 15.260 ;
        RECT 1869.970 15.060 1876.730 15.200 ;
        RECT 1869.970 15.000 1870.290 15.060 ;
        RECT 1876.410 15.000 1876.730 15.060 ;
      LAYER via ;
        RECT 766.920 123.800 767.180 124.060 ;
        RECT 1870.000 123.800 1870.260 124.060 ;
        RECT 1870.000 15.000 1870.260 15.260 ;
        RECT 1876.440 15.000 1876.700 15.260 ;
      LAYER met2 ;
        RECT 766.350 400.250 766.630 404.000 ;
        RECT 766.350 400.110 767.120 400.250 ;
        RECT 766.350 400.000 766.630 400.110 ;
        RECT 766.980 124.090 767.120 400.110 ;
        RECT 766.920 123.770 767.180 124.090 ;
        RECT 1870.000 123.770 1870.260 124.090 ;
        RECT 1870.060 15.290 1870.200 123.770 ;
        RECT 1870.000 14.970 1870.260 15.290 ;
        RECT 1876.440 14.970 1876.700 15.290 ;
        RECT 1876.500 2.400 1876.640 14.970 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.430 386.140 766.750 386.200 ;
        RECT 770.570 386.140 770.890 386.200 ;
        RECT 766.430 386.000 770.890 386.140 ;
        RECT 766.430 385.940 766.750 386.000 ;
        RECT 770.570 385.940 770.890 386.000 ;
        RECT 766.430 123.660 766.750 123.720 ;
        RECT 1890.670 123.660 1890.990 123.720 ;
        RECT 766.430 123.520 1890.990 123.660 ;
        RECT 766.430 123.460 766.750 123.520 ;
        RECT 1890.670 123.460 1890.990 123.520 ;
      LAYER via ;
        RECT 766.460 385.940 766.720 386.200 ;
        RECT 770.600 385.940 770.860 386.200 ;
        RECT 766.460 123.460 766.720 123.720 ;
        RECT 1890.700 123.460 1890.960 123.720 ;
      LAYER met2 ;
        RECT 771.870 400.250 772.150 404.000 ;
        RECT 770.660 400.110 772.150 400.250 ;
        RECT 770.660 386.230 770.800 400.110 ;
        RECT 771.870 400.000 772.150 400.110 ;
        RECT 766.460 385.910 766.720 386.230 ;
        RECT 770.600 385.910 770.860 386.230 ;
        RECT 766.520 123.750 766.660 385.910 ;
        RECT 766.460 123.430 766.720 123.750 ;
        RECT 1890.700 123.430 1890.960 123.750 ;
        RECT 1890.760 82.870 1890.900 123.430 ;
        RECT 1890.760 82.730 1892.280 82.870 ;
        RECT 1892.140 1.770 1892.280 82.730 ;
        RECT 1894.230 1.770 1894.790 2.400 ;
        RECT 1892.140 1.630 1894.790 1.770 ;
        RECT 1894.230 -4.800 1894.790 1.630 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.330 123.320 773.650 123.380 ;
        RECT 1911.830 123.320 1912.150 123.380 ;
        RECT 773.330 123.180 1912.150 123.320 ;
        RECT 773.330 123.120 773.650 123.180 ;
        RECT 1911.830 123.120 1912.150 123.180 ;
      LAYER via ;
        RECT 773.360 123.120 773.620 123.380 ;
        RECT 1911.860 123.120 1912.120 123.380 ;
      LAYER met2 ;
        RECT 777.390 400.250 777.670 404.000 ;
        RECT 776.180 400.110 777.670 400.250 ;
        RECT 776.180 385.970 776.320 400.110 ;
        RECT 777.390 400.000 777.670 400.110 ;
        RECT 773.420 385.830 776.320 385.970 ;
        RECT 773.420 123.410 773.560 385.830 ;
        RECT 773.360 123.090 773.620 123.410 ;
        RECT 1911.860 123.090 1912.120 123.410 ;
        RECT 1911.920 2.400 1912.060 123.090 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.690 122.980 781.010 123.040 ;
        RECT 1925.170 122.980 1925.490 123.040 ;
        RECT 780.690 122.840 1925.490 122.980 ;
        RECT 780.690 122.780 781.010 122.840 ;
        RECT 1925.170 122.780 1925.490 122.840 ;
      LAYER via ;
        RECT 780.720 122.780 780.980 123.040 ;
        RECT 1925.200 122.780 1925.460 123.040 ;
      LAYER met2 ;
        RECT 782.450 400.250 782.730 404.000 ;
        RECT 781.240 400.110 782.730 400.250 ;
        RECT 781.240 324.370 781.380 400.110 ;
        RECT 782.450 400.000 782.730 400.110 ;
        RECT 780.780 324.230 781.380 324.370 ;
        RECT 780.780 123.070 780.920 324.230 ;
        RECT 780.720 122.750 780.980 123.070 ;
        RECT 1925.200 122.750 1925.460 123.070 ;
        RECT 1925.260 82.870 1925.400 122.750 ;
        RECT 1925.260 82.730 1928.160 82.870 ;
        RECT 1928.020 17.410 1928.160 82.730 ;
        RECT 1928.020 17.270 1930.000 17.410 ;
        RECT 1929.860 2.400 1930.000 17.270 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.130 122.640 787.450 122.700 ;
        RECT 1945.870 122.640 1946.190 122.700 ;
        RECT 787.130 122.500 1946.190 122.640 ;
        RECT 787.130 122.440 787.450 122.500 ;
        RECT 1945.870 122.440 1946.190 122.500 ;
      LAYER via ;
        RECT 787.160 122.440 787.420 122.700 ;
        RECT 1945.900 122.440 1946.160 122.700 ;
      LAYER met2 ;
        RECT 787.970 400.250 788.250 404.000 ;
        RECT 787.220 400.110 788.250 400.250 ;
        RECT 787.220 122.730 787.360 400.110 ;
        RECT 787.970 400.000 788.250 400.110 ;
        RECT 787.160 122.410 787.420 122.730 ;
        RECT 1945.900 122.410 1946.160 122.730 ;
        RECT 1945.960 82.870 1946.100 122.410 ;
        RECT 1945.960 82.730 1947.480 82.870 ;
        RECT 1947.340 2.400 1947.480 82.730 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.030 78.100 794.350 78.160 ;
        RECT 1962.890 78.100 1963.210 78.160 ;
        RECT 794.030 77.960 1963.210 78.100 ;
        RECT 794.030 77.900 794.350 77.960 ;
        RECT 1962.890 77.900 1963.210 77.960 ;
      LAYER via ;
        RECT 794.060 77.900 794.320 78.160 ;
        RECT 1962.920 77.900 1963.180 78.160 ;
      LAYER met2 ;
        RECT 793.490 400.250 793.770 404.000 ;
        RECT 793.490 400.110 794.260 400.250 ;
        RECT 793.490 400.000 793.770 400.110 ;
        RECT 794.120 78.190 794.260 400.110 ;
        RECT 794.060 77.870 794.320 78.190 ;
        RECT 1962.920 77.870 1963.180 78.190 ;
        RECT 1962.980 1.770 1963.120 77.870 ;
        RECT 1965.070 1.770 1965.630 2.400 ;
        RECT 1962.980 1.630 1965.630 1.770 ;
        RECT 1965.070 -4.800 1965.630 1.630 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.490 78.440 794.810 78.500 ;
        RECT 1980.370 78.440 1980.690 78.500 ;
        RECT 794.490 78.300 1980.690 78.440 ;
        RECT 794.490 78.240 794.810 78.300 ;
        RECT 1980.370 78.240 1980.690 78.300 ;
      LAYER via ;
        RECT 794.520 78.240 794.780 78.500 ;
        RECT 1980.400 78.240 1980.660 78.500 ;
      LAYER met2 ;
        RECT 798.550 400.250 798.830 404.000 ;
        RECT 797.340 400.110 798.830 400.250 ;
        RECT 797.340 324.370 797.480 400.110 ;
        RECT 798.550 400.000 798.830 400.110 ;
        RECT 794.580 324.230 797.480 324.370 ;
        RECT 794.580 78.530 794.720 324.230 ;
        RECT 794.520 78.210 794.780 78.530 ;
        RECT 1980.400 78.210 1980.660 78.530 ;
        RECT 1980.460 1.770 1980.600 78.210 ;
        RECT 1982.550 1.770 1983.110 2.400 ;
        RECT 1980.460 1.630 1983.110 1.770 ;
        RECT 1982.550 -4.800 1983.110 1.630 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.930 78.780 801.250 78.840 ;
        RECT 1994.170 78.780 1994.490 78.840 ;
        RECT 800.930 78.640 1994.490 78.780 ;
        RECT 800.930 78.580 801.250 78.640 ;
        RECT 1994.170 78.580 1994.490 78.640 ;
        RECT 1994.170 15.200 1994.490 15.260 ;
        RECT 2000.610 15.200 2000.930 15.260 ;
        RECT 1994.170 15.060 2000.930 15.200 ;
        RECT 1994.170 15.000 1994.490 15.060 ;
        RECT 2000.610 15.000 2000.930 15.060 ;
      LAYER via ;
        RECT 800.960 78.580 801.220 78.840 ;
        RECT 1994.200 78.580 1994.460 78.840 ;
        RECT 1994.200 15.000 1994.460 15.260 ;
        RECT 2000.640 15.000 2000.900 15.260 ;
      LAYER met2 ;
        RECT 804.070 400.250 804.350 404.000 ;
        RECT 802.860 400.110 804.350 400.250 ;
        RECT 802.860 385.290 803.000 400.110 ;
        RECT 804.070 400.000 804.350 400.110 ;
        RECT 801.020 385.150 803.000 385.290 ;
        RECT 801.020 78.870 801.160 385.150 ;
        RECT 800.960 78.550 801.220 78.870 ;
        RECT 1994.200 78.550 1994.460 78.870 ;
        RECT 1994.260 15.290 1994.400 78.550 ;
        RECT 1994.200 14.970 1994.460 15.290 ;
        RECT 2000.640 14.970 2000.900 15.290 ;
        RECT 2000.700 2.400 2000.840 14.970 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 808.290 79.120 808.610 79.180 ;
        RECT 2018.090 79.120 2018.410 79.180 ;
        RECT 808.290 78.980 2018.410 79.120 ;
        RECT 808.290 78.920 808.610 78.980 ;
        RECT 2018.090 78.920 2018.410 78.980 ;
      LAYER via ;
        RECT 808.320 78.920 808.580 79.180 ;
        RECT 2018.120 78.920 2018.380 79.180 ;
      LAYER met2 ;
        RECT 809.590 400.250 809.870 404.000 ;
        RECT 808.380 400.110 809.870 400.250 ;
        RECT 808.380 79.210 808.520 400.110 ;
        RECT 809.590 400.000 809.870 400.110 ;
        RECT 808.320 78.890 808.580 79.210 ;
        RECT 2018.120 78.890 2018.380 79.210 ;
        RECT 2018.180 2.400 2018.320 78.890 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 815.190 82.860 815.510 82.920 ;
        RECT 2036.030 82.860 2036.350 82.920 ;
        RECT 815.190 82.720 2036.350 82.860 ;
        RECT 815.190 82.660 815.510 82.720 ;
        RECT 2036.030 82.660 2036.350 82.720 ;
      LAYER via ;
        RECT 815.220 82.660 815.480 82.920 ;
        RECT 2036.060 82.660 2036.320 82.920 ;
      LAYER met2 ;
        RECT 814.650 400.250 814.930 404.000 ;
        RECT 814.650 400.110 815.420 400.250 ;
        RECT 814.650 400.000 814.930 400.110 ;
        RECT 815.280 82.950 815.420 400.110 ;
        RECT 815.220 82.630 815.480 82.950 ;
        RECT 2036.060 82.630 2036.320 82.950 ;
        RECT 2036.120 2.400 2036.260 82.630 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.790 45.460 429.110 45.520 ;
        RECT 759.070 45.460 759.390 45.520 ;
        RECT 428.790 45.320 759.390 45.460 ;
        RECT 428.790 45.260 429.110 45.320 ;
        RECT 759.070 45.260 759.390 45.320 ;
      LAYER via ;
        RECT 428.820 45.260 429.080 45.520 ;
        RECT 759.100 45.260 759.360 45.520 ;
      LAYER met2 ;
        RECT 429.170 400.250 429.450 404.000 ;
        RECT 428.880 400.110 429.450 400.250 ;
        RECT 428.880 45.550 429.020 400.110 ;
        RECT 429.170 400.000 429.450 400.110 ;
        RECT 428.820 45.230 429.080 45.550 ;
        RECT 759.100 45.230 759.360 45.550 ;
        RECT 759.160 2.400 759.300 45.230 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.730 386.140 815.050 386.200 ;
        RECT 818.870 386.140 819.190 386.200 ;
        RECT 814.730 386.000 819.190 386.140 ;
        RECT 814.730 385.940 815.050 386.000 ;
        RECT 818.870 385.940 819.190 386.000 ;
        RECT 814.730 82.520 815.050 82.580 ;
        RECT 2053.970 82.520 2054.290 82.580 ;
        RECT 814.730 82.380 2054.290 82.520 ;
        RECT 814.730 82.320 815.050 82.380 ;
        RECT 2053.970 82.320 2054.290 82.380 ;
      LAYER via ;
        RECT 814.760 385.940 815.020 386.200 ;
        RECT 818.900 385.940 819.160 386.200 ;
        RECT 814.760 82.320 815.020 82.580 ;
        RECT 2054.000 82.320 2054.260 82.580 ;
      LAYER met2 ;
        RECT 820.170 400.250 820.450 404.000 ;
        RECT 818.960 400.110 820.450 400.250 ;
        RECT 818.960 386.230 819.100 400.110 ;
        RECT 820.170 400.000 820.450 400.110 ;
        RECT 814.760 385.910 815.020 386.230 ;
        RECT 818.900 385.910 819.160 386.230 ;
        RECT 814.820 82.610 814.960 385.910 ;
        RECT 814.760 82.290 815.020 82.610 ;
        RECT 2054.000 82.290 2054.260 82.610 ;
        RECT 2054.060 2.400 2054.200 82.290 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.630 382.740 821.950 382.800 ;
        RECT 824.390 382.740 824.710 382.800 ;
        RECT 821.630 382.600 824.710 382.740 ;
        RECT 821.630 382.540 821.950 382.600 ;
        RECT 824.390 382.540 824.710 382.600 ;
        RECT 821.630 82.180 821.950 82.240 ;
        RECT 2071.450 82.180 2071.770 82.240 ;
        RECT 821.630 82.040 2071.770 82.180 ;
        RECT 821.630 81.980 821.950 82.040 ;
        RECT 2071.450 81.980 2071.770 82.040 ;
      LAYER via ;
        RECT 821.660 382.540 821.920 382.800 ;
        RECT 824.420 382.540 824.680 382.800 ;
        RECT 821.660 81.980 821.920 82.240 ;
        RECT 2071.480 81.980 2071.740 82.240 ;
      LAYER met2 ;
        RECT 825.690 400.250 825.970 404.000 ;
        RECT 824.480 400.110 825.970 400.250 ;
        RECT 824.480 382.830 824.620 400.110 ;
        RECT 825.690 400.000 825.970 400.110 ;
        RECT 821.660 382.510 821.920 382.830 ;
        RECT 824.420 382.510 824.680 382.830 ;
        RECT 821.720 82.270 821.860 382.510 ;
        RECT 821.660 81.950 821.920 82.270 ;
        RECT 2071.480 81.950 2071.740 82.270 ;
        RECT 2071.540 2.400 2071.680 81.950 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.990 81.840 829.310 81.900 ;
        RECT 2087.090 81.840 2087.410 81.900 ;
        RECT 828.990 81.700 2087.410 81.840 ;
        RECT 828.990 81.640 829.310 81.700 ;
        RECT 2087.090 81.640 2087.410 81.700 ;
      LAYER via ;
        RECT 829.020 81.640 829.280 81.900 ;
        RECT 2087.120 81.640 2087.380 81.900 ;
      LAYER met2 ;
        RECT 830.750 400.250 831.030 404.000 ;
        RECT 829.540 400.110 831.030 400.250 ;
        RECT 829.540 386.480 829.680 400.110 ;
        RECT 830.750 400.000 831.030 400.110 ;
        RECT 829.080 386.340 829.680 386.480 ;
        RECT 829.080 81.930 829.220 386.340 ;
        RECT 829.020 81.610 829.280 81.930 ;
        RECT 2087.120 81.610 2087.380 81.930 ;
        RECT 2087.180 1.770 2087.320 81.610 ;
        RECT 2089.270 1.770 2089.830 2.400 ;
        RECT 2087.180 1.630 2089.830 1.770 ;
        RECT 2089.270 -4.800 2089.830 1.630 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 834.970 81.500 835.290 81.560 ;
        RECT 2104.570 81.500 2104.890 81.560 ;
        RECT 834.970 81.360 2104.890 81.500 ;
        RECT 834.970 81.300 835.290 81.360 ;
        RECT 2104.570 81.300 2104.890 81.360 ;
      LAYER via ;
        RECT 835.000 81.300 835.260 81.560 ;
        RECT 2104.600 81.300 2104.860 81.560 ;
      LAYER met2 ;
        RECT 836.270 400.250 836.550 404.000 ;
        RECT 835.060 400.110 836.550 400.250 ;
        RECT 835.060 81.590 835.200 400.110 ;
        RECT 836.270 400.000 836.550 400.110 ;
        RECT 835.000 81.270 835.260 81.590 ;
        RECT 2104.600 81.270 2104.860 81.590 ;
        RECT 2104.660 1.770 2104.800 81.270 ;
        RECT 2106.750 1.770 2107.310 2.400 ;
        RECT 2104.660 1.630 2107.310 1.770 ;
        RECT 2106.750 -4.800 2107.310 1.630 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.430 376.280 835.750 376.340 ;
        RECT 840.490 376.280 840.810 376.340 ;
        RECT 835.430 376.140 840.810 376.280 ;
        RECT 835.430 376.080 835.750 376.140 ;
        RECT 840.490 376.080 840.810 376.140 ;
        RECT 835.430 81.160 835.750 81.220 ;
        RECT 2118.830 81.160 2119.150 81.220 ;
        RECT 835.430 81.020 2119.150 81.160 ;
        RECT 835.430 80.960 835.750 81.020 ;
        RECT 2118.830 80.960 2119.150 81.020 ;
        RECT 2118.830 15.880 2119.150 15.940 ;
        RECT 2124.810 15.880 2125.130 15.940 ;
        RECT 2118.830 15.740 2125.130 15.880 ;
        RECT 2118.830 15.680 2119.150 15.740 ;
        RECT 2124.810 15.680 2125.130 15.740 ;
      LAYER via ;
        RECT 835.460 376.080 835.720 376.340 ;
        RECT 840.520 376.080 840.780 376.340 ;
        RECT 835.460 80.960 835.720 81.220 ;
        RECT 2118.860 80.960 2119.120 81.220 ;
        RECT 2118.860 15.680 2119.120 15.940 ;
        RECT 2124.840 15.680 2125.100 15.940 ;
      LAYER met2 ;
        RECT 841.330 400.250 841.610 404.000 ;
        RECT 840.580 400.110 841.610 400.250 ;
        RECT 840.580 376.370 840.720 400.110 ;
        RECT 841.330 400.000 841.610 400.110 ;
        RECT 835.460 376.050 835.720 376.370 ;
        RECT 840.520 376.050 840.780 376.370 ;
        RECT 835.520 81.250 835.660 376.050 ;
        RECT 835.460 80.930 835.720 81.250 ;
        RECT 2118.860 80.930 2119.120 81.250 ;
        RECT 2118.920 15.970 2119.060 80.930 ;
        RECT 2118.860 15.650 2119.120 15.970 ;
        RECT 2124.840 15.650 2125.100 15.970 ;
        RECT 2124.900 2.400 2125.040 15.650 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.330 376.280 842.650 376.340 ;
        RECT 845.550 376.280 845.870 376.340 ;
        RECT 842.330 376.140 845.870 376.280 ;
        RECT 842.330 376.080 842.650 376.140 ;
        RECT 845.550 376.080 845.870 376.140 ;
        RECT 842.330 80.820 842.650 80.880 ;
        RECT 2142.290 80.820 2142.610 80.880 ;
        RECT 842.330 80.680 2142.610 80.820 ;
        RECT 842.330 80.620 842.650 80.680 ;
        RECT 2142.290 80.620 2142.610 80.680 ;
      LAYER via ;
        RECT 842.360 376.080 842.620 376.340 ;
        RECT 845.580 376.080 845.840 376.340 ;
        RECT 842.360 80.620 842.620 80.880 ;
        RECT 2142.320 80.620 2142.580 80.880 ;
      LAYER met2 ;
        RECT 846.850 400.250 847.130 404.000 ;
        RECT 845.640 400.110 847.130 400.250 ;
        RECT 845.640 376.370 845.780 400.110 ;
        RECT 846.850 400.000 847.130 400.110 ;
        RECT 842.360 376.050 842.620 376.370 ;
        RECT 845.580 376.050 845.840 376.370 ;
        RECT 842.420 80.910 842.560 376.050 ;
        RECT 842.360 80.590 842.620 80.910 ;
        RECT 2142.320 80.590 2142.580 80.910 ;
        RECT 2142.380 2.400 2142.520 80.590 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 849.690 376.280 850.010 376.340 ;
        RECT 851.070 376.280 851.390 376.340 ;
        RECT 849.690 376.140 851.390 376.280 ;
        RECT 849.690 376.080 850.010 376.140 ;
        RECT 851.070 376.080 851.390 376.140 ;
        RECT 849.690 80.480 850.010 80.540 ;
        RECT 2160.230 80.480 2160.550 80.540 ;
        RECT 849.690 80.340 2160.550 80.480 ;
        RECT 849.690 80.280 850.010 80.340 ;
        RECT 2160.230 80.280 2160.550 80.340 ;
      LAYER via ;
        RECT 849.720 376.080 849.980 376.340 ;
        RECT 851.100 376.080 851.360 376.340 ;
        RECT 849.720 80.280 849.980 80.540 ;
        RECT 2160.260 80.280 2160.520 80.540 ;
      LAYER met2 ;
        RECT 852.370 400.250 852.650 404.000 ;
        RECT 851.160 400.110 852.650 400.250 ;
        RECT 851.160 376.370 851.300 400.110 ;
        RECT 852.370 400.000 852.650 400.110 ;
        RECT 849.720 376.050 849.980 376.370 ;
        RECT 851.100 376.050 851.360 376.370 ;
        RECT 849.780 80.570 849.920 376.050 ;
        RECT 849.720 80.250 849.980 80.570 ;
        RECT 2160.260 80.250 2160.520 80.570 ;
        RECT 2160.320 2.400 2160.460 80.250 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.130 376.280 856.450 376.340 ;
        RECT 857.050 376.280 857.370 376.340 ;
        RECT 856.130 376.140 857.370 376.280 ;
        RECT 856.130 376.080 856.450 376.140 ;
        RECT 857.050 376.080 857.370 376.140 ;
        RECT 856.130 80.140 856.450 80.200 ;
        RECT 2175.410 80.140 2175.730 80.200 ;
        RECT 856.130 80.000 2175.730 80.140 ;
        RECT 856.130 79.940 856.450 80.000 ;
        RECT 2175.410 79.940 2175.730 80.000 ;
      LAYER via ;
        RECT 856.160 376.080 856.420 376.340 ;
        RECT 857.080 376.080 857.340 376.340 ;
        RECT 856.160 79.940 856.420 80.200 ;
        RECT 2175.440 79.940 2175.700 80.200 ;
      LAYER met2 ;
        RECT 857.430 400.250 857.710 404.000 ;
        RECT 857.140 400.110 857.710 400.250 ;
        RECT 857.140 376.370 857.280 400.110 ;
        RECT 857.430 400.000 857.710 400.110 ;
        RECT 856.160 376.050 856.420 376.370 ;
        RECT 857.080 376.050 857.340 376.370 ;
        RECT 856.220 80.230 856.360 376.050 ;
        RECT 856.160 79.910 856.420 80.230 ;
        RECT 2175.440 79.910 2175.700 80.230 ;
        RECT 2175.500 1.770 2175.640 79.910 ;
        RECT 2177.590 1.770 2178.150 2.400 ;
        RECT 2175.500 1.630 2178.150 1.770 ;
        RECT 2177.590 -4.800 2178.150 1.630 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.950 79.800 864.270 79.860 ;
        RECT 2195.650 79.800 2195.970 79.860 ;
        RECT 863.950 79.660 2195.970 79.800 ;
        RECT 863.950 79.600 864.270 79.660 ;
        RECT 2195.650 79.600 2195.970 79.660 ;
      LAYER via ;
        RECT 863.980 79.600 864.240 79.860 ;
        RECT 2195.680 79.600 2195.940 79.860 ;
      LAYER met2 ;
        RECT 862.950 400.250 863.230 404.000 ;
        RECT 862.950 400.110 864.180 400.250 ;
        RECT 862.950 400.000 863.230 400.110 ;
        RECT 864.040 79.890 864.180 400.110 ;
        RECT 863.980 79.570 864.240 79.890 ;
        RECT 2195.680 79.570 2195.940 79.890 ;
        RECT 2195.740 2.400 2195.880 79.570 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.490 376.280 863.810 376.340 ;
        RECT 867.170 376.280 867.490 376.340 ;
        RECT 863.490 376.140 867.490 376.280 ;
        RECT 863.490 376.080 863.810 376.140 ;
        RECT 867.170 376.080 867.490 376.140 ;
        RECT 863.490 79.460 863.810 79.520 ;
        RECT 2213.130 79.460 2213.450 79.520 ;
        RECT 863.490 79.320 2213.450 79.460 ;
        RECT 863.490 79.260 863.810 79.320 ;
        RECT 2213.130 79.260 2213.450 79.320 ;
      LAYER via ;
        RECT 863.520 376.080 863.780 376.340 ;
        RECT 867.200 376.080 867.460 376.340 ;
        RECT 863.520 79.260 863.780 79.520 ;
        RECT 2213.160 79.260 2213.420 79.520 ;
      LAYER met2 ;
        RECT 868.470 400.250 868.750 404.000 ;
        RECT 867.260 400.110 868.750 400.250 ;
        RECT 867.260 376.370 867.400 400.110 ;
        RECT 868.470 400.000 868.750 400.110 ;
        RECT 863.520 376.050 863.780 376.370 ;
        RECT 867.200 376.050 867.460 376.370 ;
        RECT 863.580 79.550 863.720 376.050 ;
        RECT 863.520 79.230 863.780 79.550 ;
        RECT 2213.160 79.230 2213.420 79.550 ;
        RECT 2213.220 2.400 2213.360 79.230 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 429.250 45.120 429.570 45.180 ;
        RECT 777.010 45.120 777.330 45.180 ;
        RECT 429.250 44.980 777.330 45.120 ;
        RECT 429.250 44.920 429.570 44.980 ;
        RECT 777.010 44.920 777.330 44.980 ;
      LAYER via ;
        RECT 429.280 44.920 429.540 45.180 ;
        RECT 777.040 44.920 777.300 45.180 ;
      LAYER met2 ;
        RECT 434.230 400.250 434.510 404.000 ;
        RECT 433.020 400.110 434.510 400.250 ;
        RECT 433.020 324.370 433.160 400.110 ;
        RECT 434.230 400.000 434.510 400.110 ;
        RECT 429.340 324.230 433.160 324.370 ;
        RECT 429.340 45.210 429.480 324.230 ;
        RECT 429.280 44.890 429.540 45.210 ;
        RECT 777.040 44.890 777.300 45.210 ;
        RECT 777.100 2.400 777.240 44.890 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.530 400.250 873.810 404.000 ;
        RECT 872.320 400.110 873.810 400.250 ;
        RECT 872.320 324.370 872.460 400.110 ;
        RECT 873.530 400.000 873.810 400.110 ;
        RECT 870.940 324.230 872.460 324.370 ;
        RECT 870.940 80.085 871.080 324.230 ;
        RECT 870.870 79.715 871.150 80.085 ;
        RECT 2228.790 79.715 2229.070 80.085 ;
        RECT 2228.860 1.770 2229.000 79.715 ;
        RECT 2230.950 1.770 2231.510 2.400 ;
        RECT 2228.860 1.630 2231.510 1.770 ;
        RECT 2230.950 -4.800 2231.510 1.630 ;
      LAYER via2 ;
        RECT 870.870 79.760 871.150 80.040 ;
        RECT 2228.790 79.760 2229.070 80.040 ;
      LAYER met3 ;
        RECT 870.845 80.050 871.175 80.065 ;
        RECT 2228.765 80.050 2229.095 80.065 ;
        RECT 870.845 79.750 2229.095 80.050 ;
        RECT 870.845 79.735 871.175 79.750 ;
        RECT 2228.765 79.735 2229.095 79.750 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2242.570 16.900 2242.890 16.960 ;
        RECT 2249.010 16.900 2249.330 16.960 ;
        RECT 2242.570 16.760 2249.330 16.900 ;
        RECT 2242.570 16.700 2242.890 16.760 ;
        RECT 2249.010 16.700 2249.330 16.760 ;
      LAYER via ;
        RECT 2242.600 16.700 2242.860 16.960 ;
        RECT 2249.040 16.700 2249.300 16.960 ;
      LAYER met2 ;
        RECT 879.050 400.250 879.330 404.000 ;
        RECT 877.840 400.110 879.330 400.250 ;
        RECT 877.840 79.405 877.980 400.110 ;
        RECT 879.050 400.000 879.330 400.110 ;
        RECT 877.770 79.035 878.050 79.405 ;
        RECT 2242.590 79.035 2242.870 79.405 ;
        RECT 2242.660 16.990 2242.800 79.035 ;
        RECT 2242.600 16.670 2242.860 16.990 ;
        RECT 2249.040 16.670 2249.300 16.990 ;
        RECT 2249.100 2.400 2249.240 16.670 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
      LAYER via2 ;
        RECT 877.770 79.080 878.050 79.360 ;
        RECT 2242.590 79.080 2242.870 79.360 ;
      LAYER met3 ;
        RECT 877.745 79.370 878.075 79.385 ;
        RECT 2242.565 79.370 2242.895 79.385 ;
        RECT 877.745 79.070 2242.895 79.370 ;
        RECT 877.745 79.055 878.075 79.070 ;
        RECT 2242.565 79.055 2242.895 79.070 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 884.650 122.300 884.970 122.360 ;
        RECT 2263.270 122.300 2263.590 122.360 ;
        RECT 884.650 122.160 2263.590 122.300 ;
        RECT 884.650 122.100 884.970 122.160 ;
        RECT 2263.270 122.100 2263.590 122.160 ;
      LAYER via ;
        RECT 884.680 122.100 884.940 122.360 ;
        RECT 2263.300 122.100 2263.560 122.360 ;
      LAYER met2 ;
        RECT 884.570 400.180 884.850 404.000 ;
        RECT 884.570 400.000 884.880 400.180 ;
        RECT 884.740 122.390 884.880 400.000 ;
        RECT 884.680 122.070 884.940 122.390 ;
        RECT 2263.300 122.070 2263.560 122.390 ;
        RECT 2263.360 82.870 2263.500 122.070 ;
        RECT 2263.360 82.730 2266.720 82.870 ;
        RECT 2266.580 2.400 2266.720 82.730 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 884.190 375.940 884.510 376.000 ;
        RECT 888.330 375.940 888.650 376.000 ;
        RECT 884.190 375.800 888.650 375.940 ;
        RECT 884.190 375.740 884.510 375.800 ;
        RECT 888.330 375.740 888.650 375.800 ;
        RECT 884.190 121.960 884.510 122.020 ;
        RECT 2284.430 121.960 2284.750 122.020 ;
        RECT 884.190 121.820 2284.750 121.960 ;
        RECT 884.190 121.760 884.510 121.820 ;
        RECT 2284.430 121.760 2284.750 121.820 ;
      LAYER via ;
        RECT 884.220 375.740 884.480 376.000 ;
        RECT 888.360 375.740 888.620 376.000 ;
        RECT 884.220 121.760 884.480 122.020 ;
        RECT 2284.460 121.760 2284.720 122.020 ;
      LAYER met2 ;
        RECT 889.630 400.250 889.910 404.000 ;
        RECT 888.420 400.110 889.910 400.250 ;
        RECT 888.420 376.030 888.560 400.110 ;
        RECT 889.630 400.000 889.910 400.110 ;
        RECT 884.220 375.710 884.480 376.030 ;
        RECT 888.360 375.710 888.620 376.030 ;
        RECT 884.280 122.050 884.420 375.710 ;
        RECT 884.220 121.730 884.480 122.050 ;
        RECT 2284.460 121.730 2284.720 122.050 ;
        RECT 2284.520 2.400 2284.660 121.730 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 891.090 121.620 891.410 121.680 ;
        RECT 2297.770 121.620 2298.090 121.680 ;
        RECT 891.090 121.480 2298.090 121.620 ;
        RECT 891.090 121.420 891.410 121.480 ;
        RECT 2297.770 121.420 2298.090 121.480 ;
      LAYER via ;
        RECT 891.120 121.420 891.380 121.680 ;
        RECT 2297.800 121.420 2298.060 121.680 ;
      LAYER met2 ;
        RECT 895.150 400.250 895.430 404.000 ;
        RECT 893.940 400.110 895.430 400.250 ;
        RECT 893.940 324.370 894.080 400.110 ;
        RECT 895.150 400.000 895.430 400.110 ;
        RECT 891.180 324.230 894.080 324.370 ;
        RECT 891.180 121.710 891.320 324.230 ;
        RECT 891.120 121.390 891.380 121.710 ;
        RECT 2297.800 121.390 2298.060 121.710 ;
        RECT 2297.860 82.870 2298.000 121.390 ;
        RECT 2297.860 82.730 2299.840 82.870 ;
        RECT 2299.700 1.770 2299.840 82.730 ;
        RECT 2301.790 1.770 2302.350 2.400 ;
        RECT 2299.700 1.630 2302.350 1.770 ;
        RECT 2301.790 -4.800 2302.350 1.630 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 898.450 121.280 898.770 121.340 ;
        RECT 2318.470 121.280 2318.790 121.340 ;
        RECT 898.450 121.140 2318.790 121.280 ;
        RECT 898.450 121.080 898.770 121.140 ;
        RECT 2318.470 121.080 2318.790 121.140 ;
      LAYER via ;
        RECT 898.480 121.080 898.740 121.340 ;
        RECT 2318.500 121.080 2318.760 121.340 ;
      LAYER met2 ;
        RECT 900.670 400.250 900.950 404.000 ;
        RECT 899.460 400.110 900.950 400.250 ;
        RECT 899.460 324.370 899.600 400.110 ;
        RECT 900.670 400.000 900.950 400.110 ;
        RECT 898.540 324.230 899.600 324.370 ;
        RECT 898.540 121.370 898.680 324.230 ;
        RECT 898.480 121.050 898.740 121.370 ;
        RECT 2318.500 121.050 2318.760 121.370 ;
        RECT 2318.560 82.870 2318.700 121.050 ;
        RECT 2318.560 82.730 2320.080 82.870 ;
        RECT 2319.940 2.400 2320.080 82.730 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 905.350 120.940 905.670 121.000 ;
        RECT 2332.270 120.940 2332.590 121.000 ;
        RECT 905.350 120.800 2332.590 120.940 ;
        RECT 905.350 120.740 905.670 120.800 ;
        RECT 2332.270 120.740 2332.590 120.800 ;
      LAYER via ;
        RECT 905.380 120.740 905.640 121.000 ;
        RECT 2332.300 120.740 2332.560 121.000 ;
      LAYER met2 ;
        RECT 905.730 400.250 906.010 404.000 ;
        RECT 905.440 400.110 906.010 400.250 ;
        RECT 905.440 121.030 905.580 400.110 ;
        RECT 905.730 400.000 906.010 400.110 ;
        RECT 905.380 120.710 905.640 121.030 ;
        RECT 2332.300 120.710 2332.560 121.030 ;
        RECT 2332.360 82.870 2332.500 120.710 ;
        RECT 2332.360 82.730 2337.560 82.870 ;
        RECT 2337.420 2.400 2337.560 82.730 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.790 84.900 912.110 84.960 ;
        RECT 2352.970 84.900 2353.290 84.960 ;
        RECT 911.790 84.760 2353.290 84.900 ;
        RECT 911.790 84.700 912.110 84.760 ;
        RECT 2352.970 84.700 2353.290 84.760 ;
      LAYER via ;
        RECT 911.820 84.700 912.080 84.960 ;
        RECT 2353.000 84.700 2353.260 84.960 ;
      LAYER met2 ;
        RECT 911.250 400.250 911.530 404.000 ;
        RECT 911.250 400.110 912.020 400.250 ;
        RECT 911.250 400.000 911.530 400.110 ;
        RECT 911.880 84.990 912.020 400.110 ;
        RECT 911.820 84.670 912.080 84.990 ;
        RECT 2353.000 84.670 2353.260 84.990 ;
        RECT 2353.060 1.770 2353.200 84.670 ;
        RECT 2355.150 1.770 2355.710 2.400 ;
        RECT 2353.060 1.630 2355.710 1.770 ;
        RECT 2355.150 -4.800 2355.710 1.630 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 912.250 85.240 912.570 85.300 ;
        RECT 2366.770 85.240 2367.090 85.300 ;
        RECT 912.250 85.100 2367.090 85.240 ;
        RECT 912.250 85.040 912.570 85.100 ;
        RECT 2366.770 85.040 2367.090 85.100 ;
        RECT 2366.770 17.580 2367.090 17.640 ;
        RECT 2370.910 17.580 2371.230 17.640 ;
        RECT 2366.770 17.440 2371.230 17.580 ;
        RECT 2366.770 17.380 2367.090 17.440 ;
        RECT 2370.910 17.380 2371.230 17.440 ;
      LAYER via ;
        RECT 912.280 85.040 912.540 85.300 ;
        RECT 2366.800 85.040 2367.060 85.300 ;
        RECT 2366.800 17.380 2367.060 17.640 ;
        RECT 2370.940 17.380 2371.200 17.640 ;
      LAYER met2 ;
        RECT 916.770 400.250 917.050 404.000 ;
        RECT 915.560 400.110 917.050 400.250 ;
        RECT 915.560 324.370 915.700 400.110 ;
        RECT 916.770 400.000 917.050 400.110 ;
        RECT 912.340 324.230 915.700 324.370 ;
        RECT 912.340 85.330 912.480 324.230 ;
        RECT 912.280 85.010 912.540 85.330 ;
        RECT 2366.800 85.010 2367.060 85.330 ;
        RECT 2366.860 17.670 2367.000 85.010 ;
        RECT 2366.800 17.350 2367.060 17.670 ;
        RECT 2370.940 17.350 2371.200 17.670 ;
        RECT 2371.000 1.770 2371.140 17.350 ;
        RECT 2372.630 1.770 2373.190 2.400 ;
        RECT 2371.000 1.630 2373.190 1.770 ;
        RECT 2372.630 -4.800 2373.190 1.630 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 919.150 85.580 919.470 85.640 ;
        RECT 2387.470 85.580 2387.790 85.640 ;
        RECT 919.150 85.440 2387.790 85.580 ;
        RECT 919.150 85.380 919.470 85.440 ;
        RECT 2387.470 85.380 2387.790 85.440 ;
      LAYER via ;
        RECT 919.180 85.380 919.440 85.640 ;
        RECT 2387.500 85.380 2387.760 85.640 ;
      LAYER met2 ;
        RECT 921.830 400.250 922.110 404.000 ;
        RECT 920.620 400.110 922.110 400.250 ;
        RECT 920.620 324.370 920.760 400.110 ;
        RECT 921.830 400.000 922.110 400.110 ;
        RECT 919.240 324.230 920.760 324.370 ;
        RECT 919.240 85.670 919.380 324.230 ;
        RECT 919.180 85.350 919.440 85.670 ;
        RECT 2387.500 85.350 2387.760 85.670 ;
        RECT 2387.560 82.870 2387.700 85.350 ;
        RECT 2387.560 82.730 2390.920 82.870 ;
        RECT 2390.780 2.400 2390.920 82.730 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.690 44.780 436.010 44.840 ;
        RECT 794.490 44.780 794.810 44.840 ;
        RECT 435.690 44.640 794.810 44.780 ;
        RECT 435.690 44.580 436.010 44.640 ;
        RECT 794.490 44.580 794.810 44.640 ;
      LAYER via ;
        RECT 435.720 44.580 435.980 44.840 ;
        RECT 794.520 44.580 794.780 44.840 ;
      LAYER met2 ;
        RECT 439.750 400.250 440.030 404.000 ;
        RECT 438.540 400.110 440.030 400.250 ;
        RECT 438.540 324.370 438.680 400.110 ;
        RECT 439.750 400.000 440.030 400.110 ;
        RECT 435.780 324.230 438.680 324.370 ;
        RECT 435.780 44.870 435.920 324.230 ;
        RECT 435.720 44.550 435.980 44.870 ;
        RECT 794.520 44.550 794.780 44.870 ;
        RECT 794.580 2.400 794.720 44.550 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.290 39.340 394.610 39.400 ;
        RECT 640.850 39.340 641.170 39.400 ;
        RECT 394.290 39.200 641.170 39.340 ;
        RECT 394.290 39.140 394.610 39.200 ;
        RECT 640.850 39.140 641.170 39.200 ;
      LAYER via ;
        RECT 394.320 39.140 394.580 39.400 ;
        RECT 640.880 39.140 641.140 39.400 ;
      LAYER met2 ;
        RECT 393.290 400.250 393.570 404.000 ;
        RECT 393.290 400.110 394.520 400.250 ;
        RECT 393.290 400.000 393.570 400.110 ;
        RECT 394.380 39.430 394.520 400.110 ;
        RECT 394.320 39.110 394.580 39.430 ;
        RECT 640.880 39.110 641.140 39.430 ;
        RECT 640.940 2.400 641.080 39.110 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.130 376.280 925.450 376.340 ;
        RECT 927.890 376.280 928.210 376.340 ;
        RECT 925.130 376.140 928.210 376.280 ;
        RECT 925.130 376.080 925.450 376.140 ;
        RECT 927.890 376.080 928.210 376.140 ;
        RECT 925.130 85.920 925.450 85.980 ;
        RECT 2408.170 85.920 2408.490 85.980 ;
        RECT 925.130 85.780 2408.490 85.920 ;
        RECT 925.130 85.720 925.450 85.780 ;
        RECT 2408.170 85.720 2408.490 85.780 ;
        RECT 2408.170 17.580 2408.490 17.640 ;
        RECT 2412.310 17.580 2412.630 17.640 ;
        RECT 2408.170 17.440 2412.630 17.580 ;
        RECT 2408.170 17.380 2408.490 17.440 ;
        RECT 2412.310 17.380 2412.630 17.440 ;
      LAYER via ;
        RECT 925.160 376.080 925.420 376.340 ;
        RECT 927.920 376.080 928.180 376.340 ;
        RECT 925.160 85.720 925.420 85.980 ;
        RECT 2408.200 85.720 2408.460 85.980 ;
        RECT 2408.200 17.380 2408.460 17.640 ;
        RECT 2412.340 17.380 2412.600 17.640 ;
      LAYER met2 ;
        RECT 929.190 400.250 929.470 404.000 ;
        RECT 927.980 400.110 929.470 400.250 ;
        RECT 927.980 376.370 928.120 400.110 ;
        RECT 929.190 400.000 929.470 400.110 ;
        RECT 925.160 376.050 925.420 376.370 ;
        RECT 927.920 376.050 928.180 376.370 ;
        RECT 925.220 86.010 925.360 376.050 ;
        RECT 925.160 85.690 925.420 86.010 ;
        RECT 2408.200 85.690 2408.460 86.010 ;
        RECT 2408.260 17.670 2408.400 85.690 ;
        RECT 2408.200 17.350 2408.460 17.670 ;
        RECT 2412.340 17.350 2412.600 17.670 ;
        RECT 2412.400 1.770 2412.540 17.350 ;
        RECT 2414.030 1.770 2414.590 2.400 ;
        RECT 2412.400 1.630 2414.590 1.770 ;
        RECT 2414.030 -4.800 2414.590 1.630 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.490 89.660 932.810 89.720 ;
        RECT 2428.870 89.660 2429.190 89.720 ;
        RECT 932.490 89.520 2429.190 89.660 ;
        RECT 932.490 89.460 932.810 89.520 ;
        RECT 2428.870 89.460 2429.190 89.520 ;
      LAYER via ;
        RECT 932.520 89.460 932.780 89.720 ;
        RECT 2428.900 89.460 2429.160 89.720 ;
      LAYER met2 ;
        RECT 934.250 400.250 934.530 404.000 ;
        RECT 933.500 400.110 934.530 400.250 ;
        RECT 933.500 351.970 933.640 400.110 ;
        RECT 934.250 400.000 934.530 400.110 ;
        RECT 932.580 351.830 933.640 351.970 ;
        RECT 932.580 89.750 932.720 351.830 ;
        RECT 932.520 89.430 932.780 89.750 ;
        RECT 2428.900 89.430 2429.160 89.750 ;
        RECT 2428.960 82.870 2429.100 89.430 ;
        RECT 2428.960 82.730 2432.320 82.870 ;
        RECT 2432.180 2.400 2432.320 82.730 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.930 89.320 939.250 89.380 ;
        RECT 2450.030 89.320 2450.350 89.380 ;
        RECT 938.930 89.180 2450.350 89.320 ;
        RECT 938.930 89.120 939.250 89.180 ;
        RECT 2450.030 89.120 2450.350 89.180 ;
      LAYER via ;
        RECT 938.960 89.120 939.220 89.380 ;
        RECT 2450.060 89.120 2450.320 89.380 ;
      LAYER met2 ;
        RECT 939.770 400.250 940.050 404.000 ;
        RECT 939.020 400.110 940.050 400.250 ;
        RECT 939.020 89.410 939.160 400.110 ;
        RECT 939.770 400.000 940.050 400.110 ;
        RECT 938.960 89.090 939.220 89.410 ;
        RECT 2450.060 89.090 2450.320 89.410 ;
        RECT 2450.120 16.730 2450.260 89.090 ;
        RECT 2449.660 16.590 2450.260 16.730 ;
        RECT 2449.660 2.400 2449.800 16.590 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.830 88.980 946.150 89.040 ;
        RECT 2463.370 88.980 2463.690 89.040 ;
        RECT 945.830 88.840 2463.690 88.980 ;
        RECT 945.830 88.780 946.150 88.840 ;
        RECT 2463.370 88.780 2463.690 88.840 ;
      LAYER via ;
        RECT 945.860 88.780 946.120 89.040 ;
        RECT 2463.400 88.780 2463.660 89.040 ;
      LAYER met2 ;
        RECT 945.290 400.250 945.570 404.000 ;
        RECT 945.290 400.110 946.060 400.250 ;
        RECT 945.290 400.000 945.570 400.110 ;
        RECT 945.920 89.070 946.060 400.110 ;
        RECT 945.860 88.750 946.120 89.070 ;
        RECT 2463.400 88.750 2463.660 89.070 ;
        RECT 2463.460 82.870 2463.600 88.750 ;
        RECT 2463.460 82.730 2465.440 82.870 ;
        RECT 2465.300 1.770 2465.440 82.730 ;
        RECT 2467.390 1.770 2467.950 2.400 ;
        RECT 2465.300 1.630 2467.950 1.770 ;
        RECT 2467.390 -4.800 2467.950 1.630 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.290 376.280 946.610 376.340 ;
        RECT 949.050 376.280 949.370 376.340 ;
        RECT 946.290 376.140 949.370 376.280 ;
        RECT 946.290 376.080 946.610 376.140 ;
        RECT 949.050 376.080 949.370 376.140 ;
        RECT 946.290 88.640 946.610 88.700 ;
        RECT 2484.070 88.640 2484.390 88.700 ;
        RECT 946.290 88.500 2484.390 88.640 ;
        RECT 946.290 88.440 946.610 88.500 ;
        RECT 2484.070 88.440 2484.390 88.500 ;
      LAYER via ;
        RECT 946.320 376.080 946.580 376.340 ;
        RECT 949.080 376.080 949.340 376.340 ;
        RECT 946.320 88.440 946.580 88.700 ;
        RECT 2484.100 88.440 2484.360 88.700 ;
      LAYER met2 ;
        RECT 950.350 400.250 950.630 404.000 ;
        RECT 949.140 400.110 950.630 400.250 ;
        RECT 949.140 376.370 949.280 400.110 ;
        RECT 950.350 400.000 950.630 400.110 ;
        RECT 946.320 376.050 946.580 376.370 ;
        RECT 949.080 376.050 949.340 376.370 ;
        RECT 946.380 88.730 946.520 376.050 ;
        RECT 946.320 88.410 946.580 88.730 ;
        RECT 2484.100 88.410 2484.360 88.730 ;
        RECT 2484.160 82.870 2484.300 88.410 ;
        RECT 2484.160 82.730 2485.680 82.870 ;
        RECT 2485.540 2.400 2485.680 82.730 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 953.650 88.300 953.970 88.360 ;
        RECT 2497.870 88.300 2498.190 88.360 ;
        RECT 953.650 88.160 2498.190 88.300 ;
        RECT 953.650 88.100 953.970 88.160 ;
        RECT 2497.870 88.100 2498.190 88.160 ;
      LAYER via ;
        RECT 953.680 88.100 953.940 88.360 ;
        RECT 2497.900 88.100 2498.160 88.360 ;
      LAYER met2 ;
        RECT 955.870 400.250 956.150 404.000 ;
        RECT 954.660 400.110 956.150 400.250 ;
        RECT 954.660 324.370 954.800 400.110 ;
        RECT 955.870 400.000 956.150 400.110 ;
        RECT 953.740 324.230 954.800 324.370 ;
        RECT 953.740 88.390 953.880 324.230 ;
        RECT 953.680 88.070 953.940 88.390 ;
        RECT 2497.900 88.070 2498.160 88.390 ;
        RECT 2497.960 82.870 2498.100 88.070 ;
        RECT 2497.960 82.730 2503.160 82.870 ;
        RECT 2503.020 2.400 2503.160 82.730 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.630 87.960 959.950 88.020 ;
        RECT 2518.570 87.960 2518.890 88.020 ;
        RECT 959.630 87.820 2518.890 87.960 ;
        RECT 959.630 87.760 959.950 87.820 ;
        RECT 2518.570 87.760 2518.890 87.820 ;
      LAYER via ;
        RECT 959.660 87.760 959.920 88.020 ;
        RECT 2518.600 87.760 2518.860 88.020 ;
      LAYER met2 ;
        RECT 961.390 400.250 961.670 404.000 ;
        RECT 960.180 400.110 961.670 400.250 ;
        RECT 960.180 392.090 960.320 400.110 ;
        RECT 961.390 400.000 961.670 400.110 ;
        RECT 959.720 391.950 960.320 392.090 ;
        RECT 959.720 88.050 959.860 391.950 ;
        RECT 959.660 87.730 959.920 88.050 ;
        RECT 2518.600 87.730 2518.860 88.050 ;
        RECT 2518.660 1.770 2518.800 87.730 ;
        RECT 2520.750 1.770 2521.310 2.400 ;
        RECT 2518.660 1.630 2521.310 1.770 ;
        RECT 2520.750 -4.800 2521.310 1.630 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.990 87.620 967.310 87.680 ;
        RECT 2532.830 87.620 2533.150 87.680 ;
        RECT 966.990 87.480 2533.150 87.620 ;
        RECT 966.990 87.420 967.310 87.480 ;
        RECT 2532.830 87.420 2533.150 87.480 ;
      LAYER via ;
        RECT 967.020 87.420 967.280 87.680 ;
        RECT 2532.860 87.420 2533.120 87.680 ;
      LAYER met2 ;
        RECT 966.450 400.250 966.730 404.000 ;
        RECT 966.450 400.110 967.220 400.250 ;
        RECT 966.450 400.000 966.730 400.110 ;
        RECT 967.080 87.710 967.220 400.110 ;
        RECT 967.020 87.390 967.280 87.710 ;
        RECT 2532.860 87.390 2533.120 87.710 ;
        RECT 2532.920 82.870 2533.060 87.390 ;
        RECT 2532.920 82.730 2536.280 82.870 ;
        RECT 2536.140 1.770 2536.280 82.730 ;
        RECT 2538.230 1.770 2538.790 2.400 ;
        RECT 2536.140 1.630 2538.790 1.770 ;
        RECT 2538.230 -4.800 2538.790 1.630 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.530 375.940 966.850 376.000 ;
        RECT 970.670 375.940 970.990 376.000 ;
        RECT 966.530 375.800 970.990 375.940 ;
        RECT 966.530 375.740 966.850 375.800 ;
        RECT 970.670 375.740 970.990 375.800 ;
        RECT 966.530 87.280 966.850 87.340 ;
        RECT 2553.070 87.280 2553.390 87.340 ;
        RECT 966.530 87.140 2553.390 87.280 ;
        RECT 966.530 87.080 966.850 87.140 ;
        RECT 2553.070 87.080 2553.390 87.140 ;
      LAYER via ;
        RECT 966.560 375.740 966.820 376.000 ;
        RECT 970.700 375.740 970.960 376.000 ;
        RECT 966.560 87.080 966.820 87.340 ;
        RECT 2553.100 87.080 2553.360 87.340 ;
      LAYER met2 ;
        RECT 971.970 400.250 972.250 404.000 ;
        RECT 970.760 400.110 972.250 400.250 ;
        RECT 970.760 376.030 970.900 400.110 ;
        RECT 971.970 400.000 972.250 400.110 ;
        RECT 966.560 375.710 966.820 376.030 ;
        RECT 970.700 375.710 970.960 376.030 ;
        RECT 966.620 87.370 966.760 375.710 ;
        RECT 966.560 87.050 966.820 87.370 ;
        RECT 2553.100 87.050 2553.360 87.370 ;
        RECT 2553.160 82.870 2553.300 87.050 ;
        RECT 2553.160 82.730 2556.520 82.870 ;
        RECT 2556.380 2.400 2556.520 82.730 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.890 376.280 974.210 376.340 ;
        RECT 976.190 376.280 976.510 376.340 ;
        RECT 973.890 376.140 976.510 376.280 ;
        RECT 973.890 376.080 974.210 376.140 ;
        RECT 976.190 376.080 976.510 376.140 ;
        RECT 973.890 86.940 974.210 87.000 ;
        RECT 2573.770 86.940 2574.090 87.000 ;
        RECT 973.890 86.800 2574.090 86.940 ;
        RECT 973.890 86.740 974.210 86.800 ;
        RECT 2573.770 86.740 2574.090 86.800 ;
      LAYER via ;
        RECT 973.920 376.080 974.180 376.340 ;
        RECT 976.220 376.080 976.480 376.340 ;
        RECT 973.920 86.740 974.180 87.000 ;
        RECT 2573.800 86.740 2574.060 87.000 ;
      LAYER met2 ;
        RECT 977.490 400.250 977.770 404.000 ;
        RECT 976.280 400.110 977.770 400.250 ;
        RECT 976.280 376.370 976.420 400.110 ;
        RECT 977.490 400.000 977.770 400.110 ;
        RECT 973.920 376.050 974.180 376.370 ;
        RECT 976.220 376.050 976.480 376.370 ;
        RECT 973.980 87.030 974.120 376.050 ;
        RECT 973.920 86.710 974.180 87.030 ;
        RECT 2573.800 86.710 2574.060 87.030 ;
        RECT 2573.860 2.400 2574.000 86.710 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 39.680 443.370 39.740 ;
        RECT 651.430 39.680 651.750 39.740 ;
        RECT 443.050 39.540 651.750 39.680 ;
        RECT 443.050 39.480 443.370 39.540 ;
        RECT 651.430 39.480 651.750 39.540 ;
        RECT 651.430 18.940 651.750 19.000 ;
        RECT 818.410 18.940 818.730 19.000 ;
        RECT 651.430 18.800 818.730 18.940 ;
        RECT 651.430 18.740 651.750 18.800 ;
        RECT 818.410 18.740 818.730 18.800 ;
      LAYER via ;
        RECT 443.080 39.480 443.340 39.740 ;
        RECT 651.460 39.480 651.720 39.740 ;
        RECT 651.460 18.740 651.720 19.000 ;
        RECT 818.440 18.740 818.700 19.000 ;
      LAYER met2 ;
        RECT 446.650 400.250 446.930 404.000 ;
        RECT 445.440 400.110 446.930 400.250 ;
        RECT 445.440 387.330 445.580 400.110 ;
        RECT 446.650 400.000 446.930 400.110 ;
        RECT 443.140 387.190 445.580 387.330 ;
        RECT 443.140 39.770 443.280 387.190 ;
        RECT 443.080 39.450 443.340 39.770 ;
        RECT 651.460 39.450 651.720 39.770 ;
        RECT 651.520 19.030 651.660 39.450 ;
        RECT 651.460 18.710 651.720 19.030 ;
        RECT 818.440 18.710 818.700 19.030 ;
        RECT 818.500 2.400 818.640 18.710 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 981.250 86.600 981.570 86.660 ;
        RECT 2587.570 86.600 2587.890 86.660 ;
        RECT 981.250 86.460 2587.890 86.600 ;
        RECT 981.250 86.400 981.570 86.460 ;
        RECT 2587.570 86.400 2587.890 86.460 ;
      LAYER via ;
        RECT 981.280 86.400 981.540 86.660 ;
        RECT 2587.600 86.400 2587.860 86.660 ;
      LAYER met2 ;
        RECT 982.550 400.250 982.830 404.000 ;
        RECT 981.340 400.110 982.830 400.250 ;
        RECT 981.340 86.690 981.480 400.110 ;
        RECT 982.550 400.000 982.830 400.110 ;
        RECT 981.280 86.370 981.540 86.690 ;
        RECT 2587.600 86.370 2587.860 86.690 ;
        RECT 2587.660 82.870 2587.800 86.370 ;
        RECT 2587.660 82.730 2589.640 82.870 ;
        RECT 2589.500 1.770 2589.640 82.730 ;
        RECT 2591.590 1.770 2592.150 2.400 ;
        RECT 2589.500 1.630 2592.150 1.770 ;
        RECT 2591.590 -4.800 2592.150 1.630 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.690 86.260 988.010 86.320 ;
        RECT 2608.270 86.260 2608.590 86.320 ;
        RECT 987.690 86.120 2608.590 86.260 ;
        RECT 987.690 86.060 988.010 86.120 ;
        RECT 2608.270 86.060 2608.590 86.120 ;
      LAYER via ;
        RECT 987.720 86.060 987.980 86.320 ;
        RECT 2608.300 86.060 2608.560 86.320 ;
      LAYER met2 ;
        RECT 988.070 400.250 988.350 404.000 ;
        RECT 987.780 400.110 988.350 400.250 ;
        RECT 987.780 86.350 987.920 400.110 ;
        RECT 988.070 400.000 988.350 400.110 ;
        RECT 987.720 86.030 987.980 86.350 ;
        RECT 2608.300 86.030 2608.560 86.350 ;
        RECT 2608.360 1.770 2608.500 86.030 ;
        RECT 2609.070 1.770 2609.630 2.400 ;
        RECT 2608.360 1.630 2609.630 1.770 ;
        RECT 2609.070 -4.800 2609.630 1.630 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.590 387.840 994.910 387.900 ;
        RECT 995.970 387.840 996.290 387.900 ;
        RECT 994.590 387.700 996.290 387.840 ;
        RECT 994.590 387.640 994.910 387.700 ;
        RECT 995.970 387.640 996.290 387.700 ;
      LAYER via ;
        RECT 994.620 387.640 994.880 387.900 ;
        RECT 996.000 387.640 996.260 387.900 ;
      LAYER met2 ;
        RECT 993.590 400.250 993.870 404.000 ;
        RECT 993.590 400.110 994.820 400.250 ;
        RECT 993.590 400.000 993.870 400.110 ;
        RECT 994.680 387.930 994.820 400.110 ;
        RECT 994.620 387.610 994.880 387.930 ;
        RECT 996.000 387.610 996.260 387.930 ;
        RECT 996.060 384.610 996.200 387.610 ;
        RECT 994.680 384.470 996.200 384.610 ;
        RECT 994.680 86.885 994.820 384.470 ;
        RECT 994.610 86.515 994.890 86.885 ;
        RECT 2622.090 86.515 2622.370 86.885 ;
        RECT 2622.160 82.870 2622.300 86.515 ;
        RECT 2622.160 82.730 2627.360 82.870 ;
        RECT 2627.220 2.400 2627.360 82.730 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
      LAYER via2 ;
        RECT 994.610 86.560 994.890 86.840 ;
        RECT 2622.090 86.560 2622.370 86.840 ;
      LAYER met3 ;
        RECT 994.585 86.850 994.915 86.865 ;
        RECT 2622.065 86.850 2622.395 86.865 ;
        RECT 994.585 86.550 2622.395 86.850 ;
        RECT 994.585 86.535 994.915 86.550 ;
        RECT 2622.065 86.535 2622.395 86.550 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.650 400.250 998.930 404.000 ;
        RECT 997.440 400.110 998.930 400.250 ;
        RECT 997.440 324.370 997.580 400.110 ;
        RECT 998.650 400.000 998.930 400.110 ;
        RECT 995.600 324.230 997.580 324.370 ;
        RECT 995.600 86.205 995.740 324.230 ;
        RECT 995.530 85.835 995.810 86.205 ;
        RECT 2642.790 85.835 2643.070 86.205 ;
        RECT 2642.860 1.770 2643.000 85.835 ;
        RECT 2644.950 1.770 2645.510 2.400 ;
        RECT 2642.860 1.630 2645.510 1.770 ;
        RECT 2644.950 -4.800 2645.510 1.630 ;
      LAYER via2 ;
        RECT 995.530 85.880 995.810 86.160 ;
        RECT 2642.790 85.880 2643.070 86.160 ;
      LAYER met3 ;
        RECT 995.505 86.170 995.835 86.185 ;
        RECT 2642.765 86.170 2643.095 86.185 ;
        RECT 995.505 85.870 2643.095 86.170 ;
        RECT 995.505 85.855 995.835 85.870 ;
        RECT 2642.765 85.855 2643.095 85.870 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.950 120.600 1002.270 120.660 ;
        RECT 2656.570 120.600 2656.890 120.660 ;
        RECT 1001.950 120.460 2656.890 120.600 ;
        RECT 1001.950 120.400 1002.270 120.460 ;
        RECT 2656.570 120.400 2656.890 120.460 ;
        RECT 2656.570 17.580 2656.890 17.640 ;
        RECT 2660.710 17.580 2661.030 17.640 ;
        RECT 2656.570 17.440 2661.030 17.580 ;
        RECT 2656.570 17.380 2656.890 17.440 ;
        RECT 2660.710 17.380 2661.030 17.440 ;
      LAYER via ;
        RECT 1001.980 120.400 1002.240 120.660 ;
        RECT 2656.600 120.400 2656.860 120.660 ;
        RECT 2656.600 17.380 2656.860 17.640 ;
        RECT 2660.740 17.380 2661.000 17.640 ;
      LAYER met2 ;
        RECT 1004.170 400.250 1004.450 404.000 ;
        RECT 1002.960 400.110 1004.450 400.250 ;
        RECT 1002.960 324.370 1003.100 400.110 ;
        RECT 1004.170 400.000 1004.450 400.110 ;
        RECT 1002.040 324.230 1003.100 324.370 ;
        RECT 1002.040 120.690 1002.180 324.230 ;
        RECT 1001.980 120.370 1002.240 120.690 ;
        RECT 2656.600 120.370 2656.860 120.690 ;
        RECT 2656.660 17.670 2656.800 120.370 ;
        RECT 2656.600 17.350 2656.860 17.670 ;
        RECT 2660.740 17.350 2661.000 17.670 ;
        RECT 2660.800 1.770 2660.940 17.350 ;
        RECT 2662.430 1.770 2662.990 2.400 ;
        RECT 2660.800 1.630 2662.990 1.770 ;
        RECT 2662.430 -4.800 2662.990 1.630 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.230 400.250 1009.510 404.000 ;
        RECT 1008.940 400.110 1009.510 400.250 ;
        RECT 1008.940 121.565 1009.080 400.110 ;
        RECT 1009.230 400.000 1009.510 400.110 ;
        RECT 1008.870 121.195 1009.150 121.565 ;
        RECT 2677.290 121.195 2677.570 121.565 ;
        RECT 2677.360 82.870 2677.500 121.195 ;
        RECT 2677.360 82.730 2680.720 82.870 ;
        RECT 2680.580 2.400 2680.720 82.730 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
      LAYER via2 ;
        RECT 1008.870 121.240 1009.150 121.520 ;
        RECT 2677.290 121.240 2677.570 121.520 ;
      LAYER met3 ;
        RECT 1008.845 121.530 1009.175 121.545 ;
        RECT 2677.265 121.530 2677.595 121.545 ;
        RECT 1008.845 121.230 2677.595 121.530 ;
        RECT 1008.845 121.215 1009.175 121.230 ;
        RECT 2677.265 121.215 2677.595 121.230 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.750 400.250 1015.030 404.000 ;
        RECT 1014.750 400.110 1015.520 400.250 ;
        RECT 1014.750 400.000 1015.030 400.110 ;
        RECT 1015.380 120.885 1015.520 400.110 ;
        RECT 1015.310 120.515 1015.590 120.885 ;
        RECT 2697.990 120.515 2698.270 120.885 ;
        RECT 2698.060 2.400 2698.200 120.515 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
      LAYER via2 ;
        RECT 1015.310 120.560 1015.590 120.840 ;
        RECT 2697.990 120.560 2698.270 120.840 ;
      LAYER met3 ;
        RECT 1015.285 120.850 1015.615 120.865 ;
        RECT 2697.965 120.850 2698.295 120.865 ;
        RECT 1015.285 120.550 2698.295 120.850 ;
        RECT 1015.285 120.535 1015.615 120.550 ;
        RECT 2697.965 120.535 2698.295 120.550 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.270 400.250 1020.550 404.000 ;
        RECT 1019.060 400.110 1020.550 400.250 ;
        RECT 1019.060 324.370 1019.200 400.110 ;
        RECT 1020.270 400.000 1020.550 400.110 ;
        RECT 1015.840 324.230 1019.200 324.370 ;
        RECT 1015.840 127.685 1015.980 324.230 ;
        RECT 1015.770 127.315 1016.050 127.685 ;
        RECT 2711.790 127.315 2712.070 127.685 ;
        RECT 2711.860 82.870 2712.000 127.315 ;
        RECT 2711.860 82.730 2713.840 82.870 ;
        RECT 2713.700 1.770 2713.840 82.730 ;
        RECT 2715.790 1.770 2716.350 2.400 ;
        RECT 2713.700 1.630 2716.350 1.770 ;
        RECT 2715.790 -4.800 2716.350 1.630 ;
      LAYER via2 ;
        RECT 1015.770 127.360 1016.050 127.640 ;
        RECT 2711.790 127.360 2712.070 127.640 ;
      LAYER met3 ;
        RECT 1015.745 127.650 1016.075 127.665 ;
        RECT 2711.765 127.650 2712.095 127.665 ;
        RECT 1015.745 127.350 2712.095 127.650 ;
        RECT 1015.745 127.335 1016.075 127.350 ;
        RECT 2711.765 127.335 2712.095 127.350 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.650 95.440 1022.970 95.500 ;
        RECT 2732.470 95.440 2732.790 95.500 ;
        RECT 1022.650 95.300 2732.790 95.440 ;
        RECT 1022.650 95.240 1022.970 95.300 ;
        RECT 2732.470 95.240 2732.790 95.300 ;
      LAYER via ;
        RECT 1022.680 95.240 1022.940 95.500 ;
        RECT 2732.500 95.240 2732.760 95.500 ;
      LAYER met2 ;
        RECT 1025.330 400.250 1025.610 404.000 ;
        RECT 1024.580 400.110 1025.610 400.250 ;
        RECT 1024.580 324.370 1024.720 400.110 ;
        RECT 1025.330 400.000 1025.610 400.110 ;
        RECT 1022.740 324.230 1024.720 324.370 ;
        RECT 1022.740 95.530 1022.880 324.230 ;
        RECT 1022.680 95.210 1022.940 95.530 ;
        RECT 2732.500 95.210 2732.760 95.530 ;
        RECT 2732.560 1.770 2732.700 95.210 ;
        RECT 2733.270 1.770 2733.830 2.400 ;
        RECT 2732.560 1.630 2733.830 1.770 ;
        RECT 2733.270 -4.800 2733.830 1.630 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1029.550 95.100 1029.870 95.160 ;
        RECT 2746.270 95.100 2746.590 95.160 ;
        RECT 1029.550 94.960 2746.590 95.100 ;
        RECT 1029.550 94.900 1029.870 94.960 ;
        RECT 2746.270 94.900 2746.590 94.960 ;
      LAYER via ;
        RECT 1029.580 94.900 1029.840 95.160 ;
        RECT 2746.300 94.900 2746.560 95.160 ;
      LAYER met2 ;
        RECT 1030.850 400.250 1031.130 404.000 ;
        RECT 1029.640 400.110 1031.130 400.250 ;
        RECT 1029.640 95.190 1029.780 400.110 ;
        RECT 1030.850 400.000 1031.130 400.110 ;
        RECT 1029.580 94.870 1029.840 95.190 ;
        RECT 2746.300 94.870 2746.560 95.190 ;
        RECT 2746.360 82.870 2746.500 94.870 ;
        RECT 2746.360 82.730 2751.560 82.870 ;
        RECT 2751.420 2.400 2751.560 82.730 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.490 53.960 449.810 54.020 ;
        RECT 835.890 53.960 836.210 54.020 ;
        RECT 449.490 53.820 836.210 53.960 ;
        RECT 449.490 53.760 449.810 53.820 ;
        RECT 835.890 53.760 836.210 53.820 ;
      LAYER via ;
        RECT 449.520 53.760 449.780 54.020 ;
        RECT 835.920 53.760 836.180 54.020 ;
      LAYER met2 ;
        RECT 452.170 400.250 452.450 404.000 ;
        RECT 450.960 400.110 452.450 400.250 ;
        RECT 450.960 324.370 451.100 400.110 ;
        RECT 452.170 400.000 452.450 400.110 ;
        RECT 449.580 324.230 451.100 324.370 ;
        RECT 449.580 54.050 449.720 324.230 ;
        RECT 449.520 53.730 449.780 54.050 ;
        RECT 835.920 53.730 836.180 54.050 ;
        RECT 835.980 2.400 836.120 53.730 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1036.450 94.760 1036.770 94.820 ;
        RECT 2766.970 94.760 2767.290 94.820 ;
        RECT 1036.450 94.620 2767.290 94.760 ;
        RECT 1036.450 94.560 1036.770 94.620 ;
        RECT 2766.970 94.560 2767.290 94.620 ;
      LAYER via ;
        RECT 1036.480 94.560 1036.740 94.820 ;
        RECT 2767.000 94.560 2767.260 94.820 ;
      LAYER met2 ;
        RECT 1036.370 400.180 1036.650 404.000 ;
        RECT 1036.370 400.000 1036.680 400.180 ;
        RECT 1036.540 94.850 1036.680 400.000 ;
        RECT 1036.480 94.530 1036.740 94.850 ;
        RECT 2767.000 94.530 2767.260 94.850 ;
        RECT 2767.060 82.870 2767.200 94.530 ;
        RECT 2767.060 82.730 2769.040 82.870 ;
        RECT 2768.900 2.400 2769.040 82.730 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.990 375.940 1036.310 376.000 ;
        RECT 1040.130 375.940 1040.450 376.000 ;
        RECT 1035.990 375.800 1040.450 375.940 ;
        RECT 1035.990 375.740 1036.310 375.800 ;
        RECT 1040.130 375.740 1040.450 375.800 ;
        RECT 1035.990 94.420 1036.310 94.480 ;
        RECT 2780.770 94.420 2781.090 94.480 ;
        RECT 1035.990 94.280 2781.090 94.420 ;
        RECT 1035.990 94.220 1036.310 94.280 ;
        RECT 2780.770 94.220 2781.090 94.280 ;
        RECT 2780.770 17.580 2781.090 17.640 ;
        RECT 2784.910 17.580 2785.230 17.640 ;
        RECT 2780.770 17.440 2785.230 17.580 ;
        RECT 2780.770 17.380 2781.090 17.440 ;
        RECT 2784.910 17.380 2785.230 17.440 ;
      LAYER via ;
        RECT 1036.020 375.740 1036.280 376.000 ;
        RECT 1040.160 375.740 1040.420 376.000 ;
        RECT 1036.020 94.220 1036.280 94.480 ;
        RECT 2780.800 94.220 2781.060 94.480 ;
        RECT 2780.800 17.380 2781.060 17.640 ;
        RECT 2784.940 17.380 2785.200 17.640 ;
      LAYER met2 ;
        RECT 1041.430 400.250 1041.710 404.000 ;
        RECT 1040.220 400.110 1041.710 400.250 ;
        RECT 1040.220 376.030 1040.360 400.110 ;
        RECT 1041.430 400.000 1041.710 400.110 ;
        RECT 1036.020 375.710 1036.280 376.030 ;
        RECT 1040.160 375.710 1040.420 376.030 ;
        RECT 1036.080 94.510 1036.220 375.710 ;
        RECT 1036.020 94.190 1036.280 94.510 ;
        RECT 2780.800 94.190 2781.060 94.510 ;
        RECT 2780.860 17.670 2781.000 94.190 ;
        RECT 2780.800 17.350 2781.060 17.670 ;
        RECT 2784.940 17.350 2785.200 17.670 ;
        RECT 2785.000 1.770 2785.140 17.350 ;
        RECT 2786.630 1.770 2787.190 2.400 ;
        RECT 2785.000 1.630 2787.190 1.770 ;
        RECT 2786.630 -4.800 2787.190 1.630 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.430 376.280 1042.750 376.340 ;
        RECT 1045.650 376.280 1045.970 376.340 ;
        RECT 1042.430 376.140 1045.970 376.280 ;
        RECT 1042.430 376.080 1042.750 376.140 ;
        RECT 1045.650 376.080 1045.970 376.140 ;
        RECT 1042.430 94.080 1042.750 94.140 ;
        RECT 2801.470 94.080 2801.790 94.140 ;
        RECT 1042.430 93.940 2801.790 94.080 ;
        RECT 1042.430 93.880 1042.750 93.940 ;
        RECT 2801.470 93.880 2801.790 93.940 ;
      LAYER via ;
        RECT 1042.460 376.080 1042.720 376.340 ;
        RECT 1045.680 376.080 1045.940 376.340 ;
        RECT 1042.460 93.880 1042.720 94.140 ;
        RECT 2801.500 93.880 2801.760 94.140 ;
      LAYER met2 ;
        RECT 1046.950 400.250 1047.230 404.000 ;
        RECT 1045.740 400.110 1047.230 400.250 ;
        RECT 1045.740 376.370 1045.880 400.110 ;
        RECT 1046.950 400.000 1047.230 400.110 ;
        RECT 1042.460 376.050 1042.720 376.370 ;
        RECT 1045.680 376.050 1045.940 376.370 ;
        RECT 1042.520 94.170 1042.660 376.050 ;
        RECT 1042.460 93.850 1042.720 94.170 ;
        RECT 2801.500 93.850 2801.760 94.170 ;
        RECT 2801.560 82.870 2801.700 93.850 ;
        RECT 2801.560 82.730 2802.160 82.870 ;
        RECT 2802.020 1.770 2802.160 82.730 ;
        RECT 2804.110 1.770 2804.670 2.400 ;
        RECT 2802.020 1.630 2804.670 1.770 ;
        RECT 2804.110 -4.800 2804.670 1.630 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.330 376.280 1049.650 376.340 ;
        RECT 1051.170 376.280 1051.490 376.340 ;
        RECT 1049.330 376.140 1051.490 376.280 ;
        RECT 1049.330 376.080 1049.650 376.140 ;
        RECT 1051.170 376.080 1051.490 376.140 ;
        RECT 1049.330 93.740 1049.650 93.800 ;
        RECT 2822.630 93.740 2822.950 93.800 ;
        RECT 1049.330 93.600 2822.950 93.740 ;
        RECT 1049.330 93.540 1049.650 93.600 ;
        RECT 2822.630 93.540 2822.950 93.600 ;
      LAYER via ;
        RECT 1049.360 376.080 1049.620 376.340 ;
        RECT 1051.200 376.080 1051.460 376.340 ;
        RECT 1049.360 93.540 1049.620 93.800 ;
        RECT 2822.660 93.540 2822.920 93.800 ;
      LAYER met2 ;
        RECT 1052.470 400.250 1052.750 404.000 ;
        RECT 1051.260 400.110 1052.750 400.250 ;
        RECT 1051.260 376.370 1051.400 400.110 ;
        RECT 1052.470 400.000 1052.750 400.110 ;
        RECT 1049.360 376.050 1049.620 376.370 ;
        RECT 1051.200 376.050 1051.460 376.370 ;
        RECT 1049.420 93.830 1049.560 376.050 ;
        RECT 1049.360 93.510 1049.620 93.830 ;
        RECT 2822.660 93.510 2822.920 93.830 ;
        RECT 2822.720 16.730 2822.860 93.510 ;
        RECT 2822.260 16.590 2822.860 16.730 ;
        RECT 2822.260 2.400 2822.400 16.590 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1056.690 93.400 1057.010 93.460 ;
        RECT 2835.970 93.400 2836.290 93.460 ;
        RECT 1056.690 93.260 2836.290 93.400 ;
        RECT 1056.690 93.200 1057.010 93.260 ;
        RECT 2835.970 93.200 2836.290 93.260 ;
      LAYER via ;
        RECT 1056.720 93.200 1056.980 93.460 ;
        RECT 2836.000 93.200 2836.260 93.460 ;
      LAYER met2 ;
        RECT 1057.530 400.250 1057.810 404.000 ;
        RECT 1056.780 400.110 1057.810 400.250 ;
        RECT 1056.780 93.490 1056.920 400.110 ;
        RECT 1057.530 400.000 1057.810 400.110 ;
        RECT 1056.720 93.170 1056.980 93.490 ;
        RECT 2836.000 93.170 2836.260 93.490 ;
        RECT 2836.060 82.870 2836.200 93.170 ;
        RECT 2836.060 82.730 2838.040 82.870 ;
        RECT 2837.900 1.770 2838.040 82.730 ;
        RECT 2839.990 1.770 2840.550 2.400 ;
        RECT 2837.900 1.630 2840.550 1.770 ;
        RECT 2839.990 -4.800 2840.550 1.630 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.590 93.060 1063.910 93.120 ;
        RECT 2856.670 93.060 2856.990 93.120 ;
        RECT 1063.590 92.920 2856.990 93.060 ;
        RECT 1063.590 92.860 1063.910 92.920 ;
        RECT 2856.670 92.860 2856.990 92.920 ;
      LAYER via ;
        RECT 1063.620 92.860 1063.880 93.120 ;
        RECT 2856.700 92.860 2856.960 93.120 ;
      LAYER met2 ;
        RECT 1063.050 400.250 1063.330 404.000 ;
        RECT 1063.050 400.110 1063.820 400.250 ;
        RECT 1063.050 400.000 1063.330 400.110 ;
        RECT 1063.680 93.150 1063.820 400.110 ;
        RECT 1063.620 92.830 1063.880 93.150 ;
        RECT 2856.700 92.830 2856.960 93.150 ;
        RECT 2856.760 1.770 2856.900 92.830 ;
        RECT 2857.470 1.770 2858.030 2.400 ;
        RECT 2856.760 1.630 2858.030 1.770 ;
        RECT 2857.470 -4.800 2858.030 1.630 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.570 400.250 1068.850 404.000 ;
        RECT 1067.360 400.110 1068.850 400.250 ;
        RECT 1067.360 324.370 1067.500 400.110 ;
        RECT 1068.570 400.000 1068.850 400.110 ;
        RECT 1064.140 324.230 1067.500 324.370 ;
        RECT 1064.140 93.685 1064.280 324.230 ;
        RECT 1064.070 93.315 1064.350 93.685 ;
        RECT 2870.490 93.315 2870.770 93.685 ;
        RECT 2870.560 82.870 2870.700 93.315 ;
        RECT 2870.560 82.730 2875.760 82.870 ;
        RECT 2875.620 2.400 2875.760 82.730 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
      LAYER via2 ;
        RECT 1064.070 93.360 1064.350 93.640 ;
        RECT 2870.490 93.360 2870.770 93.640 ;
      LAYER met3 ;
        RECT 1064.045 93.650 1064.375 93.665 ;
        RECT 2870.465 93.650 2870.795 93.665 ;
        RECT 1064.045 93.350 2870.795 93.650 ;
        RECT 1064.045 93.335 1064.375 93.350 ;
        RECT 2870.465 93.335 2870.795 93.350 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.630 400.250 1073.910 404.000 ;
        RECT 1072.420 400.110 1073.910 400.250 ;
        RECT 1072.420 324.370 1072.560 400.110 ;
        RECT 1073.630 400.000 1073.910 400.110 ;
        RECT 1071.500 324.230 1072.560 324.370 ;
        RECT 1071.500 93.005 1071.640 324.230 ;
        RECT 1071.430 92.635 1071.710 93.005 ;
        RECT 2891.190 92.635 2891.470 93.005 ;
        RECT 2891.260 82.870 2891.400 92.635 ;
        RECT 2891.260 82.730 2893.240 82.870 ;
        RECT 2893.100 2.400 2893.240 82.730 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 1071.430 92.680 1071.710 92.960 ;
        RECT 2891.190 92.680 2891.470 92.960 ;
      LAYER met3 ;
        RECT 1071.405 92.970 1071.735 92.985 ;
        RECT 2891.165 92.970 2891.495 92.985 ;
        RECT 1071.405 92.670 2891.495 92.970 ;
        RECT 1071.405 92.655 1071.735 92.670 ;
        RECT 2891.165 92.655 2891.495 92.670 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.930 53.620 456.250 53.680 ;
        RECT 851.530 53.620 851.850 53.680 ;
        RECT 455.930 53.480 851.850 53.620 ;
        RECT 455.930 53.420 456.250 53.480 ;
        RECT 851.530 53.420 851.850 53.480 ;
      LAYER via ;
        RECT 455.960 53.420 456.220 53.680 ;
        RECT 851.560 53.420 851.820 53.680 ;
      LAYER met2 ;
        RECT 457.690 400.250 457.970 404.000 ;
        RECT 456.480 400.110 457.970 400.250 ;
        RECT 456.480 386.480 456.620 400.110 ;
        RECT 457.690 400.000 457.970 400.110 ;
        RECT 456.020 386.340 456.620 386.480 ;
        RECT 456.020 53.710 456.160 386.340 ;
        RECT 455.960 53.390 456.220 53.710 ;
        RECT 851.560 53.390 851.820 53.710 ;
        RECT 851.620 1.770 851.760 53.390 ;
        RECT 853.710 1.770 854.270 2.400 ;
        RECT 851.620 1.630 854.270 1.770 ;
        RECT 853.710 -4.800 854.270 1.630 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.830 52.940 463.150 53.000 ;
        RECT 871.310 52.940 871.630 53.000 ;
        RECT 462.830 52.800 871.630 52.940 ;
        RECT 462.830 52.740 463.150 52.800 ;
        RECT 871.310 52.740 871.630 52.800 ;
      LAYER via ;
        RECT 462.860 52.740 463.120 53.000 ;
        RECT 871.340 52.740 871.600 53.000 ;
      LAYER met2 ;
        RECT 462.750 400.180 463.030 404.000 ;
        RECT 462.750 400.000 463.060 400.180 ;
        RECT 462.920 53.030 463.060 400.000 ;
        RECT 462.860 52.710 463.120 53.030 ;
        RECT 871.340 52.710 871.600 53.030 ;
        RECT 871.400 2.400 871.540 52.710 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 386.480 463.610 386.540 ;
        RECT 466.970 386.480 467.290 386.540 ;
        RECT 463.290 386.340 467.290 386.480 ;
        RECT 463.290 386.280 463.610 386.340 ;
        RECT 466.970 386.280 467.290 386.340 ;
        RECT 463.290 52.600 463.610 52.660 ;
        RECT 889.250 52.600 889.570 52.660 ;
        RECT 463.290 52.460 889.570 52.600 ;
        RECT 463.290 52.400 463.610 52.460 ;
        RECT 889.250 52.400 889.570 52.460 ;
      LAYER via ;
        RECT 463.320 386.280 463.580 386.540 ;
        RECT 467.000 386.280 467.260 386.540 ;
        RECT 463.320 52.400 463.580 52.660 ;
        RECT 889.280 52.400 889.540 52.660 ;
      LAYER met2 ;
        RECT 468.270 400.250 468.550 404.000 ;
        RECT 467.060 400.110 468.550 400.250 ;
        RECT 467.060 386.570 467.200 400.110 ;
        RECT 468.270 400.000 468.550 400.110 ;
        RECT 463.320 386.250 463.580 386.570 ;
        RECT 467.000 386.250 467.260 386.570 ;
        RECT 463.380 52.690 463.520 386.250 ;
        RECT 463.320 52.370 463.580 52.690 ;
        RECT 889.280 52.370 889.540 52.690 ;
        RECT 889.340 2.400 889.480 52.370 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 470.190 386.480 470.510 386.540 ;
        RECT 472.490 386.480 472.810 386.540 ;
        RECT 470.190 386.340 472.810 386.480 ;
        RECT 470.190 386.280 470.510 386.340 ;
        RECT 472.490 386.280 472.810 386.340 ;
        RECT 470.190 51.580 470.510 51.640 ;
        RECT 904.890 51.580 905.210 51.640 ;
        RECT 470.190 51.440 905.210 51.580 ;
        RECT 470.190 51.380 470.510 51.440 ;
        RECT 904.890 51.380 905.210 51.440 ;
      LAYER via ;
        RECT 470.220 386.280 470.480 386.540 ;
        RECT 472.520 386.280 472.780 386.540 ;
        RECT 470.220 51.380 470.480 51.640 ;
        RECT 904.920 51.380 905.180 51.640 ;
      LAYER met2 ;
        RECT 473.790 400.250 474.070 404.000 ;
        RECT 472.580 400.110 474.070 400.250 ;
        RECT 472.580 386.570 472.720 400.110 ;
        RECT 473.790 400.000 474.070 400.110 ;
        RECT 470.220 386.250 470.480 386.570 ;
        RECT 472.520 386.250 472.780 386.570 ;
        RECT 470.280 51.670 470.420 386.250 ;
        RECT 470.220 51.350 470.480 51.670 ;
        RECT 904.920 51.350 905.180 51.670 ;
        RECT 904.980 1.770 905.120 51.350 ;
        RECT 907.070 1.770 907.630 2.400 ;
        RECT 904.980 1.630 907.630 1.770 ;
        RECT 907.070 -4.800 907.630 1.630 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 478.930 389.880 479.250 389.940 ;
        RECT 755.390 389.880 755.710 389.940 ;
        RECT 478.930 389.740 755.710 389.880 ;
        RECT 478.930 389.680 479.250 389.740 ;
        RECT 755.390 389.680 755.710 389.740 ;
        RECT 755.390 26.760 755.710 26.820 ;
        RECT 924.670 26.760 924.990 26.820 ;
        RECT 755.390 26.620 924.990 26.760 ;
        RECT 755.390 26.560 755.710 26.620 ;
        RECT 924.670 26.560 924.990 26.620 ;
      LAYER via ;
        RECT 478.960 389.680 479.220 389.940 ;
        RECT 755.420 389.680 755.680 389.940 ;
        RECT 755.420 26.560 755.680 26.820 ;
        RECT 924.700 26.560 924.960 26.820 ;
      LAYER met2 ;
        RECT 478.850 400.180 479.130 404.000 ;
        RECT 478.850 400.000 479.160 400.180 ;
        RECT 479.020 389.970 479.160 400.000 ;
        RECT 478.960 389.650 479.220 389.970 ;
        RECT 755.420 389.650 755.680 389.970 ;
        RECT 755.480 26.850 755.620 389.650 ;
        RECT 755.420 26.530 755.680 26.850 ;
        RECT 924.700 26.530 924.960 26.850 ;
        RECT 924.760 2.400 924.900 26.530 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 49.540 483.850 49.600 ;
        RECT 942.610 49.540 942.930 49.600 ;
        RECT 483.530 49.400 942.930 49.540 ;
        RECT 483.530 49.340 483.850 49.400 ;
        RECT 942.610 49.340 942.930 49.400 ;
      LAYER via ;
        RECT 483.560 49.340 483.820 49.600 ;
        RECT 942.640 49.340 942.900 49.600 ;
      LAYER met2 ;
        RECT 484.370 400.250 484.650 404.000 ;
        RECT 483.620 400.110 484.650 400.250 ;
        RECT 483.620 49.630 483.760 400.110 ;
        RECT 484.370 400.000 484.650 400.110 ;
        RECT 483.560 49.310 483.820 49.630 ;
        RECT 942.640 49.310 942.900 49.630 ;
        RECT 942.700 2.400 942.840 49.310 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.890 60.420 491.210 60.480 ;
        RECT 960.090 60.420 960.410 60.480 ;
        RECT 490.890 60.280 960.410 60.420 ;
        RECT 490.890 60.220 491.210 60.280 ;
        RECT 960.090 60.220 960.410 60.280 ;
      LAYER via ;
        RECT 490.920 60.220 491.180 60.480 ;
        RECT 960.120 60.220 960.380 60.480 ;
      LAYER met2 ;
        RECT 489.890 400.250 490.170 404.000 ;
        RECT 489.890 400.110 491.120 400.250 ;
        RECT 489.890 400.000 490.170 400.110 ;
        RECT 490.980 60.510 491.120 400.110 ;
        RECT 490.920 60.190 491.180 60.510 ;
        RECT 960.120 60.190 960.380 60.510 ;
        RECT 960.180 2.400 960.320 60.190 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 386.140 490.750 386.200 ;
        RECT 493.650 386.140 493.970 386.200 ;
        RECT 490.430 386.000 493.970 386.140 ;
        RECT 490.430 385.940 490.750 386.000 ;
        RECT 493.650 385.940 493.970 386.000 ;
        RECT 490.430 60.080 490.750 60.140 ;
        RECT 975.730 60.080 976.050 60.140 ;
        RECT 490.430 59.940 976.050 60.080 ;
        RECT 490.430 59.880 490.750 59.940 ;
        RECT 975.730 59.880 976.050 59.940 ;
      LAYER via ;
        RECT 490.460 385.940 490.720 386.200 ;
        RECT 493.680 385.940 493.940 386.200 ;
        RECT 490.460 59.880 490.720 60.140 ;
        RECT 975.760 59.880 976.020 60.140 ;
      LAYER met2 ;
        RECT 494.950 400.250 495.230 404.000 ;
        RECT 493.740 400.110 495.230 400.250 ;
        RECT 493.740 386.230 493.880 400.110 ;
        RECT 494.950 400.000 495.230 400.110 ;
        RECT 490.460 385.910 490.720 386.230 ;
        RECT 493.680 385.910 493.940 386.230 ;
        RECT 490.520 60.170 490.660 385.910 ;
        RECT 490.460 59.850 490.720 60.170 ;
        RECT 975.760 59.850 976.020 60.170 ;
        RECT 975.820 1.770 975.960 59.850 ;
        RECT 977.910 1.770 978.470 2.400 ;
        RECT 975.820 1.630 978.470 1.770 ;
        RECT 977.910 -4.800 978.470 1.630 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.830 376.280 394.150 376.340 ;
        RECT 397.510 376.280 397.830 376.340 ;
        RECT 393.830 376.140 397.830 376.280 ;
        RECT 393.830 376.080 394.150 376.140 ;
        RECT 397.510 376.080 397.830 376.140 ;
        RECT 393.830 38.660 394.150 38.720 ;
        RECT 658.330 38.660 658.650 38.720 ;
        RECT 393.830 38.520 658.650 38.660 ;
        RECT 393.830 38.460 394.150 38.520 ;
        RECT 658.330 38.460 658.650 38.520 ;
      LAYER via ;
        RECT 393.860 376.080 394.120 376.340 ;
        RECT 397.540 376.080 397.800 376.340 ;
        RECT 393.860 38.460 394.120 38.720 ;
        RECT 658.360 38.460 658.620 38.720 ;
      LAYER met2 ;
        RECT 398.810 400.250 399.090 404.000 ;
        RECT 397.600 400.110 399.090 400.250 ;
        RECT 397.600 376.370 397.740 400.110 ;
        RECT 398.810 400.000 399.090 400.110 ;
        RECT 393.860 376.050 394.120 376.370 ;
        RECT 397.540 376.050 397.800 376.370 ;
        RECT 393.920 38.750 394.060 376.050 ;
        RECT 393.860 38.430 394.120 38.750 ;
        RECT 658.360 38.430 658.620 38.750 ;
        RECT 658.420 17.410 658.560 38.430 ;
        RECT 658.420 17.270 659.020 17.410 ;
        RECT 658.880 2.400 659.020 17.270 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.250 59.400 498.570 59.460 ;
        RECT 994.590 59.400 994.910 59.460 ;
        RECT 498.250 59.260 994.910 59.400 ;
        RECT 498.250 59.200 498.570 59.260 ;
        RECT 994.590 59.200 994.910 59.260 ;
      LAYER via ;
        RECT 498.280 59.200 498.540 59.460 ;
        RECT 994.620 59.200 994.880 59.460 ;
      LAYER met2 ;
        RECT 500.470 400.250 500.750 404.000 ;
        RECT 499.260 400.110 500.750 400.250 ;
        RECT 499.260 324.370 499.400 400.110 ;
        RECT 500.470 400.000 500.750 400.110 ;
        RECT 498.340 324.230 499.400 324.370 ;
        RECT 498.340 59.490 498.480 324.230 ;
        RECT 498.280 59.170 498.540 59.490 ;
        RECT 994.620 59.170 994.880 59.490 ;
        RECT 994.680 1.770 994.820 59.170 ;
        RECT 995.390 1.770 995.950 2.400 ;
        RECT 994.680 1.630 995.950 1.770 ;
        RECT 995.390 -4.800 995.950 1.630 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 59.060 504.550 59.120 ;
        RECT 1013.450 59.060 1013.770 59.120 ;
        RECT 504.230 58.920 1013.770 59.060 ;
        RECT 504.230 58.860 504.550 58.920 ;
        RECT 1013.450 58.860 1013.770 58.920 ;
      LAYER via ;
        RECT 504.260 58.860 504.520 59.120 ;
        RECT 1013.480 58.860 1013.740 59.120 ;
      LAYER met2 ;
        RECT 505.530 400.250 505.810 404.000 ;
        RECT 504.780 400.110 505.810 400.250 ;
        RECT 504.780 324.370 504.920 400.110 ;
        RECT 505.530 400.000 505.810 400.110 ;
        RECT 504.320 324.230 504.920 324.370 ;
        RECT 504.320 59.150 504.460 324.230 ;
        RECT 504.260 58.830 504.520 59.150 ;
        RECT 1013.480 58.830 1013.740 59.150 ;
        RECT 1013.540 2.400 1013.680 58.830 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 512.050 58.720 512.370 58.780 ;
        RECT 1030.930 58.720 1031.250 58.780 ;
        RECT 512.050 58.580 1031.250 58.720 ;
        RECT 512.050 58.520 512.370 58.580 ;
        RECT 1030.930 58.520 1031.250 58.580 ;
      LAYER via ;
        RECT 512.080 58.520 512.340 58.780 ;
        RECT 1030.960 58.520 1031.220 58.780 ;
      LAYER met2 ;
        RECT 511.050 400.250 511.330 404.000 ;
        RECT 511.050 400.110 512.280 400.250 ;
        RECT 511.050 400.000 511.330 400.110 ;
        RECT 512.140 58.810 512.280 400.110 ;
        RECT 512.080 58.490 512.340 58.810 ;
        RECT 1030.960 58.490 1031.220 58.810 ;
        RECT 1031.020 2.400 1031.160 58.490 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 386.480 511.910 386.540 ;
        RECT 515.270 386.480 515.590 386.540 ;
        RECT 511.590 386.340 515.590 386.480 ;
        RECT 511.590 386.280 511.910 386.340 ;
        RECT 515.270 386.280 515.590 386.340 ;
        RECT 511.590 56.340 511.910 56.400 ;
        RECT 1048.870 56.340 1049.190 56.400 ;
        RECT 511.590 56.200 1049.190 56.340 ;
        RECT 511.590 56.140 511.910 56.200 ;
        RECT 1048.870 56.140 1049.190 56.200 ;
      LAYER via ;
        RECT 511.620 386.280 511.880 386.540 ;
        RECT 515.300 386.280 515.560 386.540 ;
        RECT 511.620 56.140 511.880 56.400 ;
        RECT 1048.900 56.140 1049.160 56.400 ;
      LAYER met2 ;
        RECT 516.570 400.250 516.850 404.000 ;
        RECT 515.360 400.110 516.850 400.250 ;
        RECT 515.360 386.570 515.500 400.110 ;
        RECT 516.570 400.000 516.850 400.110 ;
        RECT 511.620 386.250 511.880 386.570 ;
        RECT 515.300 386.250 515.560 386.570 ;
        RECT 511.680 56.430 511.820 386.250 ;
        RECT 511.620 56.110 511.880 56.430 ;
        RECT 1048.900 56.110 1049.160 56.430 ;
        RECT 1048.960 2.400 1049.100 56.110 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 56.680 518.350 56.740 ;
        RECT 1066.810 56.680 1067.130 56.740 ;
        RECT 518.030 56.540 1067.130 56.680 ;
        RECT 518.030 56.480 518.350 56.540 ;
        RECT 1066.810 56.480 1067.130 56.540 ;
      LAYER via ;
        RECT 518.060 56.480 518.320 56.740 ;
        RECT 1066.840 56.480 1067.100 56.740 ;
      LAYER met2 ;
        RECT 521.630 400.250 521.910 404.000 ;
        RECT 520.880 400.110 521.910 400.250 ;
        RECT 520.880 386.480 521.020 400.110 ;
        RECT 521.630 400.000 521.910 400.110 ;
        RECT 518.120 386.340 521.020 386.480 ;
        RECT 518.120 56.770 518.260 386.340 ;
        RECT 518.060 56.450 518.320 56.770 ;
        RECT 1066.840 56.450 1067.100 56.770 ;
        RECT 1066.900 2.400 1067.040 56.450 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 77.760 525.250 77.820 ;
        RECT 1084.290 77.760 1084.610 77.820 ;
        RECT 524.930 77.620 1084.610 77.760 ;
        RECT 524.930 77.560 525.250 77.620 ;
        RECT 1084.290 77.560 1084.610 77.620 ;
      LAYER via ;
        RECT 524.960 77.560 525.220 77.820 ;
        RECT 1084.320 77.560 1084.580 77.820 ;
      LAYER met2 ;
        RECT 527.150 400.250 527.430 404.000 ;
        RECT 525.940 400.110 527.430 400.250 ;
        RECT 525.940 386.470 526.080 400.110 ;
        RECT 527.150 400.000 527.430 400.110 ;
        RECT 525.020 386.330 526.080 386.470 ;
        RECT 525.020 77.850 525.160 386.330 ;
        RECT 524.960 77.530 525.220 77.850 ;
        RECT 1084.320 77.530 1084.580 77.850 ;
        RECT 1084.380 2.400 1084.520 77.530 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 84.560 531.690 84.620 ;
        RECT 1097.170 84.560 1097.490 84.620 ;
        RECT 531.370 84.420 1097.490 84.560 ;
        RECT 531.370 84.360 531.690 84.420 ;
        RECT 1097.170 84.360 1097.490 84.420 ;
      LAYER via ;
        RECT 531.400 84.360 531.660 84.620 ;
        RECT 1097.200 84.360 1097.460 84.620 ;
      LAYER met2 ;
        RECT 532.670 400.250 532.950 404.000 ;
        RECT 531.460 400.110 532.950 400.250 ;
        RECT 531.460 84.650 531.600 400.110 ;
        RECT 532.670 400.000 532.950 400.110 ;
        RECT 531.400 84.330 531.660 84.650 ;
        RECT 1097.200 84.330 1097.460 84.650 ;
        RECT 1097.260 82.870 1097.400 84.330 ;
        RECT 1097.260 82.730 1100.160 82.870 ;
        RECT 1100.020 1.770 1100.160 82.730 ;
        RECT 1102.110 1.770 1102.670 2.400 ;
        RECT 1100.020 1.630 1102.670 1.770 ;
        RECT 1102.110 -4.800 1102.670 1.630 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 386.480 532.150 386.540 ;
        RECT 536.430 386.480 536.750 386.540 ;
        RECT 531.830 386.340 536.750 386.480 ;
        RECT 531.830 386.280 532.150 386.340 ;
        RECT 536.430 386.280 536.750 386.340 ;
        RECT 531.830 91.360 532.150 91.420 ;
        RECT 1117.870 91.360 1118.190 91.420 ;
        RECT 531.830 91.220 1118.190 91.360 ;
        RECT 531.830 91.160 532.150 91.220 ;
        RECT 1117.870 91.160 1118.190 91.220 ;
      LAYER via ;
        RECT 531.860 386.280 532.120 386.540 ;
        RECT 536.460 386.280 536.720 386.540 ;
        RECT 531.860 91.160 532.120 91.420 ;
        RECT 1117.900 91.160 1118.160 91.420 ;
      LAYER met2 ;
        RECT 537.730 400.250 538.010 404.000 ;
        RECT 536.520 400.110 538.010 400.250 ;
        RECT 536.520 386.570 536.660 400.110 ;
        RECT 537.730 400.000 538.010 400.110 ;
        RECT 531.860 386.250 532.120 386.570 ;
        RECT 536.460 386.250 536.720 386.570 ;
        RECT 531.920 91.450 532.060 386.250 ;
        RECT 531.860 91.130 532.120 91.450 ;
        RECT 1117.900 91.130 1118.160 91.450 ;
        RECT 1117.960 1.770 1118.100 91.130 ;
        RECT 1119.590 1.770 1120.150 2.400 ;
        RECT 1117.960 1.630 1120.150 1.770 ;
        RECT 1119.590 -4.800 1120.150 1.630 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 386.480 539.050 386.540 ;
        RECT 541.950 386.480 542.270 386.540 ;
        RECT 538.730 386.340 542.270 386.480 ;
        RECT 538.730 386.280 539.050 386.340 ;
        RECT 541.950 386.280 542.270 386.340 ;
        RECT 538.730 91.700 539.050 91.760 ;
        RECT 1132.130 91.700 1132.450 91.760 ;
        RECT 538.730 91.560 1132.450 91.700 ;
        RECT 538.730 91.500 539.050 91.560 ;
        RECT 1132.130 91.500 1132.450 91.560 ;
      LAYER via ;
        RECT 538.760 386.280 539.020 386.540 ;
        RECT 541.980 386.280 542.240 386.540 ;
        RECT 538.760 91.500 539.020 91.760 ;
        RECT 1132.160 91.500 1132.420 91.760 ;
      LAYER met2 ;
        RECT 543.250 400.250 543.530 404.000 ;
        RECT 542.040 400.110 543.530 400.250 ;
        RECT 542.040 386.570 542.180 400.110 ;
        RECT 543.250 400.000 543.530 400.110 ;
        RECT 538.760 386.250 539.020 386.570 ;
        RECT 541.980 386.250 542.240 386.570 ;
        RECT 538.820 91.790 538.960 386.250 ;
        RECT 538.760 91.470 539.020 91.790 ;
        RECT 1132.160 91.470 1132.420 91.790 ;
        RECT 1132.220 82.870 1132.360 91.470 ;
        RECT 1132.220 82.730 1137.880 82.870 ;
        RECT 1137.740 2.400 1137.880 82.730 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.090 376.280 546.410 376.340 ;
        RECT 547.470 376.280 547.790 376.340 ;
        RECT 546.090 376.140 547.790 376.280 ;
        RECT 546.090 376.080 546.410 376.140 ;
        RECT 547.470 376.080 547.790 376.140 ;
        RECT 546.090 92.040 546.410 92.100 ;
        RECT 1152.370 92.040 1152.690 92.100 ;
        RECT 546.090 91.900 1152.690 92.040 ;
        RECT 546.090 91.840 546.410 91.900 ;
        RECT 1152.370 91.840 1152.690 91.900 ;
      LAYER via ;
        RECT 546.120 376.080 546.380 376.340 ;
        RECT 547.500 376.080 547.760 376.340 ;
        RECT 546.120 91.840 546.380 92.100 ;
        RECT 1152.400 91.840 1152.660 92.100 ;
      LAYER met2 ;
        RECT 548.770 400.250 549.050 404.000 ;
        RECT 547.560 400.110 549.050 400.250 ;
        RECT 547.560 376.370 547.700 400.110 ;
        RECT 548.770 400.000 549.050 400.110 ;
        RECT 546.120 376.050 546.380 376.370 ;
        RECT 547.500 376.050 547.760 376.370 ;
        RECT 546.180 92.130 546.320 376.050 ;
        RECT 546.120 91.810 546.380 92.130 ;
        RECT 1152.400 91.810 1152.660 92.130 ;
        RECT 1152.460 82.870 1152.600 91.810 ;
        RECT 1152.460 82.730 1155.360 82.870 ;
        RECT 1155.220 2.400 1155.360 82.730 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 401.190 374.240 401.510 374.300 ;
        RECT 402.570 374.240 402.890 374.300 ;
        RECT 401.190 374.100 402.890 374.240 ;
        RECT 401.190 374.040 401.510 374.100 ;
        RECT 402.570 374.040 402.890 374.100 ;
        RECT 401.190 32.540 401.510 32.600 ;
        RECT 558.970 32.540 559.290 32.600 ;
        RECT 401.190 32.400 559.290 32.540 ;
        RECT 401.190 32.340 401.510 32.400 ;
        RECT 558.970 32.340 559.290 32.400 ;
        RECT 558.970 15.880 559.290 15.940 ;
        RECT 676.270 15.880 676.590 15.940 ;
        RECT 558.970 15.740 676.590 15.880 ;
        RECT 558.970 15.680 559.290 15.740 ;
        RECT 676.270 15.680 676.590 15.740 ;
      LAYER via ;
        RECT 401.220 374.040 401.480 374.300 ;
        RECT 402.600 374.040 402.860 374.300 ;
        RECT 401.220 32.340 401.480 32.600 ;
        RECT 559.000 32.340 559.260 32.600 ;
        RECT 559.000 15.680 559.260 15.940 ;
        RECT 676.300 15.680 676.560 15.940 ;
      LAYER met2 ;
        RECT 403.870 400.250 404.150 404.000 ;
        RECT 402.660 400.110 404.150 400.250 ;
        RECT 402.660 374.330 402.800 400.110 ;
        RECT 403.870 400.000 404.150 400.110 ;
        RECT 401.220 374.010 401.480 374.330 ;
        RECT 402.600 374.010 402.860 374.330 ;
        RECT 401.280 32.630 401.420 374.010 ;
        RECT 401.220 32.310 401.480 32.630 ;
        RECT 559.000 32.310 559.260 32.630 ;
        RECT 559.060 15.970 559.200 32.310 ;
        RECT 559.000 15.650 559.260 15.970 ;
        RECT 676.300 15.650 676.560 15.970 ;
        RECT 676.360 2.400 676.500 15.650 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.990 399.880 553.310 400.140 ;
        RECT 553.080 399.120 553.220 399.880 ;
        RECT 552.990 398.860 553.310 399.120 ;
        RECT 552.990 92.380 553.310 92.440 ;
        RECT 1173.070 92.380 1173.390 92.440 ;
        RECT 552.990 92.240 1173.390 92.380 ;
        RECT 552.990 92.180 553.310 92.240 ;
        RECT 1173.070 92.180 1173.390 92.240 ;
      LAYER via ;
        RECT 553.020 399.880 553.280 400.140 ;
        RECT 553.020 398.860 553.280 399.120 ;
        RECT 553.020 92.180 553.280 92.440 ;
        RECT 1173.100 92.180 1173.360 92.440 ;
      LAYER met2 ;
        RECT 553.830 400.930 554.110 404.000 ;
        RECT 553.080 400.790 554.110 400.930 ;
        RECT 553.080 400.170 553.220 400.790 ;
        RECT 553.020 399.850 553.280 400.170 ;
        RECT 553.830 400.000 554.110 400.790 ;
        RECT 553.020 398.830 553.280 399.150 ;
        RECT 553.080 92.470 553.220 398.830 ;
        RECT 553.020 92.150 553.280 92.470 ;
        RECT 1173.100 92.150 1173.360 92.470 ;
        RECT 1173.160 2.400 1173.300 92.150 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.890 92.720 560.210 92.780 ;
        RECT 1186.870 92.720 1187.190 92.780 ;
        RECT 559.890 92.580 1187.190 92.720 ;
        RECT 559.890 92.520 560.210 92.580 ;
        RECT 1186.870 92.520 1187.190 92.580 ;
      LAYER via ;
        RECT 559.920 92.520 560.180 92.780 ;
        RECT 1186.900 92.520 1187.160 92.780 ;
      LAYER met2 ;
        RECT 559.350 400.250 559.630 404.000 ;
        RECT 559.060 400.110 559.630 400.250 ;
        RECT 559.060 398.890 559.200 400.110 ;
        RECT 559.350 400.000 559.630 400.110 ;
        RECT 559.060 398.750 559.660 398.890 ;
        RECT 559.520 377.810 559.660 398.750 ;
        RECT 559.520 377.670 560.120 377.810 ;
        RECT 559.980 92.810 560.120 377.670 ;
        RECT 559.920 92.490 560.180 92.810 ;
        RECT 1186.900 92.490 1187.160 92.810 ;
        RECT 1186.960 82.870 1187.100 92.490 ;
        RECT 1186.960 82.730 1188.480 82.870 ;
        RECT 1188.340 1.770 1188.480 82.730 ;
        RECT 1190.430 1.770 1190.990 2.400 ;
        RECT 1188.340 1.630 1190.990 1.770 ;
        RECT 1190.430 -4.800 1190.990 1.630 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.350 96.460 560.670 96.520 ;
        RECT 1207.570 96.460 1207.890 96.520 ;
        RECT 560.350 96.320 1207.890 96.460 ;
        RECT 560.350 96.260 560.670 96.320 ;
        RECT 1207.570 96.260 1207.890 96.320 ;
      LAYER via ;
        RECT 560.380 96.260 560.640 96.520 ;
        RECT 1207.600 96.260 1207.860 96.520 ;
      LAYER met2 ;
        RECT 564.870 400.250 565.150 404.000 ;
        RECT 563.660 400.110 565.150 400.250 ;
        RECT 563.660 324.370 563.800 400.110 ;
        RECT 564.870 400.000 565.150 400.110 ;
        RECT 560.440 324.230 563.800 324.370 ;
        RECT 560.440 96.550 560.580 324.230 ;
        RECT 560.380 96.230 560.640 96.550 ;
        RECT 1207.600 96.230 1207.860 96.550 ;
        RECT 1207.660 82.870 1207.800 96.230 ;
        RECT 1207.660 82.730 1208.720 82.870 ;
        RECT 1208.580 2.400 1208.720 82.730 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.250 96.120 567.570 96.180 ;
        RECT 1221.370 96.120 1221.690 96.180 ;
        RECT 567.250 95.980 1221.690 96.120 ;
        RECT 567.250 95.920 567.570 95.980 ;
        RECT 1221.370 95.920 1221.690 95.980 ;
      LAYER via ;
        RECT 567.280 95.920 567.540 96.180 ;
        RECT 1221.400 95.920 1221.660 96.180 ;
      LAYER met2 ;
        RECT 569.930 400.250 570.210 404.000 ;
        RECT 568.720 400.110 570.210 400.250 ;
        RECT 568.720 324.370 568.860 400.110 ;
        RECT 569.930 400.000 570.210 400.110 ;
        RECT 567.340 324.230 568.860 324.370 ;
        RECT 567.340 96.210 567.480 324.230 ;
        RECT 567.280 95.890 567.540 96.210 ;
        RECT 1221.400 95.890 1221.660 96.210 ;
        RECT 1221.460 82.870 1221.600 95.890 ;
        RECT 1221.460 82.730 1226.200 82.870 ;
        RECT 1226.060 2.400 1226.200 82.730 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 574.150 95.780 574.470 95.840 ;
        RECT 1242.070 95.780 1242.390 95.840 ;
        RECT 574.150 95.640 1242.390 95.780 ;
        RECT 574.150 95.580 574.470 95.640 ;
        RECT 1242.070 95.580 1242.390 95.640 ;
      LAYER via ;
        RECT 574.180 95.580 574.440 95.840 ;
        RECT 1242.100 95.580 1242.360 95.840 ;
      LAYER met2 ;
        RECT 575.450 400.250 575.730 404.000 ;
        RECT 574.240 400.110 575.730 400.250 ;
        RECT 574.240 95.870 574.380 400.110 ;
        RECT 575.450 400.000 575.730 400.110 ;
        RECT 574.180 95.550 574.440 95.870 ;
        RECT 1242.100 95.550 1242.360 95.870 ;
        RECT 1242.160 1.770 1242.300 95.550 ;
        RECT 1243.790 1.770 1244.350 2.400 ;
        RECT 1242.160 1.630 1244.350 1.770 ;
        RECT 1243.790 -4.800 1244.350 1.630 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 117.200 580.910 117.260 ;
        RECT 1255.870 117.200 1256.190 117.260 ;
        RECT 580.590 117.060 1256.190 117.200 ;
        RECT 580.590 117.000 580.910 117.060 ;
        RECT 1255.870 117.000 1256.190 117.060 ;
        RECT 1255.870 20.980 1256.190 21.040 ;
        RECT 1261.850 20.980 1262.170 21.040 ;
        RECT 1255.870 20.840 1262.170 20.980 ;
        RECT 1255.870 20.780 1256.190 20.840 ;
        RECT 1261.850 20.780 1262.170 20.840 ;
      LAYER via ;
        RECT 580.620 117.000 580.880 117.260 ;
        RECT 1255.900 117.000 1256.160 117.260 ;
        RECT 1255.900 20.780 1256.160 21.040 ;
        RECT 1261.880 20.780 1262.140 21.040 ;
      LAYER met2 ;
        RECT 580.970 400.250 581.250 404.000 ;
        RECT 580.680 400.110 581.250 400.250 ;
        RECT 580.680 117.290 580.820 400.110 ;
        RECT 580.970 400.000 581.250 400.110 ;
        RECT 580.620 116.970 580.880 117.290 ;
        RECT 1255.900 116.970 1256.160 117.290 ;
        RECT 1255.960 21.070 1256.100 116.970 ;
        RECT 1255.900 20.750 1256.160 21.070 ;
        RECT 1261.880 20.750 1262.140 21.070 ;
        RECT 1261.940 2.400 1262.080 20.750 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.050 118.900 581.370 118.960 ;
        RECT 1276.570 118.900 1276.890 118.960 ;
        RECT 581.050 118.760 1276.890 118.900 ;
        RECT 581.050 118.700 581.370 118.760 ;
        RECT 1276.570 118.700 1276.890 118.760 ;
      LAYER via ;
        RECT 581.080 118.700 581.340 118.960 ;
        RECT 1276.600 118.700 1276.860 118.960 ;
      LAYER met2 ;
        RECT 586.030 400.250 586.310 404.000 ;
        RECT 584.820 400.110 586.310 400.250 ;
        RECT 584.820 324.370 584.960 400.110 ;
        RECT 586.030 400.000 586.310 400.110 ;
        RECT 581.140 324.230 584.960 324.370 ;
        RECT 581.140 118.990 581.280 324.230 ;
        RECT 581.080 118.670 581.340 118.990 ;
        RECT 1276.600 118.670 1276.860 118.990 ;
        RECT 1276.660 82.870 1276.800 118.670 ;
        RECT 1276.660 82.730 1279.560 82.870 ;
        RECT 1279.420 2.400 1279.560 82.730 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.490 98.160 587.810 98.220 ;
        RECT 1297.270 98.160 1297.590 98.220 ;
        RECT 587.490 98.020 1297.590 98.160 ;
        RECT 587.490 97.960 587.810 98.020 ;
        RECT 1297.270 97.960 1297.590 98.020 ;
      LAYER via ;
        RECT 587.520 97.960 587.780 98.220 ;
        RECT 1297.300 97.960 1297.560 98.220 ;
      LAYER met2 ;
        RECT 591.550 400.250 591.830 404.000 ;
        RECT 590.340 400.110 591.830 400.250 ;
        RECT 590.340 351.970 590.480 400.110 ;
        RECT 591.550 400.000 591.830 400.110 ;
        RECT 587.580 351.830 590.480 351.970 ;
        RECT 587.580 98.250 587.720 351.830 ;
        RECT 587.520 97.930 587.780 98.250 ;
        RECT 1297.300 97.930 1297.560 98.250 ;
        RECT 1297.360 2.400 1297.500 97.930 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.850 98.500 595.170 98.560 ;
        RECT 1311.070 98.500 1311.390 98.560 ;
        RECT 594.850 98.360 1311.390 98.500 ;
        RECT 594.850 98.300 595.170 98.360 ;
        RECT 1311.070 98.300 1311.390 98.360 ;
      LAYER via ;
        RECT 594.880 98.300 595.140 98.560 ;
        RECT 1311.100 98.300 1311.360 98.560 ;
      LAYER met2 ;
        RECT 597.070 400.250 597.350 404.000 ;
        RECT 595.860 400.110 597.350 400.250 ;
        RECT 595.860 324.370 596.000 400.110 ;
        RECT 597.070 400.000 597.350 400.110 ;
        RECT 594.940 324.230 596.000 324.370 ;
        RECT 594.940 98.590 595.080 324.230 ;
        RECT 594.880 98.270 595.140 98.590 ;
        RECT 1311.100 98.270 1311.360 98.590 ;
        RECT 1311.160 82.870 1311.300 98.270 ;
        RECT 1311.160 82.730 1312.680 82.870 ;
        RECT 1312.540 1.770 1312.680 82.730 ;
        RECT 1314.630 1.770 1315.190 2.400 ;
        RECT 1312.540 1.630 1315.190 1.770 ;
        RECT 1314.630 -4.800 1315.190 1.630 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.290 98.840 601.610 98.900 ;
        RECT 1331.770 98.840 1332.090 98.900 ;
        RECT 601.290 98.700 1332.090 98.840 ;
        RECT 601.290 98.640 601.610 98.700 ;
        RECT 1331.770 98.640 1332.090 98.700 ;
      LAYER via ;
        RECT 601.320 98.640 601.580 98.900 ;
        RECT 1331.800 98.640 1332.060 98.900 ;
      LAYER met2 ;
        RECT 602.130 400.250 602.410 404.000 ;
        RECT 601.380 400.110 602.410 400.250 ;
        RECT 601.380 98.930 601.520 400.110 ;
        RECT 602.130 400.000 602.410 400.110 ;
        RECT 601.320 98.610 601.580 98.930 ;
        RECT 1331.800 98.610 1332.060 98.930 ;
        RECT 1331.860 82.870 1332.000 98.610 ;
        RECT 1331.860 82.730 1332.920 82.870 ;
        RECT 1332.780 2.400 1332.920 82.730 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.630 32.880 407.950 32.940 ;
        RECT 564.490 32.880 564.810 32.940 ;
        RECT 407.630 32.740 564.810 32.880 ;
        RECT 407.630 32.680 407.950 32.740 ;
        RECT 564.490 32.680 564.810 32.740 ;
        RECT 564.490 16.220 564.810 16.280 ;
        RECT 694.210 16.220 694.530 16.280 ;
        RECT 564.490 16.080 694.530 16.220 ;
        RECT 564.490 16.020 564.810 16.080 ;
        RECT 694.210 16.020 694.530 16.080 ;
      LAYER via ;
        RECT 407.660 32.680 407.920 32.940 ;
        RECT 564.520 32.680 564.780 32.940 ;
        RECT 564.520 16.020 564.780 16.280 ;
        RECT 694.240 16.020 694.500 16.280 ;
      LAYER met2 ;
        RECT 409.390 400.250 409.670 404.000 ;
        RECT 408.180 400.110 409.670 400.250 ;
        RECT 408.180 386.650 408.320 400.110 ;
        RECT 409.390 400.000 409.670 400.110 ;
        RECT 407.720 386.510 408.320 386.650 ;
        RECT 407.720 32.970 407.860 386.510 ;
        RECT 407.660 32.650 407.920 32.970 ;
        RECT 564.520 32.650 564.780 32.970 ;
        RECT 564.580 16.310 564.720 32.650 ;
        RECT 564.520 15.990 564.780 16.310 ;
        RECT 694.240 15.990 694.500 16.310 ;
        RECT 694.300 2.400 694.440 15.990 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 99.180 608.510 99.240 ;
        RECT 1345.570 99.180 1345.890 99.240 ;
        RECT 608.190 99.040 1345.890 99.180 ;
        RECT 608.190 98.980 608.510 99.040 ;
        RECT 1345.570 98.980 1345.890 99.040 ;
      LAYER via ;
        RECT 608.220 98.980 608.480 99.240 ;
        RECT 1345.600 98.980 1345.860 99.240 ;
      LAYER met2 ;
        RECT 607.650 400.250 607.930 404.000 ;
        RECT 607.650 400.110 608.420 400.250 ;
        RECT 607.650 400.000 607.930 400.110 ;
        RECT 608.280 99.270 608.420 400.110 ;
        RECT 608.220 98.950 608.480 99.270 ;
        RECT 1345.600 98.950 1345.860 99.270 ;
        RECT 1345.660 82.870 1345.800 98.950 ;
        RECT 1345.660 82.730 1350.400 82.870 ;
        RECT 1350.260 2.400 1350.400 82.730 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 375.940 608.050 376.000 ;
        RECT 611.870 375.940 612.190 376.000 ;
        RECT 607.730 375.800 612.190 375.940 ;
        RECT 607.730 375.740 608.050 375.800 ;
        RECT 611.870 375.740 612.190 375.800 ;
        RECT 607.730 99.520 608.050 99.580 ;
        RECT 1366.270 99.520 1366.590 99.580 ;
        RECT 607.730 99.380 1366.590 99.520 ;
        RECT 607.730 99.320 608.050 99.380 ;
        RECT 1366.270 99.320 1366.590 99.380 ;
      LAYER via ;
        RECT 607.760 375.740 608.020 376.000 ;
        RECT 611.900 375.740 612.160 376.000 ;
        RECT 607.760 99.320 608.020 99.580 ;
        RECT 1366.300 99.320 1366.560 99.580 ;
      LAYER met2 ;
        RECT 612.710 400.250 612.990 404.000 ;
        RECT 611.960 400.110 612.990 400.250 ;
        RECT 611.960 376.030 612.100 400.110 ;
        RECT 612.710 400.000 612.990 400.110 ;
        RECT 607.760 375.710 608.020 376.030 ;
        RECT 611.900 375.710 612.160 376.030 ;
        RECT 607.820 99.610 607.960 375.710 ;
        RECT 607.760 99.290 608.020 99.610 ;
        RECT 1366.300 99.290 1366.560 99.610 ;
        RECT 1366.360 1.770 1366.500 99.290 ;
        RECT 1367.990 1.770 1368.550 2.400 ;
        RECT 1366.360 1.630 1368.550 1.770 ;
        RECT 1367.990 -4.800 1368.550 1.630 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.630 375.940 614.950 376.000 ;
        RECT 616.930 375.940 617.250 376.000 ;
        RECT 614.630 375.800 617.250 375.940 ;
        RECT 614.630 375.740 614.950 375.800 ;
        RECT 616.930 375.740 617.250 375.800 ;
        RECT 614.630 103.260 614.950 103.320 ;
        RECT 1380.070 103.260 1380.390 103.320 ;
        RECT 614.630 103.120 1380.390 103.260 ;
        RECT 614.630 103.060 614.950 103.120 ;
        RECT 1380.070 103.060 1380.390 103.120 ;
        RECT 1380.070 20.980 1380.390 21.040 ;
        RECT 1383.750 20.980 1384.070 21.040 ;
        RECT 1380.070 20.840 1384.070 20.980 ;
        RECT 1380.070 20.780 1380.390 20.840 ;
        RECT 1383.750 20.780 1384.070 20.840 ;
      LAYER via ;
        RECT 614.660 375.740 614.920 376.000 ;
        RECT 616.960 375.740 617.220 376.000 ;
        RECT 614.660 103.060 614.920 103.320 ;
        RECT 1380.100 103.060 1380.360 103.320 ;
        RECT 1380.100 20.780 1380.360 21.040 ;
        RECT 1383.780 20.780 1384.040 21.040 ;
      LAYER met2 ;
        RECT 618.230 400.250 618.510 404.000 ;
        RECT 617.020 400.110 618.510 400.250 ;
        RECT 617.020 376.030 617.160 400.110 ;
        RECT 618.230 400.000 618.510 400.110 ;
        RECT 614.660 375.710 614.920 376.030 ;
        RECT 616.960 375.710 617.220 376.030 ;
        RECT 614.720 103.350 614.860 375.710 ;
        RECT 614.660 103.030 614.920 103.350 ;
        RECT 1380.100 103.030 1380.360 103.350 ;
        RECT 1380.160 21.070 1380.300 103.030 ;
        RECT 1380.100 20.750 1380.360 21.070 ;
        RECT 1383.780 20.750 1384.040 21.070 ;
        RECT 1383.840 1.770 1383.980 20.750 ;
        RECT 1385.470 1.770 1386.030 2.400 ;
        RECT 1383.840 1.630 1386.030 1.770 ;
        RECT 1385.470 -4.800 1386.030 1.630 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 102.920 622.310 102.980 ;
        RECT 1400.770 102.920 1401.090 102.980 ;
        RECT 621.990 102.780 1401.090 102.920 ;
        RECT 621.990 102.720 622.310 102.780 ;
        RECT 1400.770 102.720 1401.090 102.780 ;
      LAYER via ;
        RECT 622.020 102.720 622.280 102.980 ;
        RECT 1400.800 102.720 1401.060 102.980 ;
      LAYER met2 ;
        RECT 623.750 400.250 624.030 404.000 ;
        RECT 622.540 400.110 624.030 400.250 ;
        RECT 622.540 351.970 622.680 400.110 ;
        RECT 623.750 400.000 624.030 400.110 ;
        RECT 622.080 351.830 622.680 351.970 ;
        RECT 622.080 103.010 622.220 351.830 ;
        RECT 622.020 102.690 622.280 103.010 ;
        RECT 1400.800 102.690 1401.060 103.010 ;
        RECT 1400.860 82.870 1401.000 102.690 ;
        RECT 1400.860 82.730 1403.760 82.870 ;
        RECT 1403.620 2.400 1403.760 82.730 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.350 102.580 629.670 102.640 ;
        RECT 1421.470 102.580 1421.790 102.640 ;
        RECT 629.350 102.440 1421.790 102.580 ;
        RECT 629.350 102.380 629.670 102.440 ;
        RECT 1421.470 102.380 1421.790 102.440 ;
      LAYER via ;
        RECT 629.380 102.380 629.640 102.640 ;
        RECT 1421.500 102.380 1421.760 102.640 ;
      LAYER met2 ;
        RECT 628.810 400.250 629.090 404.000 ;
        RECT 628.810 400.110 629.580 400.250 ;
        RECT 628.810 400.000 629.090 400.110 ;
        RECT 629.440 102.670 629.580 400.110 ;
        RECT 629.380 102.350 629.640 102.670 ;
        RECT 1421.500 102.350 1421.760 102.670 ;
        RECT 1421.560 2.400 1421.700 102.350 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.890 376.620 629.210 376.680 ;
        RECT 633.030 376.620 633.350 376.680 ;
        RECT 628.890 376.480 633.350 376.620 ;
        RECT 628.890 376.420 629.210 376.480 ;
        RECT 633.030 376.420 633.350 376.480 ;
        RECT 628.890 102.240 629.210 102.300 ;
        RECT 1435.270 102.240 1435.590 102.300 ;
        RECT 628.890 102.100 1435.590 102.240 ;
        RECT 628.890 102.040 629.210 102.100 ;
        RECT 1435.270 102.040 1435.590 102.100 ;
      LAYER via ;
        RECT 628.920 376.420 629.180 376.680 ;
        RECT 633.060 376.420 633.320 376.680 ;
        RECT 628.920 102.040 629.180 102.300 ;
        RECT 1435.300 102.040 1435.560 102.300 ;
      LAYER met2 ;
        RECT 634.330 400.250 634.610 404.000 ;
        RECT 633.120 400.110 634.610 400.250 ;
        RECT 633.120 376.710 633.260 400.110 ;
        RECT 634.330 400.000 634.610 400.110 ;
        RECT 628.920 376.390 629.180 376.710 ;
        RECT 633.060 376.390 633.320 376.710 ;
        RECT 628.980 102.330 629.120 376.390 ;
        RECT 628.920 102.010 629.180 102.330 ;
        RECT 1435.300 102.010 1435.560 102.330 ;
        RECT 1435.360 82.870 1435.500 102.010 ;
        RECT 1435.360 82.730 1436.880 82.870 ;
        RECT 1436.740 1.770 1436.880 82.730 ;
        RECT 1438.830 1.770 1439.390 2.400 ;
        RECT 1436.740 1.630 1439.390 1.770 ;
        RECT 1438.830 -4.800 1439.390 1.630 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.790 101.900 636.110 101.960 ;
        RECT 1455.970 101.900 1456.290 101.960 ;
        RECT 635.790 101.760 1456.290 101.900 ;
        RECT 635.790 101.700 636.110 101.760 ;
        RECT 1455.970 101.700 1456.290 101.760 ;
      LAYER via ;
        RECT 635.820 101.700 636.080 101.960 ;
        RECT 1456.000 101.700 1456.260 101.960 ;
      LAYER met2 ;
        RECT 639.850 400.250 640.130 404.000 ;
        RECT 638.640 400.110 640.130 400.250 ;
        RECT 638.640 399.570 638.780 400.110 ;
        RECT 639.850 400.000 640.130 400.110 ;
        RECT 637.720 399.430 638.780 399.570 ;
        RECT 637.720 351.970 637.860 399.430 ;
        RECT 635.880 351.830 637.860 351.970 ;
        RECT 635.880 101.990 636.020 351.830 ;
        RECT 635.820 101.670 636.080 101.990 ;
        RECT 1456.000 101.670 1456.260 101.990 ;
        RECT 1456.060 82.870 1456.200 101.670 ;
        RECT 1456.060 82.730 1457.120 82.870 ;
        RECT 1456.980 2.400 1457.120 82.730 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 643.150 101.560 643.470 101.620 ;
        RECT 1469.770 101.560 1470.090 101.620 ;
        RECT 643.150 101.420 1470.090 101.560 ;
        RECT 643.150 101.360 643.470 101.420 ;
        RECT 1469.770 101.360 1470.090 101.420 ;
      LAYER via ;
        RECT 643.180 101.360 643.440 101.620 ;
        RECT 1469.800 101.360 1470.060 101.620 ;
      LAYER met2 ;
        RECT 644.910 400.250 645.190 404.000 ;
        RECT 643.700 400.110 645.190 400.250 ;
        RECT 643.700 324.370 643.840 400.110 ;
        RECT 644.910 400.000 645.190 400.110 ;
        RECT 643.240 324.230 643.840 324.370 ;
        RECT 643.240 101.650 643.380 324.230 ;
        RECT 643.180 101.330 643.440 101.650 ;
        RECT 1469.800 101.330 1470.060 101.650 ;
        RECT 1469.860 82.870 1470.000 101.330 ;
        RECT 1469.860 82.730 1474.600 82.870 ;
        RECT 1474.460 2.400 1474.600 82.730 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.130 101.220 649.450 101.280 ;
        RECT 1490.470 101.220 1490.790 101.280 ;
        RECT 649.130 101.080 1490.790 101.220 ;
        RECT 649.130 101.020 649.450 101.080 ;
        RECT 1490.470 101.020 1490.790 101.080 ;
      LAYER via ;
        RECT 649.160 101.020 649.420 101.280 ;
        RECT 1490.500 101.020 1490.760 101.280 ;
      LAYER met2 ;
        RECT 650.430 400.250 650.710 404.000 ;
        RECT 649.220 400.110 650.710 400.250 ;
        RECT 649.220 101.310 649.360 400.110 ;
        RECT 650.430 400.000 650.710 400.110 ;
        RECT 649.160 100.990 649.420 101.310 ;
        RECT 1490.500 100.990 1490.760 101.310 ;
        RECT 1490.560 1.770 1490.700 100.990 ;
        RECT 1492.190 1.770 1492.750 2.400 ;
        RECT 1490.560 1.630 1492.750 1.770 ;
        RECT 1492.190 -4.800 1492.750 1.630 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.490 100.880 656.810 100.940 ;
        RECT 1504.270 100.880 1504.590 100.940 ;
        RECT 656.490 100.740 1504.590 100.880 ;
        RECT 656.490 100.680 656.810 100.740 ;
        RECT 1504.270 100.680 1504.590 100.740 ;
      LAYER via ;
        RECT 656.520 100.680 656.780 100.940 ;
        RECT 1504.300 100.680 1504.560 100.940 ;
      LAYER met2 ;
        RECT 655.950 400.180 656.230 404.000 ;
        RECT 655.950 400.000 656.260 400.180 ;
        RECT 656.120 396.850 656.260 400.000 ;
        RECT 656.120 396.710 656.720 396.850 ;
        RECT 656.580 100.970 656.720 396.710 ;
        RECT 656.520 100.650 656.780 100.970 ;
        RECT 1504.300 100.650 1504.560 100.970 ;
        RECT 1504.360 82.870 1504.500 100.650 ;
        RECT 1504.360 82.730 1507.720 82.870 ;
        RECT 1507.580 1.770 1507.720 82.730 ;
        RECT 1509.670 1.770 1510.230 2.400 ;
        RECT 1507.580 1.630 1510.230 1.770 ;
        RECT 1509.670 -4.800 1510.230 1.630 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.530 33.560 414.850 33.620 ;
        RECT 552.990 33.560 553.310 33.620 ;
        RECT 414.530 33.420 553.310 33.560 ;
        RECT 414.530 33.360 414.850 33.420 ;
        RECT 552.990 33.360 553.310 33.420 ;
        RECT 552.990 16.560 553.310 16.620 ;
        RECT 712.150 16.560 712.470 16.620 ;
        RECT 552.990 16.420 712.470 16.560 ;
        RECT 552.990 16.360 553.310 16.420 ;
        RECT 712.150 16.360 712.470 16.420 ;
      LAYER via ;
        RECT 414.560 33.360 414.820 33.620 ;
        RECT 553.020 33.360 553.280 33.620 ;
        RECT 553.020 16.360 553.280 16.620 ;
        RECT 712.180 16.360 712.440 16.620 ;
      LAYER met2 ;
        RECT 414.450 400.180 414.730 404.000 ;
        RECT 414.450 400.000 414.760 400.180 ;
        RECT 414.620 33.650 414.760 400.000 ;
        RECT 414.560 33.330 414.820 33.650 ;
        RECT 553.020 33.330 553.280 33.650 ;
        RECT 553.080 16.650 553.220 33.330 ;
        RECT 553.020 16.330 553.280 16.650 ;
        RECT 712.180 16.330 712.440 16.650 ;
        RECT 712.240 2.400 712.380 16.330 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.030 396.340 656.350 396.400 ;
        RECT 659.710 396.340 660.030 396.400 ;
        RECT 656.030 396.200 660.030 396.340 ;
        RECT 656.030 396.140 656.350 396.200 ;
        RECT 659.710 396.140 660.030 396.200 ;
        RECT 656.030 100.540 656.350 100.600 ;
        RECT 1524.970 100.540 1525.290 100.600 ;
        RECT 656.030 100.400 1525.290 100.540 ;
        RECT 656.030 100.340 656.350 100.400 ;
        RECT 1524.970 100.340 1525.290 100.400 ;
      LAYER via ;
        RECT 656.060 396.140 656.320 396.400 ;
        RECT 659.740 396.140 660.000 396.400 ;
        RECT 656.060 100.340 656.320 100.600 ;
        RECT 1525.000 100.340 1525.260 100.600 ;
      LAYER met2 ;
        RECT 661.010 400.250 661.290 404.000 ;
        RECT 659.800 400.110 661.290 400.250 ;
        RECT 659.800 396.430 659.940 400.110 ;
        RECT 661.010 400.000 661.290 400.110 ;
        RECT 656.060 396.110 656.320 396.430 ;
        RECT 659.740 396.110 660.000 396.430 ;
        RECT 656.120 100.630 656.260 396.110 ;
        RECT 656.060 100.310 656.320 100.630 ;
        RECT 1525.000 100.310 1525.260 100.630 ;
        RECT 1525.060 82.870 1525.200 100.310 ;
        RECT 1525.060 82.730 1527.960 82.870 ;
        RECT 1527.820 2.400 1527.960 82.730 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 375.940 663.710 376.000 ;
        RECT 665.230 375.940 665.550 376.000 ;
        RECT 663.390 375.800 665.550 375.940 ;
        RECT 663.390 375.740 663.710 375.800 ;
        RECT 665.230 375.740 665.550 375.800 ;
        RECT 663.390 100.200 663.710 100.260 ;
        RECT 1539.230 100.200 1539.550 100.260 ;
        RECT 663.390 100.060 1539.550 100.200 ;
        RECT 663.390 100.000 663.710 100.060 ;
        RECT 1539.230 100.000 1539.550 100.060 ;
        RECT 1539.230 20.980 1539.550 21.040 ;
        RECT 1545.210 20.980 1545.530 21.040 ;
        RECT 1539.230 20.840 1545.530 20.980 ;
        RECT 1539.230 20.780 1539.550 20.840 ;
        RECT 1545.210 20.780 1545.530 20.840 ;
      LAYER via ;
        RECT 663.420 375.740 663.680 376.000 ;
        RECT 665.260 375.740 665.520 376.000 ;
        RECT 663.420 100.000 663.680 100.260 ;
        RECT 1539.260 100.000 1539.520 100.260 ;
        RECT 1539.260 20.780 1539.520 21.040 ;
        RECT 1545.240 20.780 1545.500 21.040 ;
      LAYER met2 ;
        RECT 666.530 400.250 666.810 404.000 ;
        RECT 665.320 400.110 666.810 400.250 ;
        RECT 665.320 376.030 665.460 400.110 ;
        RECT 666.530 400.000 666.810 400.110 ;
        RECT 663.420 375.710 663.680 376.030 ;
        RECT 665.260 375.710 665.520 376.030 ;
        RECT 663.480 100.290 663.620 375.710 ;
        RECT 663.420 99.970 663.680 100.290 ;
        RECT 1539.260 99.970 1539.520 100.290 ;
        RECT 1539.320 21.070 1539.460 99.970 ;
        RECT 1539.260 20.750 1539.520 21.070 ;
        RECT 1545.240 20.750 1545.500 21.070 ;
        RECT 1545.300 2.400 1545.440 20.750 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.290 376.280 670.610 376.340 ;
        RECT 671.210 376.280 671.530 376.340 ;
        RECT 670.290 376.140 671.530 376.280 ;
        RECT 670.290 376.080 670.610 376.140 ;
        RECT 671.210 376.080 671.530 376.140 ;
        RECT 670.290 99.860 670.610 99.920 ;
        RECT 1559.470 99.860 1559.790 99.920 ;
        RECT 670.290 99.720 1559.790 99.860 ;
        RECT 670.290 99.660 670.610 99.720 ;
        RECT 1559.470 99.660 1559.790 99.720 ;
      LAYER via ;
        RECT 670.320 376.080 670.580 376.340 ;
        RECT 671.240 376.080 671.500 376.340 ;
        RECT 670.320 99.660 670.580 99.920 ;
        RECT 1559.500 99.660 1559.760 99.920 ;
      LAYER met2 ;
        RECT 672.050 400.250 672.330 404.000 ;
        RECT 671.300 400.110 672.330 400.250 ;
        RECT 671.300 376.370 671.440 400.110 ;
        RECT 672.050 400.000 672.330 400.110 ;
        RECT 670.320 376.050 670.580 376.370 ;
        RECT 671.240 376.050 671.500 376.370 ;
        RECT 670.380 99.950 670.520 376.050 ;
        RECT 670.320 99.630 670.580 99.950 ;
        RECT 1559.500 99.630 1559.760 99.950 ;
        RECT 1559.560 82.870 1559.700 99.630 ;
        RECT 1559.560 82.730 1561.080 82.870 ;
        RECT 1560.940 1.770 1561.080 82.730 ;
        RECT 1563.030 1.770 1563.590 2.400 ;
        RECT 1560.940 1.630 1563.590 1.770 ;
        RECT 1563.030 -4.800 1563.590 1.630 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 677.190 126.040 677.510 126.100 ;
        RECT 1580.170 126.040 1580.490 126.100 ;
        RECT 677.190 125.900 1580.490 126.040 ;
        RECT 677.190 125.840 677.510 125.900 ;
        RECT 1580.170 125.840 1580.490 125.900 ;
      LAYER via ;
        RECT 677.220 125.840 677.480 126.100 ;
        RECT 1580.200 125.840 1580.460 126.100 ;
      LAYER met2 ;
        RECT 677.110 400.180 677.390 404.000 ;
        RECT 677.110 400.000 677.420 400.180 ;
        RECT 677.280 126.130 677.420 400.000 ;
        RECT 677.220 125.810 677.480 126.130 ;
        RECT 1580.200 125.810 1580.460 126.130 ;
        RECT 1580.260 82.870 1580.400 125.810 ;
        RECT 1580.260 82.730 1581.320 82.870 ;
        RECT 1581.180 2.400 1581.320 82.730 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 677.650 126.380 677.970 126.440 ;
        RECT 1593.970 126.380 1594.290 126.440 ;
        RECT 677.650 126.240 1594.290 126.380 ;
        RECT 677.650 126.180 677.970 126.240 ;
        RECT 1593.970 126.180 1594.290 126.240 ;
      LAYER via ;
        RECT 677.680 126.180 677.940 126.440 ;
        RECT 1594.000 126.180 1594.260 126.440 ;
      LAYER met2 ;
        RECT 682.630 400.250 682.910 404.000 ;
        RECT 681.420 400.110 682.910 400.250 ;
        RECT 681.420 324.370 681.560 400.110 ;
        RECT 682.630 400.000 682.910 400.110 ;
        RECT 677.740 324.230 681.560 324.370 ;
        RECT 677.740 126.470 677.880 324.230 ;
        RECT 677.680 126.150 677.940 126.470 ;
        RECT 1594.000 126.150 1594.260 126.470 ;
        RECT 1594.060 82.870 1594.200 126.150 ;
        RECT 1594.060 82.730 1598.800 82.870 ;
        RECT 1598.660 2.400 1598.800 82.730 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.550 126.720 684.870 126.780 ;
        RECT 1614.670 126.720 1614.990 126.780 ;
        RECT 684.550 126.580 1614.990 126.720 ;
        RECT 684.550 126.520 684.870 126.580 ;
        RECT 1614.670 126.520 1614.990 126.580 ;
      LAYER via ;
        RECT 684.580 126.520 684.840 126.780 ;
        RECT 1614.700 126.520 1614.960 126.780 ;
      LAYER met2 ;
        RECT 688.150 400.250 688.430 404.000 ;
        RECT 686.940 400.110 688.430 400.250 ;
        RECT 686.940 324.370 687.080 400.110 ;
        RECT 688.150 400.000 688.430 400.110 ;
        RECT 684.640 324.230 687.080 324.370 ;
        RECT 684.640 126.810 684.780 324.230 ;
        RECT 684.580 126.490 684.840 126.810 ;
        RECT 1614.700 126.490 1614.960 126.810 ;
        RECT 1614.760 1.770 1614.900 126.490 ;
        RECT 1616.390 1.770 1616.950 2.400 ;
        RECT 1614.760 1.630 1616.950 1.770 ;
        RECT 1616.390 -4.800 1616.950 1.630 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.990 127.060 691.310 127.120 ;
        RECT 1628.470 127.060 1628.790 127.120 ;
        RECT 690.990 126.920 1628.790 127.060 ;
        RECT 690.990 126.860 691.310 126.920 ;
        RECT 1628.470 126.860 1628.790 126.920 ;
      LAYER via ;
        RECT 691.020 126.860 691.280 127.120 ;
        RECT 1628.500 126.860 1628.760 127.120 ;
      LAYER met2 ;
        RECT 693.210 400.250 693.490 404.000 ;
        RECT 692.000 400.110 693.490 400.250 ;
        RECT 692.000 324.370 692.140 400.110 ;
        RECT 693.210 400.000 693.490 400.110 ;
        RECT 691.080 324.230 692.140 324.370 ;
        RECT 691.080 127.150 691.220 324.230 ;
        RECT 691.020 126.830 691.280 127.150 ;
        RECT 1628.500 126.830 1628.760 127.150 ;
        RECT 1628.560 82.870 1628.700 126.830 ;
        RECT 1628.560 82.730 1631.920 82.870 ;
        RECT 1631.780 1.770 1631.920 82.730 ;
        RECT 1633.870 1.770 1634.430 2.400 ;
        RECT 1631.780 1.630 1634.430 1.770 ;
        RECT 1633.870 -4.800 1634.430 1.630 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 698.350 127.400 698.670 127.460 ;
        RECT 1649.170 127.400 1649.490 127.460 ;
        RECT 698.350 127.260 1649.490 127.400 ;
        RECT 698.350 127.200 698.670 127.260 ;
        RECT 1649.170 127.200 1649.490 127.260 ;
      LAYER via ;
        RECT 698.380 127.200 698.640 127.460 ;
        RECT 1649.200 127.200 1649.460 127.460 ;
      LAYER met2 ;
        RECT 698.730 400.250 699.010 404.000 ;
        RECT 698.440 400.110 699.010 400.250 ;
        RECT 698.440 127.490 698.580 400.110 ;
        RECT 698.730 400.000 699.010 400.110 ;
        RECT 698.380 127.170 698.640 127.490 ;
        RECT 1649.200 127.170 1649.460 127.490 ;
        RECT 1649.260 82.870 1649.400 127.170 ;
        RECT 1649.260 82.730 1652.160 82.870 ;
        RECT 1652.020 2.400 1652.160 82.730 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.410 385.460 703.730 385.520 ;
        RECT 704.790 385.460 705.110 385.520 ;
        RECT 703.410 385.320 705.110 385.460 ;
        RECT 703.410 385.260 703.730 385.320 ;
        RECT 704.790 385.260 705.110 385.320 ;
        RECT 704.790 131.140 705.110 131.200 ;
        RECT 1662.970 131.140 1663.290 131.200 ;
        RECT 704.790 131.000 1663.290 131.140 ;
        RECT 704.790 130.940 705.110 131.000 ;
        RECT 1662.970 130.940 1663.290 131.000 ;
        RECT 1662.970 15.200 1663.290 15.260 ;
        RECT 1669.410 15.200 1669.730 15.260 ;
        RECT 1662.970 15.060 1669.730 15.200 ;
        RECT 1662.970 15.000 1663.290 15.060 ;
        RECT 1669.410 15.000 1669.730 15.060 ;
      LAYER via ;
        RECT 703.440 385.260 703.700 385.520 ;
        RECT 704.820 385.260 705.080 385.520 ;
        RECT 704.820 130.940 705.080 131.200 ;
        RECT 1663.000 130.940 1663.260 131.200 ;
        RECT 1663.000 15.000 1663.260 15.260 ;
        RECT 1669.440 15.000 1669.700 15.260 ;
      LAYER met2 ;
        RECT 703.790 400.180 704.070 404.000 ;
        RECT 703.790 400.000 704.100 400.180 ;
        RECT 703.960 388.690 704.100 400.000 ;
        RECT 703.500 388.550 704.100 388.690 ;
        RECT 703.500 385.550 703.640 388.550 ;
        RECT 703.440 385.230 703.700 385.550 ;
        RECT 704.820 385.230 705.080 385.550 ;
        RECT 704.880 131.230 705.020 385.230 ;
        RECT 704.820 130.910 705.080 131.230 ;
        RECT 1663.000 130.910 1663.260 131.230 ;
        RECT 1663.060 15.290 1663.200 130.910 ;
        RECT 1663.000 14.970 1663.260 15.290 ;
        RECT 1669.440 14.970 1669.700 15.290 ;
        RECT 1669.500 2.400 1669.640 14.970 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 705.250 130.800 705.570 130.860 ;
        RECT 1683.670 130.800 1683.990 130.860 ;
        RECT 705.250 130.660 1683.990 130.800 ;
        RECT 705.250 130.600 705.570 130.660 ;
        RECT 1683.670 130.600 1683.990 130.660 ;
      LAYER via ;
        RECT 705.280 130.600 705.540 130.860 ;
        RECT 1683.700 130.600 1683.960 130.860 ;
      LAYER met2 ;
        RECT 709.310 400.250 709.590 404.000 ;
        RECT 708.100 400.110 709.590 400.250 ;
        RECT 708.100 324.370 708.240 400.110 ;
        RECT 709.310 400.000 709.590 400.110 ;
        RECT 705.340 324.230 708.240 324.370 ;
        RECT 705.340 130.890 705.480 324.230 ;
        RECT 705.280 130.570 705.540 130.890 ;
        RECT 1683.700 130.570 1683.960 130.890 ;
        RECT 1683.760 82.870 1683.900 130.570 ;
        RECT 1683.760 82.730 1685.280 82.870 ;
        RECT 1685.140 1.770 1685.280 82.730 ;
        RECT 1687.230 1.770 1687.790 2.400 ;
        RECT 1685.140 1.630 1687.790 1.770 ;
        RECT 1687.230 -4.800 1687.790 1.630 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.990 386.480 415.310 386.540 ;
        RECT 418.670 386.480 418.990 386.540 ;
        RECT 414.990 386.340 418.990 386.480 ;
        RECT 414.990 386.280 415.310 386.340 ;
        RECT 418.670 386.280 418.990 386.340 ;
        RECT 414.990 33.900 415.310 33.960 ;
        RECT 552.530 33.900 552.850 33.960 ;
        RECT 414.990 33.760 552.850 33.900 ;
        RECT 414.990 33.700 415.310 33.760 ;
        RECT 552.530 33.700 552.850 33.760 ;
        RECT 552.530 20.300 552.850 20.360 ;
        RECT 729.630 20.300 729.950 20.360 ;
        RECT 552.530 20.160 729.950 20.300 ;
        RECT 552.530 20.100 552.850 20.160 ;
        RECT 729.630 20.100 729.950 20.160 ;
      LAYER via ;
        RECT 415.020 386.280 415.280 386.540 ;
        RECT 418.700 386.280 418.960 386.540 ;
        RECT 415.020 33.700 415.280 33.960 ;
        RECT 552.560 33.700 552.820 33.960 ;
        RECT 552.560 20.100 552.820 20.360 ;
        RECT 729.660 20.100 729.920 20.360 ;
      LAYER met2 ;
        RECT 419.970 400.250 420.250 404.000 ;
        RECT 418.760 400.110 420.250 400.250 ;
        RECT 418.760 386.570 418.900 400.110 ;
        RECT 419.970 400.000 420.250 400.110 ;
        RECT 415.020 386.250 415.280 386.570 ;
        RECT 418.700 386.250 418.960 386.570 ;
        RECT 415.080 33.990 415.220 386.250 ;
        RECT 415.020 33.670 415.280 33.990 ;
        RECT 552.560 33.670 552.820 33.990 ;
        RECT 552.620 20.390 552.760 33.670 ;
        RECT 552.560 20.070 552.820 20.390 ;
        RECT 729.660 20.070 729.920 20.390 ;
        RECT 729.720 2.400 729.860 20.070 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 712.150 130.460 712.470 130.520 ;
        RECT 1704.370 130.460 1704.690 130.520 ;
        RECT 712.150 130.320 1704.690 130.460 ;
        RECT 712.150 130.260 712.470 130.320 ;
        RECT 1704.370 130.260 1704.690 130.320 ;
      LAYER via ;
        RECT 712.180 130.260 712.440 130.520 ;
        RECT 1704.400 130.260 1704.660 130.520 ;
      LAYER met2 ;
        RECT 714.830 400.250 715.110 404.000 ;
        RECT 713.620 400.110 715.110 400.250 ;
        RECT 713.620 324.370 713.760 400.110 ;
        RECT 714.830 400.000 715.110 400.110 ;
        RECT 712.240 324.230 713.760 324.370 ;
        RECT 712.240 130.550 712.380 324.230 ;
        RECT 712.180 130.230 712.440 130.550 ;
        RECT 1704.400 130.230 1704.660 130.550 ;
        RECT 1704.460 82.870 1704.600 130.230 ;
        RECT 1704.460 82.730 1705.060 82.870 ;
        RECT 1704.920 2.400 1705.060 82.730 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 719.050 130.120 719.370 130.180 ;
        RECT 1718.170 130.120 1718.490 130.180 ;
        RECT 719.050 129.980 1718.490 130.120 ;
        RECT 719.050 129.920 719.370 129.980 ;
        RECT 1718.170 129.920 1718.490 129.980 ;
      LAYER via ;
        RECT 719.080 129.920 719.340 130.180 ;
        RECT 1718.200 129.920 1718.460 130.180 ;
      LAYER met2 ;
        RECT 719.890 400.250 720.170 404.000 ;
        RECT 719.140 400.110 720.170 400.250 ;
        RECT 719.140 130.210 719.280 400.110 ;
        RECT 719.890 400.000 720.170 400.110 ;
        RECT 719.080 129.890 719.340 130.210 ;
        RECT 1718.200 129.890 1718.460 130.210 ;
        RECT 1718.260 82.870 1718.400 129.890 ;
        RECT 1718.260 82.730 1723.000 82.870 ;
        RECT 1722.860 2.400 1723.000 82.730 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.490 129.780 725.810 129.840 ;
        RECT 1738.870 129.780 1739.190 129.840 ;
        RECT 725.490 129.640 1739.190 129.780 ;
        RECT 725.490 129.580 725.810 129.640 ;
        RECT 1738.870 129.580 1739.190 129.640 ;
      LAYER via ;
        RECT 725.520 129.580 725.780 129.840 ;
        RECT 1738.900 129.580 1739.160 129.840 ;
      LAYER met2 ;
        RECT 725.410 400.180 725.690 404.000 ;
        RECT 725.410 400.000 725.720 400.180 ;
        RECT 725.580 129.870 725.720 400.000 ;
        RECT 725.520 129.550 725.780 129.870 ;
        RECT 1738.900 129.550 1739.160 129.870 ;
        RECT 1738.960 82.870 1739.100 129.550 ;
        RECT 1738.960 82.730 1740.480 82.870 ;
        RECT 1740.340 2.400 1740.480 82.730 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.950 385.800 726.270 385.860 ;
        RECT 729.630 385.800 729.950 385.860 ;
        RECT 725.950 385.660 729.950 385.800 ;
        RECT 725.950 385.600 726.270 385.660 ;
        RECT 729.630 385.600 729.950 385.660 ;
        RECT 725.950 129.440 726.270 129.500 ;
        RECT 1752.670 129.440 1752.990 129.500 ;
        RECT 725.950 129.300 1752.990 129.440 ;
        RECT 725.950 129.240 726.270 129.300 ;
        RECT 1752.670 129.240 1752.990 129.300 ;
      LAYER via ;
        RECT 725.980 385.600 726.240 385.860 ;
        RECT 729.660 385.600 729.920 385.860 ;
        RECT 725.980 129.240 726.240 129.500 ;
        RECT 1752.700 129.240 1752.960 129.500 ;
      LAYER met2 ;
        RECT 730.930 400.250 731.210 404.000 ;
        RECT 729.720 400.110 731.210 400.250 ;
        RECT 729.720 385.890 729.860 400.110 ;
        RECT 730.930 400.000 731.210 400.110 ;
        RECT 725.980 385.570 726.240 385.890 ;
        RECT 729.660 385.570 729.920 385.890 ;
        RECT 726.040 129.530 726.180 385.570 ;
        RECT 725.980 129.210 726.240 129.530 ;
        RECT 1752.700 129.210 1752.960 129.530 ;
        RECT 1752.760 82.870 1752.900 129.210 ;
        RECT 1752.760 82.730 1756.120 82.870 ;
        RECT 1755.980 1.770 1756.120 82.730 ;
        RECT 1758.070 1.770 1758.630 2.400 ;
        RECT 1755.980 1.630 1758.630 1.770 ;
        RECT 1758.070 -4.800 1758.630 1.630 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.850 129.100 733.170 129.160 ;
        RECT 1773.370 129.100 1773.690 129.160 ;
        RECT 732.850 128.960 1773.690 129.100 ;
        RECT 732.850 128.900 733.170 128.960 ;
        RECT 1773.370 128.900 1773.690 128.960 ;
      LAYER via ;
        RECT 732.880 128.900 733.140 129.160 ;
        RECT 1773.400 128.900 1773.660 129.160 ;
      LAYER met2 ;
        RECT 735.990 400.250 736.270 404.000 ;
        RECT 734.780 400.110 736.270 400.250 ;
        RECT 734.780 324.370 734.920 400.110 ;
        RECT 735.990 400.000 736.270 400.110 ;
        RECT 732.940 324.230 734.920 324.370 ;
        RECT 732.940 129.190 733.080 324.230 ;
        RECT 732.880 128.870 733.140 129.190 ;
        RECT 1773.400 128.870 1773.660 129.190 ;
        RECT 1773.460 82.870 1773.600 128.870 ;
        RECT 1773.460 82.730 1776.360 82.870 ;
        RECT 1776.220 2.400 1776.360 82.730 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 739.290 128.760 739.610 128.820 ;
        RECT 1787.170 128.760 1787.490 128.820 ;
        RECT 739.290 128.620 1787.490 128.760 ;
        RECT 739.290 128.560 739.610 128.620 ;
        RECT 1787.170 128.560 1787.490 128.620 ;
        RECT 1787.170 15.200 1787.490 15.260 ;
        RECT 1793.610 15.200 1793.930 15.260 ;
        RECT 1787.170 15.060 1793.930 15.200 ;
        RECT 1787.170 15.000 1787.490 15.060 ;
        RECT 1793.610 15.000 1793.930 15.060 ;
      LAYER via ;
        RECT 739.320 128.560 739.580 128.820 ;
        RECT 1787.200 128.560 1787.460 128.820 ;
        RECT 1787.200 15.000 1787.460 15.260 ;
        RECT 1793.640 15.000 1793.900 15.260 ;
      LAYER met2 ;
        RECT 741.510 400.250 741.790 404.000 ;
        RECT 740.300 400.110 741.790 400.250 ;
        RECT 740.300 324.370 740.440 400.110 ;
        RECT 741.510 400.000 741.790 400.110 ;
        RECT 739.380 324.230 740.440 324.370 ;
        RECT 739.380 128.850 739.520 324.230 ;
        RECT 739.320 128.530 739.580 128.850 ;
        RECT 1787.200 128.530 1787.460 128.850 ;
        RECT 1787.260 15.290 1787.400 128.530 ;
        RECT 1787.200 14.970 1787.460 15.290 ;
        RECT 1793.640 14.970 1793.900 15.290 ;
        RECT 1793.700 2.400 1793.840 14.970 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 746.650 128.420 746.970 128.480 ;
        RECT 1807.870 128.420 1808.190 128.480 ;
        RECT 746.650 128.280 1808.190 128.420 ;
        RECT 746.650 128.220 746.970 128.280 ;
        RECT 1807.870 128.220 1808.190 128.280 ;
      LAYER via ;
        RECT 746.680 128.220 746.940 128.480 ;
        RECT 1807.900 128.220 1808.160 128.480 ;
      LAYER met2 ;
        RECT 747.030 400.250 747.310 404.000 ;
        RECT 746.740 400.110 747.310 400.250 ;
        RECT 746.740 128.510 746.880 400.110 ;
        RECT 747.030 400.000 747.310 400.110 ;
        RECT 746.680 128.190 746.940 128.510 ;
        RECT 1807.900 128.190 1808.160 128.510 ;
        RECT 1807.960 82.870 1808.100 128.190 ;
        RECT 1807.960 82.730 1809.480 82.870 ;
        RECT 1809.340 1.770 1809.480 82.730 ;
        RECT 1811.430 1.770 1811.990 2.400 ;
        RECT 1809.340 1.630 1811.990 1.770 ;
        RECT 1811.430 -4.800 1811.990 1.630 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.170 392.600 752.490 392.660 ;
        RECT 1828.570 392.600 1828.890 392.660 ;
        RECT 752.170 392.460 1828.890 392.600 ;
        RECT 752.170 392.400 752.490 392.460 ;
        RECT 1828.570 392.400 1828.890 392.460 ;
      LAYER via ;
        RECT 752.200 392.400 752.460 392.660 ;
        RECT 1828.600 392.400 1828.860 392.660 ;
      LAYER met2 ;
        RECT 752.090 400.180 752.370 404.000 ;
        RECT 752.090 400.000 752.400 400.180 ;
        RECT 752.260 392.690 752.400 400.000 ;
        RECT 752.200 392.370 752.460 392.690 ;
        RECT 1828.600 392.370 1828.860 392.690 ;
        RECT 1828.660 82.870 1828.800 392.370 ;
        RECT 1828.660 82.730 1829.260 82.870 ;
        RECT 1829.120 2.400 1829.260 82.730 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 753.090 128.080 753.410 128.140 ;
        RECT 1842.370 128.080 1842.690 128.140 ;
        RECT 753.090 127.940 1842.690 128.080 ;
        RECT 753.090 127.880 753.410 127.940 ;
        RECT 1842.370 127.880 1842.690 127.940 ;
      LAYER via ;
        RECT 753.120 127.880 753.380 128.140 ;
        RECT 1842.400 127.880 1842.660 128.140 ;
      LAYER met2 ;
        RECT 757.610 400.250 757.890 404.000 ;
        RECT 756.400 400.110 757.890 400.250 ;
        RECT 756.400 390.730 756.540 400.110 ;
        RECT 757.610 400.000 757.890 400.110 ;
        RECT 755.020 390.590 756.540 390.730 ;
        RECT 755.020 324.370 755.160 390.590 ;
        RECT 753.180 324.230 755.160 324.370 ;
        RECT 753.180 128.170 753.320 324.230 ;
        RECT 753.120 127.850 753.380 128.170 ;
        RECT 1842.400 127.850 1842.660 128.170 ;
        RECT 1842.460 82.870 1842.600 127.850 ;
        RECT 1842.460 82.730 1847.200 82.870 ;
        RECT 1847.060 2.400 1847.200 82.730 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 763.210 392.260 763.530 392.320 ;
        RECT 1863.070 392.260 1863.390 392.320 ;
        RECT 763.210 392.120 1863.390 392.260 ;
        RECT 763.210 392.060 763.530 392.120 ;
        RECT 1863.070 392.060 1863.390 392.120 ;
      LAYER via ;
        RECT 763.240 392.060 763.500 392.320 ;
        RECT 1863.100 392.060 1863.360 392.320 ;
      LAYER met2 ;
        RECT 763.130 400.180 763.410 404.000 ;
        RECT 763.130 400.000 763.440 400.180 ;
        RECT 763.300 392.350 763.440 400.000 ;
        RECT 763.240 392.030 763.500 392.350 ;
        RECT 1863.100 392.030 1863.360 392.350 ;
        RECT 1863.160 82.870 1863.300 392.030 ;
        RECT 1863.160 82.730 1864.680 82.870 ;
        RECT 1864.540 2.400 1864.680 82.730 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 386.480 421.290 386.540 ;
        RECT 424.190 386.480 424.510 386.540 ;
        RECT 420.970 386.340 424.510 386.480 ;
        RECT 420.970 386.280 421.290 386.340 ;
        RECT 424.190 386.280 424.510 386.340 ;
        RECT 420.970 17.580 421.290 17.640 ;
        RECT 747.570 17.580 747.890 17.640 ;
        RECT 420.970 17.440 440.980 17.580 ;
        RECT 420.970 17.380 421.290 17.440 ;
        RECT 440.840 17.240 440.980 17.440 ;
        RECT 452.340 17.440 747.890 17.580 ;
        RECT 452.340 17.240 452.480 17.440 ;
        RECT 747.570 17.380 747.890 17.440 ;
        RECT 440.840 17.100 452.480 17.240 ;
      LAYER via ;
        RECT 421.000 386.280 421.260 386.540 ;
        RECT 424.220 386.280 424.480 386.540 ;
        RECT 421.000 17.380 421.260 17.640 ;
        RECT 747.600 17.380 747.860 17.640 ;
      LAYER met2 ;
        RECT 425.490 400.250 425.770 404.000 ;
        RECT 424.280 400.110 425.770 400.250 ;
        RECT 424.280 386.570 424.420 400.110 ;
        RECT 425.490 400.000 425.770 400.110 ;
        RECT 421.000 386.250 421.260 386.570 ;
        RECT 424.220 386.250 424.480 386.570 ;
        RECT 421.060 17.670 421.200 386.250 ;
        RECT 421.000 17.350 421.260 17.670 ;
        RECT 747.600 17.350 747.860 17.670 ;
        RECT 747.660 2.400 747.800 17.350 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 767.350 127.740 767.670 127.800 ;
        RECT 1876.870 127.740 1877.190 127.800 ;
        RECT 767.350 127.600 1877.190 127.740 ;
        RECT 767.350 127.540 767.670 127.600 ;
        RECT 1876.870 127.540 1877.190 127.600 ;
      LAYER via ;
        RECT 767.380 127.540 767.640 127.800 ;
        RECT 1876.900 127.540 1877.160 127.800 ;
      LAYER met2 ;
        RECT 768.190 400.250 768.470 404.000 ;
        RECT 767.440 400.110 768.470 400.250 ;
        RECT 767.440 127.830 767.580 400.110 ;
        RECT 768.190 400.000 768.470 400.110 ;
        RECT 767.380 127.510 767.640 127.830 ;
        RECT 1876.900 127.510 1877.160 127.830 ;
        RECT 1876.960 82.870 1877.100 127.510 ;
        RECT 1876.960 82.730 1880.320 82.870 ;
        RECT 1880.180 1.770 1880.320 82.730 ;
        RECT 1882.270 1.770 1882.830 2.400 ;
        RECT 1880.180 1.630 1882.830 1.770 ;
        RECT 1882.270 -4.800 1882.830 1.630 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.790 391.920 774.110 391.980 ;
        RECT 1897.570 391.920 1897.890 391.980 ;
        RECT 773.790 391.780 1897.890 391.920 ;
        RECT 773.790 391.720 774.110 391.780 ;
        RECT 1897.570 391.720 1897.890 391.780 ;
      LAYER via ;
        RECT 773.820 391.720 774.080 391.980 ;
        RECT 1897.600 391.720 1897.860 391.980 ;
      LAYER met2 ;
        RECT 773.710 400.180 773.990 404.000 ;
        RECT 773.710 400.000 774.020 400.180 ;
        RECT 773.880 392.010 774.020 400.000 ;
        RECT 773.820 391.690 774.080 392.010 ;
        RECT 1897.600 391.690 1897.860 392.010 ;
        RECT 1897.660 1.770 1897.800 391.690 ;
        RECT 1899.750 1.770 1900.310 2.400 ;
        RECT 1897.660 1.630 1900.310 1.770 ;
        RECT 1899.750 -4.800 1900.310 1.630 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.790 136.240 774.110 136.300 ;
        RECT 1911.370 136.240 1911.690 136.300 ;
        RECT 773.790 136.100 1911.690 136.240 ;
        RECT 773.790 136.040 774.110 136.100 ;
        RECT 1911.370 136.040 1911.690 136.100 ;
        RECT 1911.370 15.200 1911.690 15.260 ;
        RECT 1917.810 15.200 1918.130 15.260 ;
        RECT 1911.370 15.060 1918.130 15.200 ;
        RECT 1911.370 15.000 1911.690 15.060 ;
        RECT 1917.810 15.000 1918.130 15.060 ;
      LAYER via ;
        RECT 773.820 136.040 774.080 136.300 ;
        RECT 1911.400 136.040 1911.660 136.300 ;
        RECT 1911.400 15.000 1911.660 15.260 ;
        RECT 1917.840 15.000 1918.100 15.260 ;
      LAYER met2 ;
        RECT 779.230 400.250 779.510 404.000 ;
        RECT 778.020 400.110 779.510 400.250 ;
        RECT 778.020 324.370 778.160 400.110 ;
        RECT 779.230 400.000 779.510 400.110 ;
        RECT 773.880 324.230 778.160 324.370 ;
        RECT 773.880 136.330 774.020 324.230 ;
        RECT 773.820 136.010 774.080 136.330 ;
        RECT 1911.400 136.010 1911.660 136.330 ;
        RECT 1911.460 15.290 1911.600 136.010 ;
        RECT 1911.400 14.970 1911.660 15.290 ;
        RECT 1917.840 14.970 1918.100 15.290 ;
        RECT 1917.900 2.400 1918.040 14.970 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 784.370 391.580 784.690 391.640 ;
        RECT 1932.070 391.580 1932.390 391.640 ;
        RECT 784.370 391.440 1932.390 391.580 ;
        RECT 784.370 391.380 784.690 391.440 ;
        RECT 1932.070 391.380 1932.390 391.440 ;
      LAYER via ;
        RECT 784.400 391.380 784.660 391.640 ;
        RECT 1932.100 391.380 1932.360 391.640 ;
      LAYER met2 ;
        RECT 784.290 400.180 784.570 404.000 ;
        RECT 784.290 400.000 784.600 400.180 ;
        RECT 784.460 391.670 784.600 400.000 ;
        RECT 784.400 391.350 784.660 391.670 ;
        RECT 1932.100 391.350 1932.360 391.670 ;
        RECT 1932.160 82.870 1932.300 391.350 ;
        RECT 1932.160 82.730 1933.680 82.870 ;
        RECT 1933.540 1.770 1933.680 82.730 ;
        RECT 1935.630 1.770 1936.190 2.400 ;
        RECT 1933.540 1.630 1936.190 1.770 ;
        RECT 1935.630 -4.800 1936.190 1.630 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.590 135.900 787.910 135.960 ;
        RECT 1952.770 135.900 1953.090 135.960 ;
        RECT 787.590 135.760 1953.090 135.900 ;
        RECT 787.590 135.700 787.910 135.760 ;
        RECT 1952.770 135.700 1953.090 135.760 ;
      LAYER via ;
        RECT 787.620 135.700 787.880 135.960 ;
        RECT 1952.800 135.700 1953.060 135.960 ;
      LAYER met2 ;
        RECT 789.810 400.250 790.090 404.000 ;
        RECT 788.600 400.110 790.090 400.250 ;
        RECT 788.600 324.370 788.740 400.110 ;
        RECT 789.810 400.000 790.090 400.110 ;
        RECT 787.680 324.230 788.740 324.370 ;
        RECT 787.680 135.990 787.820 324.230 ;
        RECT 787.620 135.670 787.880 135.990 ;
        RECT 1952.800 135.670 1953.060 135.990 ;
        RECT 1952.860 82.870 1953.000 135.670 ;
        RECT 1952.860 82.730 1953.460 82.870 ;
        RECT 1953.320 2.400 1953.460 82.730 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 795.410 391.240 795.730 391.300 ;
        RECT 1966.570 391.240 1966.890 391.300 ;
        RECT 795.410 391.100 1966.890 391.240 ;
        RECT 795.410 391.040 795.730 391.100 ;
        RECT 1966.570 391.040 1966.890 391.100 ;
      LAYER via ;
        RECT 795.440 391.040 795.700 391.300 ;
        RECT 1966.600 391.040 1966.860 391.300 ;
      LAYER met2 ;
        RECT 795.330 400.180 795.610 404.000 ;
        RECT 795.330 400.000 795.640 400.180 ;
        RECT 795.500 391.330 795.640 400.000 ;
        RECT 795.440 391.010 795.700 391.330 ;
        RECT 1966.600 391.010 1966.860 391.330 ;
        RECT 1966.660 82.870 1966.800 391.010 ;
        RECT 1966.660 82.730 1971.400 82.870 ;
        RECT 1971.260 2.400 1971.400 82.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.010 384.780 800.330 384.840 ;
        RECT 801.390 384.780 801.710 384.840 ;
        RECT 800.010 384.640 801.710 384.780 ;
        RECT 800.010 384.580 800.330 384.640 ;
        RECT 801.390 384.580 801.710 384.640 ;
        RECT 801.390 135.560 801.710 135.620 ;
        RECT 1987.270 135.560 1987.590 135.620 ;
        RECT 801.390 135.420 1987.590 135.560 ;
        RECT 801.390 135.360 801.710 135.420 ;
        RECT 1987.270 135.360 1987.590 135.420 ;
      LAYER via ;
        RECT 800.040 384.580 800.300 384.840 ;
        RECT 801.420 384.580 801.680 384.840 ;
        RECT 801.420 135.360 801.680 135.620 ;
        RECT 1987.300 135.360 1987.560 135.620 ;
      LAYER met2 ;
        RECT 800.390 400.180 800.670 404.000 ;
        RECT 800.390 400.000 800.700 400.180 ;
        RECT 800.560 386.470 800.700 400.000 ;
        RECT 800.100 386.330 800.700 386.470 ;
        RECT 800.100 384.870 800.240 386.330 ;
        RECT 800.040 384.550 800.300 384.870 ;
        RECT 801.420 384.550 801.680 384.870 ;
        RECT 801.480 135.650 801.620 384.550 ;
        RECT 801.420 135.330 801.680 135.650 ;
        RECT 1987.300 135.330 1987.560 135.650 ;
        RECT 1987.360 82.870 1987.500 135.330 ;
        RECT 1987.360 82.730 1988.880 82.870 ;
        RECT 1988.740 2.400 1988.880 82.730 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 805.990 390.900 806.310 390.960 ;
        RECT 2001.070 390.900 2001.390 390.960 ;
        RECT 805.990 390.760 2001.390 390.900 ;
        RECT 805.990 390.700 806.310 390.760 ;
        RECT 2001.070 390.700 2001.390 390.760 ;
      LAYER via ;
        RECT 806.020 390.700 806.280 390.960 ;
        RECT 2001.100 390.700 2001.360 390.960 ;
      LAYER met2 ;
        RECT 805.910 400.180 806.190 404.000 ;
        RECT 805.910 400.000 806.220 400.180 ;
        RECT 806.080 390.990 806.220 400.000 ;
        RECT 806.020 390.670 806.280 390.990 ;
        RECT 2001.100 390.670 2001.360 390.990 ;
        RECT 2001.160 82.870 2001.300 390.670 ;
        RECT 2001.160 82.730 2004.520 82.870 ;
        RECT 2004.380 1.770 2004.520 82.730 ;
        RECT 2006.470 1.770 2007.030 2.400 ;
        RECT 2004.380 1.630 2007.030 1.770 ;
        RECT 2006.470 -4.800 2007.030 1.630 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 808.750 135.220 809.070 135.280 ;
        RECT 2021.770 135.220 2022.090 135.280 ;
        RECT 808.750 135.080 2022.090 135.220 ;
        RECT 808.750 135.020 809.070 135.080 ;
        RECT 2021.770 135.020 2022.090 135.080 ;
      LAYER via ;
        RECT 808.780 135.020 809.040 135.280 ;
        RECT 2021.800 135.020 2022.060 135.280 ;
      LAYER met2 ;
        RECT 810.970 400.250 811.250 404.000 ;
        RECT 810.220 400.110 811.250 400.250 ;
        RECT 810.220 324.370 810.360 400.110 ;
        RECT 810.970 400.000 811.250 400.110 ;
        RECT 808.840 324.230 810.360 324.370 ;
        RECT 808.840 135.310 808.980 324.230 ;
        RECT 808.780 134.990 809.040 135.310 ;
        RECT 2021.800 134.990 2022.060 135.310 ;
        RECT 2021.860 1.770 2022.000 134.990 ;
        RECT 2023.950 1.770 2024.510 2.400 ;
        RECT 2021.860 1.630 2024.510 1.770 ;
        RECT 2023.950 -4.800 2024.510 1.630 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 816.570 390.560 816.890 390.620 ;
        RECT 2035.570 390.560 2035.890 390.620 ;
        RECT 816.570 390.420 2035.890 390.560 ;
        RECT 816.570 390.360 816.890 390.420 ;
        RECT 2035.570 390.360 2035.890 390.420 ;
        RECT 2035.570 15.200 2035.890 15.260 ;
        RECT 2042.010 15.200 2042.330 15.260 ;
        RECT 2035.570 15.060 2042.330 15.200 ;
        RECT 2035.570 15.000 2035.890 15.060 ;
        RECT 2042.010 15.000 2042.330 15.060 ;
      LAYER via ;
        RECT 816.600 390.360 816.860 390.620 ;
        RECT 2035.600 390.360 2035.860 390.620 ;
        RECT 2035.600 15.000 2035.860 15.260 ;
        RECT 2042.040 15.000 2042.300 15.260 ;
      LAYER met2 ;
        RECT 816.490 400.180 816.770 404.000 ;
        RECT 816.490 400.000 816.800 400.180 ;
        RECT 816.660 390.650 816.800 400.000 ;
        RECT 816.600 390.330 816.860 390.650 ;
        RECT 2035.600 390.330 2035.860 390.650 ;
        RECT 2035.660 15.290 2035.800 390.330 ;
        RECT 2035.600 14.970 2035.860 15.290 ;
        RECT 2042.040 14.970 2042.300 15.290 ;
        RECT 2042.100 2.400 2042.240 14.970 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 386.480 428.190 386.540 ;
        RECT 429.710 386.480 430.030 386.540 ;
        RECT 427.870 386.340 430.030 386.480 ;
        RECT 427.870 386.280 428.190 386.340 ;
        RECT 429.710 386.280 430.030 386.340 ;
        RECT 765.050 17.240 765.370 17.300 ;
        RECT 452.800 17.100 765.370 17.240 ;
        RECT 427.870 16.220 428.190 16.280 ;
        RECT 452.800 16.220 452.940 17.100 ;
        RECT 765.050 17.040 765.370 17.100 ;
        RECT 427.870 16.080 452.940 16.220 ;
        RECT 427.870 16.020 428.190 16.080 ;
      LAYER via ;
        RECT 427.900 386.280 428.160 386.540 ;
        RECT 429.740 386.280 430.000 386.540 ;
        RECT 427.900 16.020 428.160 16.280 ;
        RECT 765.080 17.040 765.340 17.300 ;
      LAYER met2 ;
        RECT 430.550 400.250 430.830 404.000 ;
        RECT 429.800 400.110 430.830 400.250 ;
        RECT 429.800 386.570 429.940 400.110 ;
        RECT 430.550 400.000 430.830 400.110 ;
        RECT 427.900 386.250 428.160 386.570 ;
        RECT 429.740 386.250 430.000 386.570 ;
        RECT 427.960 16.310 428.100 386.250 ;
        RECT 765.080 17.010 765.340 17.330 ;
        RECT 427.900 15.990 428.160 16.310 ;
        RECT 765.140 2.400 765.280 17.010 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 822.090 134.880 822.410 134.940 ;
        RECT 2056.270 134.880 2056.590 134.940 ;
        RECT 822.090 134.740 2056.590 134.880 ;
        RECT 822.090 134.680 822.410 134.740 ;
        RECT 2056.270 134.680 2056.590 134.740 ;
      LAYER via ;
        RECT 822.120 134.680 822.380 134.940 ;
        RECT 2056.300 134.680 2056.560 134.940 ;
      LAYER met2 ;
        RECT 822.010 400.180 822.290 404.000 ;
        RECT 822.010 400.000 822.320 400.180 ;
        RECT 822.180 134.970 822.320 400.000 ;
        RECT 822.120 134.650 822.380 134.970 ;
        RECT 2056.300 134.650 2056.560 134.970 ;
        RECT 2056.360 82.870 2056.500 134.650 ;
        RECT 2056.360 82.730 2059.720 82.870 ;
        RECT 2059.580 2.400 2059.720 82.730 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 827.150 390.220 827.470 390.280 ;
        RECT 2076.970 390.220 2077.290 390.280 ;
        RECT 827.150 390.080 2077.290 390.220 ;
        RECT 827.150 390.020 827.470 390.080 ;
        RECT 2076.970 390.020 2077.290 390.080 ;
      LAYER via ;
        RECT 827.180 390.020 827.440 390.280 ;
        RECT 2077.000 390.020 2077.260 390.280 ;
      LAYER met2 ;
        RECT 827.070 400.180 827.350 404.000 ;
        RECT 827.070 400.000 827.380 400.180 ;
        RECT 827.240 390.310 827.380 400.000 ;
        RECT 827.180 389.990 827.440 390.310 ;
        RECT 2077.000 389.990 2077.260 390.310 ;
        RECT 2077.060 82.870 2077.200 389.990 ;
        RECT 2077.060 82.730 2077.660 82.870 ;
        RECT 2077.520 2.400 2077.660 82.730 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 829.450 134.540 829.770 134.600 ;
        RECT 2090.770 134.540 2091.090 134.600 ;
        RECT 829.450 134.400 2091.090 134.540 ;
        RECT 829.450 134.340 829.770 134.400 ;
        RECT 2090.770 134.340 2091.090 134.400 ;
      LAYER via ;
        RECT 829.480 134.340 829.740 134.600 ;
        RECT 2090.800 134.340 2091.060 134.600 ;
      LAYER met2 ;
        RECT 832.590 400.250 832.870 404.000 ;
        RECT 831.380 400.110 832.870 400.250 ;
        RECT 831.380 324.370 831.520 400.110 ;
        RECT 832.590 400.000 832.870 400.110 ;
        RECT 829.540 324.230 831.520 324.370 ;
        RECT 829.540 134.630 829.680 324.230 ;
        RECT 829.480 134.310 829.740 134.630 ;
        RECT 2090.800 134.310 2091.060 134.630 ;
        RECT 2090.860 82.870 2091.000 134.310 ;
        RECT 2090.860 82.730 2092.840 82.870 ;
        RECT 2092.700 1.770 2092.840 82.730 ;
        RECT 2094.790 1.770 2095.350 2.400 ;
        RECT 2092.700 1.630 2095.350 1.770 ;
        RECT 2094.790 -4.800 2095.350 1.630 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 838.190 389.880 838.510 389.940 ;
        RECT 2111.470 389.880 2111.790 389.940 ;
        RECT 838.190 389.740 2111.790 389.880 ;
        RECT 838.190 389.680 838.510 389.740 ;
        RECT 2111.470 389.680 2111.790 389.740 ;
      LAYER via ;
        RECT 838.220 389.680 838.480 389.940 ;
        RECT 2111.500 389.680 2111.760 389.940 ;
      LAYER met2 ;
        RECT 838.110 400.180 838.390 404.000 ;
        RECT 838.110 400.000 838.420 400.180 ;
        RECT 838.280 389.970 838.420 400.000 ;
        RECT 838.220 389.650 838.480 389.970 ;
        RECT 2111.500 389.650 2111.760 389.970 ;
        RECT 2111.560 82.870 2111.700 389.650 ;
        RECT 2111.560 82.730 2113.080 82.870 ;
        RECT 2112.940 2.400 2113.080 82.730 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.330 15.540 842.650 15.600 ;
        RECT 842.330 15.400 2063.170 15.540 ;
        RECT 842.330 15.340 842.650 15.400 ;
        RECT 2063.030 14.860 2063.170 15.400 ;
        RECT 2130.790 14.860 2131.110 14.920 ;
        RECT 2063.030 14.720 2131.110 14.860 ;
        RECT 2130.790 14.660 2131.110 14.720 ;
      LAYER via ;
        RECT 842.360 15.340 842.620 15.600 ;
        RECT 2130.820 14.660 2131.080 14.920 ;
      LAYER met2 ;
        RECT 843.170 400.250 843.450 404.000 ;
        RECT 841.960 400.110 843.450 400.250 ;
        RECT 841.960 34.570 842.100 400.110 ;
        RECT 843.170 400.000 843.450 400.110 ;
        RECT 841.960 34.430 842.560 34.570 ;
        RECT 842.420 15.630 842.560 34.430 ;
        RECT 842.360 15.310 842.620 15.630 ;
        RECT 2130.820 14.630 2131.080 14.950 ;
        RECT 2130.880 2.400 2131.020 14.630 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 848.770 15.880 849.090 15.940 ;
        RECT 848.770 15.740 2118.140 15.880 ;
        RECT 848.770 15.680 849.090 15.740 ;
        RECT 2118.000 15.200 2118.140 15.740 ;
        RECT 2148.270 15.200 2148.590 15.260 ;
        RECT 2118.000 15.060 2148.590 15.200 ;
        RECT 2148.270 15.000 2148.590 15.060 ;
      LAYER via ;
        RECT 848.800 15.680 849.060 15.940 ;
        RECT 2148.300 15.000 2148.560 15.260 ;
      LAYER met2 ;
        RECT 848.690 400.180 848.970 404.000 ;
        RECT 848.690 400.000 849.000 400.180 ;
        RECT 848.860 15.970 849.000 400.000 ;
        RECT 848.800 15.650 849.060 15.970 ;
        RECT 2148.300 14.970 2148.560 15.290 ;
        RECT 2148.360 2.400 2148.500 14.970 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 849.230 375.940 849.550 376.000 ;
        RECT 852.910 375.940 853.230 376.000 ;
        RECT 849.230 375.800 853.230 375.940 ;
        RECT 849.230 375.740 849.550 375.800 ;
        RECT 852.910 375.740 853.230 375.800 ;
        RECT 849.230 16.220 849.550 16.280 ;
        RECT 2166.210 16.220 2166.530 16.280 ;
        RECT 849.230 16.080 2166.530 16.220 ;
        RECT 849.230 16.020 849.550 16.080 ;
        RECT 2166.210 16.020 2166.530 16.080 ;
      LAYER via ;
        RECT 849.260 375.740 849.520 376.000 ;
        RECT 852.940 375.740 853.200 376.000 ;
        RECT 849.260 16.020 849.520 16.280 ;
        RECT 2166.240 16.020 2166.500 16.280 ;
      LAYER met2 ;
        RECT 854.210 400.250 854.490 404.000 ;
        RECT 853.000 400.110 854.490 400.250 ;
        RECT 853.000 376.030 853.140 400.110 ;
        RECT 854.210 400.000 854.490 400.110 ;
        RECT 849.260 375.710 849.520 376.030 ;
        RECT 852.940 375.710 853.200 376.030 ;
        RECT 849.320 16.310 849.460 375.710 ;
        RECT 849.260 15.990 849.520 16.310 ;
        RECT 2166.240 15.990 2166.500 16.310 ;
        RECT 2166.300 2.400 2166.440 15.990 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 855.670 375.940 855.990 376.000 ;
        RECT 857.970 375.940 858.290 376.000 ;
        RECT 855.670 375.800 858.290 375.940 ;
        RECT 855.670 375.740 855.990 375.800 ;
        RECT 857.970 375.740 858.290 375.800 ;
        RECT 855.670 16.560 855.990 16.620 ;
        RECT 2183.690 16.560 2184.010 16.620 ;
        RECT 855.670 16.420 2184.010 16.560 ;
        RECT 855.670 16.360 855.990 16.420 ;
        RECT 2183.690 16.360 2184.010 16.420 ;
      LAYER via ;
        RECT 855.700 375.740 855.960 376.000 ;
        RECT 858.000 375.740 858.260 376.000 ;
        RECT 855.700 16.360 855.960 16.620 ;
        RECT 2183.720 16.360 2183.980 16.620 ;
      LAYER met2 ;
        RECT 859.270 400.250 859.550 404.000 ;
        RECT 858.060 400.110 859.550 400.250 ;
        RECT 858.060 376.030 858.200 400.110 ;
        RECT 859.270 400.000 859.550 400.110 ;
        RECT 855.700 375.710 855.960 376.030 ;
        RECT 858.000 375.710 858.260 376.030 ;
        RECT 855.760 16.650 855.900 375.710 ;
        RECT 855.700 16.330 855.960 16.650 ;
        RECT 2183.720 16.330 2183.980 16.650 ;
        RECT 2183.780 2.400 2183.920 16.330 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 862.570 375.940 862.890 376.000 ;
        RECT 864.410 375.940 864.730 376.000 ;
        RECT 862.570 375.800 864.730 375.940 ;
        RECT 862.570 375.740 862.890 375.800 ;
        RECT 864.410 375.740 864.730 375.800 ;
        RECT 862.570 16.900 862.890 16.960 ;
        RECT 2201.170 16.900 2201.490 16.960 ;
        RECT 862.570 16.760 2201.490 16.900 ;
        RECT 862.570 16.700 862.890 16.760 ;
        RECT 2201.170 16.700 2201.490 16.760 ;
      LAYER via ;
        RECT 862.600 375.740 862.860 376.000 ;
        RECT 864.440 375.740 864.700 376.000 ;
        RECT 862.600 16.700 862.860 16.960 ;
        RECT 2201.200 16.700 2201.460 16.960 ;
      LAYER met2 ;
        RECT 864.790 400.250 865.070 404.000 ;
        RECT 864.500 400.110 865.070 400.250 ;
        RECT 864.500 376.030 864.640 400.110 ;
        RECT 864.790 400.000 865.070 400.110 ;
        RECT 862.600 375.710 862.860 376.030 ;
        RECT 864.440 375.710 864.700 376.030 ;
        RECT 862.660 16.990 862.800 375.710 ;
        RECT 862.600 16.670 862.860 16.990 ;
        RECT 2201.200 16.670 2201.460 16.990 ;
        RECT 2201.260 8.570 2201.400 16.670 ;
        RECT 2201.260 8.430 2201.860 8.570 ;
        RECT 2201.720 2.400 2201.860 8.430 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.930 20.640 870.250 20.700 ;
        RECT 2219.110 20.640 2219.430 20.700 ;
        RECT 869.930 20.500 2219.430 20.640 ;
        RECT 869.930 20.440 870.250 20.500 ;
        RECT 2219.110 20.440 2219.430 20.500 ;
      LAYER via ;
        RECT 869.960 20.440 870.220 20.700 ;
        RECT 2219.140 20.440 2219.400 20.700 ;
      LAYER met2 ;
        RECT 870.310 400.250 870.590 404.000 ;
        RECT 870.020 400.110 870.590 400.250 ;
        RECT 870.020 20.730 870.160 400.110 ;
        RECT 870.310 400.000 870.590 400.110 ;
        RECT 869.960 20.410 870.220 20.730 ;
        RECT 2219.140 20.410 2219.400 20.730 ;
        RECT 2219.200 2.400 2219.340 20.410 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.070 400.250 436.350 404.000 ;
        RECT 434.860 400.110 436.350 400.250 ;
        RECT 434.860 17.525 435.000 400.110 ;
        RECT 436.070 400.000 436.350 400.110 ;
        RECT 434.790 17.155 435.070 17.525 ;
        RECT 783.010 17.155 783.290 17.525 ;
        RECT 783.080 2.400 783.220 17.155 ;
        RECT 782.870 -4.800 783.430 2.400 ;
      LAYER via2 ;
        RECT 434.790 17.200 435.070 17.480 ;
        RECT 783.010 17.200 783.290 17.480 ;
      LAYER met3 ;
        RECT 434.765 17.490 435.095 17.505 ;
        RECT 782.985 17.490 783.315 17.505 ;
        RECT 434.765 17.190 783.315 17.490 ;
        RECT 434.765 17.175 435.095 17.190 ;
        RECT 782.985 17.175 783.315 17.190 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.470 376.280 869.790 376.340 ;
        RECT 874.070 376.280 874.390 376.340 ;
        RECT 869.470 376.140 874.390 376.280 ;
        RECT 869.470 376.080 869.790 376.140 ;
        RECT 874.070 376.080 874.390 376.140 ;
        RECT 869.470 20.300 869.790 20.360 ;
        RECT 2237.050 20.300 2237.370 20.360 ;
        RECT 869.470 20.160 2237.370 20.300 ;
        RECT 869.470 20.100 869.790 20.160 ;
        RECT 2237.050 20.100 2237.370 20.160 ;
      LAYER via ;
        RECT 869.500 376.080 869.760 376.340 ;
        RECT 874.100 376.080 874.360 376.340 ;
        RECT 869.500 20.100 869.760 20.360 ;
        RECT 2237.080 20.100 2237.340 20.360 ;
      LAYER met2 ;
        RECT 875.370 400.250 875.650 404.000 ;
        RECT 874.160 400.110 875.650 400.250 ;
        RECT 874.160 376.370 874.300 400.110 ;
        RECT 875.370 400.000 875.650 400.110 ;
        RECT 869.500 376.050 869.760 376.370 ;
        RECT 874.100 376.050 874.360 376.370 ;
        RECT 869.560 20.390 869.700 376.050 ;
        RECT 869.500 20.070 869.760 20.390 ;
        RECT 2237.080 20.070 2237.340 20.390 ;
        RECT 2237.140 2.400 2237.280 20.070 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.370 375.940 876.690 376.000 ;
        RECT 879.590 375.940 879.910 376.000 ;
        RECT 876.370 375.800 879.910 375.940 ;
        RECT 876.370 375.740 876.690 375.800 ;
        RECT 879.590 375.740 879.910 375.800 ;
        RECT 876.370 19.960 876.690 20.020 ;
        RECT 2254.530 19.960 2254.850 20.020 ;
        RECT 876.370 19.820 2254.850 19.960 ;
        RECT 876.370 19.760 876.690 19.820 ;
        RECT 2254.530 19.760 2254.850 19.820 ;
      LAYER via ;
        RECT 876.400 375.740 876.660 376.000 ;
        RECT 879.620 375.740 879.880 376.000 ;
        RECT 876.400 19.760 876.660 20.020 ;
        RECT 2254.560 19.760 2254.820 20.020 ;
      LAYER met2 ;
        RECT 880.890 400.250 881.170 404.000 ;
        RECT 879.680 400.110 881.170 400.250 ;
        RECT 879.680 376.030 879.820 400.110 ;
        RECT 880.890 400.000 881.170 400.110 ;
        RECT 876.400 375.710 876.660 376.030 ;
        RECT 879.620 375.710 879.880 376.030 ;
        RECT 876.460 20.050 876.600 375.710 ;
        RECT 876.400 19.730 876.660 20.050 ;
        RECT 2254.560 19.730 2254.820 20.050 ;
        RECT 2254.620 2.400 2254.760 19.730 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.270 387.500 883.590 387.560 ;
        RECT 886.490 387.500 886.810 387.560 ;
        RECT 883.270 387.360 886.810 387.500 ;
        RECT 883.270 387.300 883.590 387.360 ;
        RECT 886.490 387.300 886.810 387.360 ;
        RECT 883.270 19.620 883.590 19.680 ;
        RECT 2272.470 19.620 2272.790 19.680 ;
        RECT 883.270 19.480 2272.790 19.620 ;
        RECT 883.270 19.420 883.590 19.480 ;
        RECT 2272.470 19.420 2272.790 19.480 ;
      LAYER via ;
        RECT 883.300 387.300 883.560 387.560 ;
        RECT 886.520 387.300 886.780 387.560 ;
        RECT 883.300 19.420 883.560 19.680 ;
        RECT 2272.500 19.420 2272.760 19.680 ;
      LAYER met2 ;
        RECT 886.410 400.180 886.690 404.000 ;
        RECT 886.410 400.000 886.720 400.180 ;
        RECT 886.580 387.590 886.720 400.000 ;
        RECT 883.300 387.270 883.560 387.590 ;
        RECT 886.520 387.270 886.780 387.590 ;
        RECT 883.360 19.710 883.500 387.270 ;
        RECT 883.300 19.390 883.560 19.710 ;
        RECT 2272.500 19.390 2272.760 19.710 ;
        RECT 2272.560 2.400 2272.700 19.390 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.170 19.280 890.490 19.340 ;
        RECT 2290.410 19.280 2290.730 19.340 ;
        RECT 890.170 19.140 2290.730 19.280 ;
        RECT 890.170 19.080 890.490 19.140 ;
        RECT 2290.410 19.080 2290.730 19.140 ;
      LAYER via ;
        RECT 890.200 19.080 890.460 19.340 ;
        RECT 2290.440 19.080 2290.700 19.340 ;
      LAYER met2 ;
        RECT 891.470 400.250 891.750 404.000 ;
        RECT 890.260 400.110 891.750 400.250 ;
        RECT 890.260 19.370 890.400 400.110 ;
        RECT 891.470 400.000 891.750 400.110 ;
        RECT 890.200 19.050 890.460 19.370 ;
        RECT 2290.440 19.050 2290.700 19.370 ;
        RECT 2290.500 2.400 2290.640 19.050 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.530 18.940 897.850 19.000 ;
        RECT 2307.890 18.940 2308.210 19.000 ;
        RECT 897.530 18.800 2308.210 18.940 ;
        RECT 897.530 18.740 897.850 18.800 ;
        RECT 2307.890 18.740 2308.210 18.800 ;
      LAYER via ;
        RECT 897.560 18.740 897.820 19.000 ;
        RECT 2307.920 18.740 2308.180 19.000 ;
      LAYER met2 ;
        RECT 896.990 400.250 897.270 404.000 ;
        RECT 896.990 400.110 897.760 400.250 ;
        RECT 896.990 400.000 897.270 400.110 ;
        RECT 897.620 19.030 897.760 400.110 ;
        RECT 897.560 18.710 897.820 19.030 ;
        RECT 2307.920 18.710 2308.180 19.030 ;
        RECT 2307.980 2.400 2308.120 18.710 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.070 376.280 897.390 376.340 ;
        RECT 901.210 376.280 901.530 376.340 ;
        RECT 897.070 376.140 901.530 376.280 ;
        RECT 897.070 376.080 897.390 376.140 ;
        RECT 901.210 376.080 901.530 376.140 ;
        RECT 897.070 18.600 897.390 18.660 ;
        RECT 2325.830 18.600 2326.150 18.660 ;
        RECT 897.070 18.460 2326.150 18.600 ;
        RECT 897.070 18.400 897.390 18.460 ;
        RECT 2325.830 18.400 2326.150 18.460 ;
      LAYER via ;
        RECT 897.100 376.080 897.360 376.340 ;
        RECT 901.240 376.080 901.500 376.340 ;
        RECT 897.100 18.400 897.360 18.660 ;
        RECT 2325.860 18.400 2326.120 18.660 ;
      LAYER met2 ;
        RECT 902.050 400.250 902.330 404.000 ;
        RECT 901.300 400.110 902.330 400.250 ;
        RECT 901.300 376.370 901.440 400.110 ;
        RECT 902.050 400.000 902.330 400.110 ;
        RECT 897.100 376.050 897.360 376.370 ;
        RECT 901.240 376.050 901.500 376.370 ;
        RECT 897.160 18.690 897.300 376.050 ;
        RECT 897.100 18.370 897.360 18.690 ;
        RECT 2325.860 18.370 2326.120 18.690 ;
        RECT 2325.920 2.400 2326.060 18.370 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 903.970 375.940 904.290 376.000 ;
        RECT 906.270 375.940 906.590 376.000 ;
        RECT 903.970 375.800 906.590 375.940 ;
        RECT 903.970 375.740 904.290 375.800 ;
        RECT 906.270 375.740 906.590 375.800 ;
        RECT 903.970 18.260 904.290 18.320 ;
        RECT 2343.310 18.260 2343.630 18.320 ;
        RECT 903.970 18.120 2343.630 18.260 ;
        RECT 903.970 18.060 904.290 18.120 ;
        RECT 2343.310 18.060 2343.630 18.120 ;
      LAYER via ;
        RECT 904.000 375.740 904.260 376.000 ;
        RECT 906.300 375.740 906.560 376.000 ;
        RECT 904.000 18.060 904.260 18.320 ;
        RECT 2343.340 18.060 2343.600 18.320 ;
      LAYER met2 ;
        RECT 907.570 400.250 907.850 404.000 ;
        RECT 906.360 400.110 907.850 400.250 ;
        RECT 906.360 376.030 906.500 400.110 ;
        RECT 907.570 400.000 907.850 400.110 ;
        RECT 904.000 375.710 904.260 376.030 ;
        RECT 906.300 375.710 906.560 376.030 ;
        RECT 904.060 18.350 904.200 375.710 ;
        RECT 904.000 18.030 904.260 18.350 ;
        RECT 2343.340 18.030 2343.600 18.350 ;
        RECT 2343.400 2.400 2343.540 18.030 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 910.870 376.280 911.190 376.340 ;
        RECT 912.250 376.280 912.570 376.340 ;
        RECT 910.870 376.140 912.570 376.280 ;
        RECT 910.870 376.080 911.190 376.140 ;
        RECT 912.250 376.080 912.570 376.140 ;
        RECT 910.870 17.920 911.190 17.980 ;
        RECT 2361.250 17.920 2361.570 17.980 ;
        RECT 910.870 17.780 2361.570 17.920 ;
        RECT 910.870 17.720 911.190 17.780 ;
        RECT 2361.250 17.720 2361.570 17.780 ;
      LAYER via ;
        RECT 910.900 376.080 911.160 376.340 ;
        RECT 912.280 376.080 912.540 376.340 ;
        RECT 910.900 17.720 911.160 17.980 ;
        RECT 2361.280 17.720 2361.540 17.980 ;
      LAYER met2 ;
        RECT 913.090 400.250 913.370 404.000 ;
        RECT 912.340 400.110 913.370 400.250 ;
        RECT 912.340 376.370 912.480 400.110 ;
        RECT 913.090 400.000 913.370 400.110 ;
        RECT 910.900 376.050 911.160 376.370 ;
        RECT 912.280 376.050 912.540 376.370 ;
        RECT 910.960 18.010 911.100 376.050 ;
        RECT 910.900 17.690 911.160 18.010 ;
        RECT 2361.280 17.690 2361.540 18.010 ;
        RECT 2361.340 2.400 2361.480 17.690 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 917.770 17.580 918.090 17.640 ;
        RECT 917.770 17.440 2366.080 17.580 ;
        RECT 917.770 17.380 918.090 17.440 ;
        RECT 2365.940 17.240 2366.080 17.440 ;
        RECT 2378.730 17.240 2379.050 17.300 ;
        RECT 2365.940 17.100 2379.050 17.240 ;
        RECT 2378.730 17.040 2379.050 17.100 ;
      LAYER via ;
        RECT 917.800 17.380 918.060 17.640 ;
        RECT 2378.760 17.040 2379.020 17.300 ;
      LAYER met2 ;
        RECT 918.150 400.250 918.430 404.000 ;
        RECT 917.860 400.110 918.430 400.250 ;
        RECT 917.860 17.670 918.000 400.110 ;
        RECT 918.150 400.000 918.430 400.110 ;
        RECT 917.800 17.350 918.060 17.670 ;
        RECT 2378.760 17.010 2379.020 17.330 ;
        RECT 2378.820 2.400 2378.960 17.010 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.230 376.280 918.550 376.340 ;
        RECT 922.370 376.280 922.690 376.340 ;
        RECT 918.230 376.140 922.690 376.280 ;
        RECT 918.230 376.080 918.550 376.140 ;
        RECT 922.370 376.080 922.690 376.140 ;
        RECT 918.230 17.240 918.550 17.300 ;
        RECT 918.230 17.100 2352.970 17.240 ;
        RECT 918.230 17.040 918.550 17.100 ;
        RECT 2352.830 16.900 2352.970 17.100 ;
        RECT 2396.670 16.900 2396.990 16.960 ;
        RECT 2352.830 16.760 2396.990 16.900 ;
        RECT 2396.670 16.700 2396.990 16.760 ;
      LAYER via ;
        RECT 918.260 376.080 918.520 376.340 ;
        RECT 922.400 376.080 922.660 376.340 ;
        RECT 918.260 17.040 918.520 17.300 ;
        RECT 2396.700 16.700 2396.960 16.960 ;
      LAYER met2 ;
        RECT 923.670 400.250 923.950 404.000 ;
        RECT 922.460 400.110 923.950 400.250 ;
        RECT 922.460 376.370 922.600 400.110 ;
        RECT 923.670 400.000 923.950 400.110 ;
        RECT 918.260 376.050 918.520 376.370 ;
        RECT 922.400 376.050 922.660 376.370 ;
        RECT 918.320 17.330 918.460 376.050 ;
        RECT 918.260 17.010 918.520 17.330 ;
        RECT 2396.700 16.670 2396.960 16.990 ;
        RECT 2396.760 2.400 2396.900 16.670 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.130 386.480 442.450 386.540 ;
        RECT 443.510 386.480 443.830 386.540 ;
        RECT 442.130 386.340 443.830 386.480 ;
        RECT 442.130 386.280 442.450 386.340 ;
        RECT 443.510 386.280 443.830 386.340 ;
      LAYER via ;
        RECT 442.160 386.280 442.420 386.540 ;
        RECT 443.540 386.280 443.800 386.540 ;
      LAYER met2 ;
        RECT 441.590 400.250 441.870 404.000 ;
        RECT 441.590 400.110 442.360 400.250 ;
        RECT 441.590 400.000 441.870 400.110 ;
        RECT 442.220 386.570 442.360 400.110 ;
        RECT 442.160 386.250 442.420 386.570 ;
        RECT 443.540 386.250 443.800 386.570 ;
        RECT 443.600 16.845 443.740 386.250 ;
        RECT 443.530 16.475 443.810 16.845 ;
        RECT 800.490 16.475 800.770 16.845 ;
        RECT 800.560 2.400 800.700 16.475 ;
        RECT 800.350 -4.800 800.910 2.400 ;
      LAYER via2 ;
        RECT 443.530 16.520 443.810 16.800 ;
        RECT 800.490 16.520 800.770 16.800 ;
      LAYER met3 ;
        RECT 443.505 16.810 443.835 16.825 ;
        RECT 800.465 16.810 800.795 16.825 ;
        RECT 443.505 16.510 800.795 16.810 ;
        RECT 443.505 16.495 443.835 16.510 ;
        RECT 800.465 16.495 800.795 16.510 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1115.110 455.500 1115.430 455.560 ;
        RECT 2652.890 455.500 2653.210 455.560 ;
        RECT 1115.110 455.360 2653.210 455.500 ;
        RECT 1115.110 455.300 1115.430 455.360 ;
        RECT 2652.890 455.300 2653.210 455.360 ;
        RECT 2652.890 17.240 2653.210 17.300 ;
        RECT 2898.990 17.240 2899.310 17.300 ;
        RECT 2652.890 17.100 2899.310 17.240 ;
        RECT 2652.890 17.040 2653.210 17.100 ;
        RECT 2898.990 17.040 2899.310 17.100 ;
      LAYER via ;
        RECT 1115.140 455.300 1115.400 455.560 ;
        RECT 2652.920 455.300 2653.180 455.560 ;
        RECT 2652.920 17.040 2653.180 17.300 ;
        RECT 2899.020 17.040 2899.280 17.300 ;
      LAYER met2 ;
        RECT 1115.130 457.795 1115.410 458.165 ;
        RECT 1115.200 455.590 1115.340 457.795 ;
        RECT 1115.140 455.270 1115.400 455.590 ;
        RECT 2652.920 455.270 2653.180 455.590 ;
        RECT 2652.980 17.330 2653.120 455.270 ;
        RECT 2652.920 17.010 2653.180 17.330 ;
        RECT 2899.020 17.010 2899.280 17.330 ;
        RECT 2899.080 2.400 2899.220 17.010 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 1115.130 457.840 1115.410 458.120 ;
      LAYER met3 ;
        RECT 1096.000 459.880 1100.000 460.480 ;
        RECT 1098.790 458.130 1099.090 459.880 ;
        RECT 1115.105 458.130 1115.435 458.145 ;
        RECT 1098.790 457.830 1115.435 458.130 ;
        RECT 1115.105 457.815 1115.435 457.830 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 579.940 1117.730 580.000 ;
        RECT 1928.390 579.940 1928.710 580.000 ;
        RECT 1117.410 579.800 1928.710 579.940 ;
        RECT 1117.410 579.740 1117.730 579.800 ;
        RECT 1928.390 579.740 1928.710 579.800 ;
      LAYER via ;
        RECT 1117.440 579.740 1117.700 580.000 ;
        RECT 1928.420 579.740 1928.680 580.000 ;
      LAYER met2 ;
        RECT 1117.430 580.875 1117.710 581.245 ;
        RECT 1117.500 580.030 1117.640 580.875 ;
        RECT 1117.440 579.710 1117.700 580.030 ;
        RECT 1928.420 579.710 1928.680 580.030 ;
        RECT 1928.480 18.205 1928.620 579.710 ;
        RECT 1928.410 17.835 1928.690 18.205 ;
        RECT 2904.990 17.155 2905.270 17.525 ;
        RECT 2905.060 2.400 2905.200 17.155 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 1117.430 580.920 1117.710 581.200 ;
        RECT 1928.410 17.880 1928.690 18.160 ;
        RECT 2904.990 17.200 2905.270 17.480 ;
      LAYER met3 ;
        RECT 1117.405 581.210 1117.735 581.225 ;
        RECT 1097.870 580.910 1117.735 581.210 ;
        RECT 1097.870 580.160 1098.170 580.910 ;
        RECT 1117.405 580.895 1117.735 580.910 ;
        RECT 1096.000 579.560 1100.000 580.160 ;
        RECT 1928.385 18.170 1928.715 18.185 ;
        RECT 1928.385 17.870 1966.650 18.170 ;
        RECT 1928.385 17.855 1928.715 17.870 ;
        RECT 1966.350 17.490 1966.650 17.870 ;
        RECT 2904.965 17.490 2905.295 17.505 ;
        RECT 1966.350 17.190 2905.295 17.490 ;
        RECT 2904.965 17.175 2905.295 17.190 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.150 400.250 1079.430 404.000 ;
        RECT 1077.940 400.110 1079.430 400.250 ;
        RECT 1077.940 324.370 1078.080 400.110 ;
        RECT 1079.150 400.000 1079.430 400.110 ;
        RECT 1076.560 324.230 1078.080 324.370 ;
        RECT 1076.560 16.845 1076.700 324.230 ;
        RECT 1076.490 16.475 1076.770 16.845 ;
        RECT 2910.970 16.475 2911.250 16.845 ;
        RECT 2911.040 2.400 2911.180 16.475 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
      LAYER via2 ;
        RECT 1076.490 16.520 1076.770 16.800 ;
        RECT 2910.970 16.520 2911.250 16.800 ;
      LAYER met3 ;
        RECT 1076.465 16.810 1076.795 16.825 ;
        RECT 2910.945 16.810 2911.275 16.825 ;
        RECT 1076.465 16.510 2911.275 16.810 ;
        RECT 1076.465 16.495 1076.795 16.510 ;
        RECT 2910.945 16.495 2911.275 16.510 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 441.475 193.110 441.845 ;
        RECT 192.900 37.925 193.040 441.475 ;
        RECT 192.830 37.555 193.110 37.925 ;
        RECT 2916.950 37.555 2917.230 37.925 ;
        RECT 2917.020 2.400 2917.160 37.555 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
      LAYER via2 ;
        RECT 192.830 441.520 193.110 441.800 ;
        RECT 192.830 37.600 193.110 37.880 ;
        RECT 2916.950 37.600 2917.230 37.880 ;
      LAYER met3 ;
        RECT 200.000 442.880 204.000 443.480 ;
        RECT 192.805 441.810 193.135 441.825 ;
        RECT 200.870 441.810 201.170 442.880 ;
        RECT 192.805 441.510 201.170 441.810 ;
        RECT 192.805 441.495 193.135 441.510 ;
        RECT 192.805 37.890 193.135 37.905 ;
        RECT 2916.925 37.890 2917.255 37.905 ;
        RECT 192.805 37.590 2917.255 37.890 ;
        RECT 192.805 37.575 193.135 37.590 ;
        RECT 2916.925 37.575 2917.255 37.590 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
        RECT 188.970 1010.000 192.070 3529.150 ;
        RECT 368.970 1010.000 372.070 3529.150 ;
        RECT 548.970 1010.000 552.070 3529.150 ;
        RECT 728.970 1010.000 732.070 3529.150 ;
        RECT 908.970 1010.000 912.070 3529.150 ;
        RECT 1088.970 1010.000 1092.070 3529.150 ;
        RECT 221.040 410.640 222.640 987.760 ;
        RECT 374.640 410.640 376.240 987.760 ;
        RECT 528.240 410.640 529.840 987.760 ;
        RECT 681.840 410.640 683.440 987.760 ;
        RECT 835.440 410.640 837.040 987.760 ;
        RECT 989.040 410.640 990.640 987.760 ;
        RECT 188.970 -9.470 192.070 390.000 ;
        RECT 368.970 -9.470 372.070 390.000 ;
        RECT 548.970 -9.470 552.070 390.000 ;
        RECT 728.970 -9.470 732.070 390.000 ;
        RECT 908.970 -9.470 912.070 390.000 ;
        RECT 1088.970 -9.470 1092.070 390.000 ;
        RECT 1268.970 -9.470 1272.070 3529.150 ;
        RECT 1448.970 -9.470 1452.070 3529.150 ;
        RECT 1628.970 -9.470 1632.070 3529.150 ;
        RECT 1808.970 -9.470 1812.070 3529.150 ;
        RECT 1988.970 -9.470 1992.070 3529.150 ;
        RECT 2168.970 -9.470 2172.070 3529.150 ;
        RECT 2348.970 -9.470 2352.070 3529.150 ;
        RECT 2528.970 -9.470 2532.070 3529.150 ;
        RECT 2708.970 -9.470 2712.070 3529.150 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER via4 ;
        RECT -9.870 3523.010 -8.690 3524.190 ;
        RECT -8.270 3523.010 -7.090 3524.190 ;
        RECT -9.870 3521.410 -8.690 3522.590 ;
        RECT -8.270 3521.410 -7.090 3522.590 ;
        RECT -9.870 3436.090 -8.690 3437.270 ;
        RECT -8.270 3436.090 -7.090 3437.270 ;
        RECT -9.870 3434.490 -8.690 3435.670 ;
        RECT -8.270 3434.490 -7.090 3435.670 ;
        RECT -9.870 3256.090 -8.690 3257.270 ;
        RECT -8.270 3256.090 -7.090 3257.270 ;
        RECT -9.870 3254.490 -8.690 3255.670 ;
        RECT -8.270 3254.490 -7.090 3255.670 ;
        RECT -9.870 3076.090 -8.690 3077.270 ;
        RECT -8.270 3076.090 -7.090 3077.270 ;
        RECT -9.870 3074.490 -8.690 3075.670 ;
        RECT -8.270 3074.490 -7.090 3075.670 ;
        RECT -9.870 2896.090 -8.690 2897.270 ;
        RECT -8.270 2896.090 -7.090 2897.270 ;
        RECT -9.870 2894.490 -8.690 2895.670 ;
        RECT -8.270 2894.490 -7.090 2895.670 ;
        RECT -9.870 2716.090 -8.690 2717.270 ;
        RECT -8.270 2716.090 -7.090 2717.270 ;
        RECT -9.870 2714.490 -8.690 2715.670 ;
        RECT -8.270 2714.490 -7.090 2715.670 ;
        RECT -9.870 2536.090 -8.690 2537.270 ;
        RECT -8.270 2536.090 -7.090 2537.270 ;
        RECT -9.870 2534.490 -8.690 2535.670 ;
        RECT -8.270 2534.490 -7.090 2535.670 ;
        RECT -9.870 2356.090 -8.690 2357.270 ;
        RECT -8.270 2356.090 -7.090 2357.270 ;
        RECT -9.870 2354.490 -8.690 2355.670 ;
        RECT -8.270 2354.490 -7.090 2355.670 ;
        RECT -9.870 2176.090 -8.690 2177.270 ;
        RECT -8.270 2176.090 -7.090 2177.270 ;
        RECT -9.870 2174.490 -8.690 2175.670 ;
        RECT -8.270 2174.490 -7.090 2175.670 ;
        RECT -9.870 1996.090 -8.690 1997.270 ;
        RECT -8.270 1996.090 -7.090 1997.270 ;
        RECT -9.870 1994.490 -8.690 1995.670 ;
        RECT -8.270 1994.490 -7.090 1995.670 ;
        RECT -9.870 1816.090 -8.690 1817.270 ;
        RECT -8.270 1816.090 -7.090 1817.270 ;
        RECT -9.870 1814.490 -8.690 1815.670 ;
        RECT -8.270 1814.490 -7.090 1815.670 ;
        RECT -9.870 1636.090 -8.690 1637.270 ;
        RECT -8.270 1636.090 -7.090 1637.270 ;
        RECT -9.870 1634.490 -8.690 1635.670 ;
        RECT -8.270 1634.490 -7.090 1635.670 ;
        RECT -9.870 1456.090 -8.690 1457.270 ;
        RECT -8.270 1456.090 -7.090 1457.270 ;
        RECT -9.870 1454.490 -8.690 1455.670 ;
        RECT -8.270 1454.490 -7.090 1455.670 ;
        RECT -9.870 1276.090 -8.690 1277.270 ;
        RECT -8.270 1276.090 -7.090 1277.270 ;
        RECT -9.870 1274.490 -8.690 1275.670 ;
        RECT -8.270 1274.490 -7.090 1275.670 ;
        RECT -9.870 1096.090 -8.690 1097.270 ;
        RECT -8.270 1096.090 -7.090 1097.270 ;
        RECT -9.870 1094.490 -8.690 1095.670 ;
        RECT -8.270 1094.490 -7.090 1095.670 ;
        RECT -9.870 916.090 -8.690 917.270 ;
        RECT -8.270 916.090 -7.090 917.270 ;
        RECT -9.870 914.490 -8.690 915.670 ;
        RECT -8.270 914.490 -7.090 915.670 ;
        RECT -9.870 736.090 -8.690 737.270 ;
        RECT -8.270 736.090 -7.090 737.270 ;
        RECT -9.870 734.490 -8.690 735.670 ;
        RECT -8.270 734.490 -7.090 735.670 ;
        RECT -9.870 556.090 -8.690 557.270 ;
        RECT -8.270 556.090 -7.090 557.270 ;
        RECT -9.870 554.490 -8.690 555.670 ;
        RECT -8.270 554.490 -7.090 555.670 ;
        RECT -9.870 376.090 -8.690 377.270 ;
        RECT -8.270 376.090 -7.090 377.270 ;
        RECT -9.870 374.490 -8.690 375.670 ;
        RECT -8.270 374.490 -7.090 375.670 ;
        RECT -9.870 196.090 -8.690 197.270 ;
        RECT -8.270 196.090 -7.090 197.270 ;
        RECT -9.870 194.490 -8.690 195.670 ;
        RECT -8.270 194.490 -7.090 195.670 ;
        RECT -9.870 16.090 -8.690 17.270 ;
        RECT -8.270 16.090 -7.090 17.270 ;
        RECT -9.870 14.490 -8.690 15.670 ;
        RECT -8.270 14.490 -7.090 15.670 ;
        RECT -9.870 -2.910 -8.690 -1.730 ;
        RECT -8.270 -2.910 -7.090 -1.730 ;
        RECT -9.870 -4.510 -8.690 -3.330 ;
        RECT -8.270 -4.510 -7.090 -3.330 ;
        RECT 9.130 3523.010 10.310 3524.190 ;
        RECT 10.730 3523.010 11.910 3524.190 ;
        RECT 9.130 3521.410 10.310 3522.590 ;
        RECT 10.730 3521.410 11.910 3522.590 ;
        RECT 9.130 3436.090 10.310 3437.270 ;
        RECT 10.730 3436.090 11.910 3437.270 ;
        RECT 9.130 3434.490 10.310 3435.670 ;
        RECT 10.730 3434.490 11.910 3435.670 ;
        RECT 9.130 3256.090 10.310 3257.270 ;
        RECT 10.730 3256.090 11.910 3257.270 ;
        RECT 9.130 3254.490 10.310 3255.670 ;
        RECT 10.730 3254.490 11.910 3255.670 ;
        RECT 9.130 3076.090 10.310 3077.270 ;
        RECT 10.730 3076.090 11.910 3077.270 ;
        RECT 9.130 3074.490 10.310 3075.670 ;
        RECT 10.730 3074.490 11.910 3075.670 ;
        RECT 9.130 2896.090 10.310 2897.270 ;
        RECT 10.730 2896.090 11.910 2897.270 ;
        RECT 9.130 2894.490 10.310 2895.670 ;
        RECT 10.730 2894.490 11.910 2895.670 ;
        RECT 9.130 2716.090 10.310 2717.270 ;
        RECT 10.730 2716.090 11.910 2717.270 ;
        RECT 9.130 2714.490 10.310 2715.670 ;
        RECT 10.730 2714.490 11.910 2715.670 ;
        RECT 9.130 2536.090 10.310 2537.270 ;
        RECT 10.730 2536.090 11.910 2537.270 ;
        RECT 9.130 2534.490 10.310 2535.670 ;
        RECT 10.730 2534.490 11.910 2535.670 ;
        RECT 9.130 2356.090 10.310 2357.270 ;
        RECT 10.730 2356.090 11.910 2357.270 ;
        RECT 9.130 2354.490 10.310 2355.670 ;
        RECT 10.730 2354.490 11.910 2355.670 ;
        RECT 9.130 2176.090 10.310 2177.270 ;
        RECT 10.730 2176.090 11.910 2177.270 ;
        RECT 9.130 2174.490 10.310 2175.670 ;
        RECT 10.730 2174.490 11.910 2175.670 ;
        RECT 9.130 1996.090 10.310 1997.270 ;
        RECT 10.730 1996.090 11.910 1997.270 ;
        RECT 9.130 1994.490 10.310 1995.670 ;
        RECT 10.730 1994.490 11.910 1995.670 ;
        RECT 9.130 1816.090 10.310 1817.270 ;
        RECT 10.730 1816.090 11.910 1817.270 ;
        RECT 9.130 1814.490 10.310 1815.670 ;
        RECT 10.730 1814.490 11.910 1815.670 ;
        RECT 9.130 1636.090 10.310 1637.270 ;
        RECT 10.730 1636.090 11.910 1637.270 ;
        RECT 9.130 1634.490 10.310 1635.670 ;
        RECT 10.730 1634.490 11.910 1635.670 ;
        RECT 9.130 1456.090 10.310 1457.270 ;
        RECT 10.730 1456.090 11.910 1457.270 ;
        RECT 9.130 1454.490 10.310 1455.670 ;
        RECT 10.730 1454.490 11.910 1455.670 ;
        RECT 9.130 1276.090 10.310 1277.270 ;
        RECT 10.730 1276.090 11.910 1277.270 ;
        RECT 9.130 1274.490 10.310 1275.670 ;
        RECT 10.730 1274.490 11.910 1275.670 ;
        RECT 9.130 1096.090 10.310 1097.270 ;
        RECT 10.730 1096.090 11.910 1097.270 ;
        RECT 9.130 1094.490 10.310 1095.670 ;
        RECT 10.730 1094.490 11.910 1095.670 ;
        RECT 189.130 3523.010 190.310 3524.190 ;
        RECT 190.730 3523.010 191.910 3524.190 ;
        RECT 189.130 3521.410 190.310 3522.590 ;
        RECT 190.730 3521.410 191.910 3522.590 ;
        RECT 189.130 3436.090 190.310 3437.270 ;
        RECT 190.730 3436.090 191.910 3437.270 ;
        RECT 189.130 3434.490 190.310 3435.670 ;
        RECT 190.730 3434.490 191.910 3435.670 ;
        RECT 189.130 3256.090 190.310 3257.270 ;
        RECT 190.730 3256.090 191.910 3257.270 ;
        RECT 189.130 3254.490 190.310 3255.670 ;
        RECT 190.730 3254.490 191.910 3255.670 ;
        RECT 189.130 3076.090 190.310 3077.270 ;
        RECT 190.730 3076.090 191.910 3077.270 ;
        RECT 189.130 3074.490 190.310 3075.670 ;
        RECT 190.730 3074.490 191.910 3075.670 ;
        RECT 189.130 2896.090 190.310 2897.270 ;
        RECT 190.730 2896.090 191.910 2897.270 ;
        RECT 189.130 2894.490 190.310 2895.670 ;
        RECT 190.730 2894.490 191.910 2895.670 ;
        RECT 189.130 2716.090 190.310 2717.270 ;
        RECT 190.730 2716.090 191.910 2717.270 ;
        RECT 189.130 2714.490 190.310 2715.670 ;
        RECT 190.730 2714.490 191.910 2715.670 ;
        RECT 189.130 2536.090 190.310 2537.270 ;
        RECT 190.730 2536.090 191.910 2537.270 ;
        RECT 189.130 2534.490 190.310 2535.670 ;
        RECT 190.730 2534.490 191.910 2535.670 ;
        RECT 189.130 2356.090 190.310 2357.270 ;
        RECT 190.730 2356.090 191.910 2357.270 ;
        RECT 189.130 2354.490 190.310 2355.670 ;
        RECT 190.730 2354.490 191.910 2355.670 ;
        RECT 189.130 2176.090 190.310 2177.270 ;
        RECT 190.730 2176.090 191.910 2177.270 ;
        RECT 189.130 2174.490 190.310 2175.670 ;
        RECT 190.730 2174.490 191.910 2175.670 ;
        RECT 189.130 1996.090 190.310 1997.270 ;
        RECT 190.730 1996.090 191.910 1997.270 ;
        RECT 189.130 1994.490 190.310 1995.670 ;
        RECT 190.730 1994.490 191.910 1995.670 ;
        RECT 189.130 1816.090 190.310 1817.270 ;
        RECT 190.730 1816.090 191.910 1817.270 ;
        RECT 189.130 1814.490 190.310 1815.670 ;
        RECT 190.730 1814.490 191.910 1815.670 ;
        RECT 189.130 1636.090 190.310 1637.270 ;
        RECT 190.730 1636.090 191.910 1637.270 ;
        RECT 189.130 1634.490 190.310 1635.670 ;
        RECT 190.730 1634.490 191.910 1635.670 ;
        RECT 189.130 1456.090 190.310 1457.270 ;
        RECT 190.730 1456.090 191.910 1457.270 ;
        RECT 189.130 1454.490 190.310 1455.670 ;
        RECT 190.730 1454.490 191.910 1455.670 ;
        RECT 189.130 1276.090 190.310 1277.270 ;
        RECT 190.730 1276.090 191.910 1277.270 ;
        RECT 189.130 1274.490 190.310 1275.670 ;
        RECT 190.730 1274.490 191.910 1275.670 ;
        RECT 189.130 1096.090 190.310 1097.270 ;
        RECT 190.730 1096.090 191.910 1097.270 ;
        RECT 189.130 1094.490 190.310 1095.670 ;
        RECT 190.730 1094.490 191.910 1095.670 ;
        RECT 369.130 3523.010 370.310 3524.190 ;
        RECT 370.730 3523.010 371.910 3524.190 ;
        RECT 369.130 3521.410 370.310 3522.590 ;
        RECT 370.730 3521.410 371.910 3522.590 ;
        RECT 369.130 3436.090 370.310 3437.270 ;
        RECT 370.730 3436.090 371.910 3437.270 ;
        RECT 369.130 3434.490 370.310 3435.670 ;
        RECT 370.730 3434.490 371.910 3435.670 ;
        RECT 369.130 3256.090 370.310 3257.270 ;
        RECT 370.730 3256.090 371.910 3257.270 ;
        RECT 369.130 3254.490 370.310 3255.670 ;
        RECT 370.730 3254.490 371.910 3255.670 ;
        RECT 369.130 3076.090 370.310 3077.270 ;
        RECT 370.730 3076.090 371.910 3077.270 ;
        RECT 369.130 3074.490 370.310 3075.670 ;
        RECT 370.730 3074.490 371.910 3075.670 ;
        RECT 369.130 2896.090 370.310 2897.270 ;
        RECT 370.730 2896.090 371.910 2897.270 ;
        RECT 369.130 2894.490 370.310 2895.670 ;
        RECT 370.730 2894.490 371.910 2895.670 ;
        RECT 369.130 2716.090 370.310 2717.270 ;
        RECT 370.730 2716.090 371.910 2717.270 ;
        RECT 369.130 2714.490 370.310 2715.670 ;
        RECT 370.730 2714.490 371.910 2715.670 ;
        RECT 369.130 2536.090 370.310 2537.270 ;
        RECT 370.730 2536.090 371.910 2537.270 ;
        RECT 369.130 2534.490 370.310 2535.670 ;
        RECT 370.730 2534.490 371.910 2535.670 ;
        RECT 369.130 2356.090 370.310 2357.270 ;
        RECT 370.730 2356.090 371.910 2357.270 ;
        RECT 369.130 2354.490 370.310 2355.670 ;
        RECT 370.730 2354.490 371.910 2355.670 ;
        RECT 369.130 2176.090 370.310 2177.270 ;
        RECT 370.730 2176.090 371.910 2177.270 ;
        RECT 369.130 2174.490 370.310 2175.670 ;
        RECT 370.730 2174.490 371.910 2175.670 ;
        RECT 369.130 1996.090 370.310 1997.270 ;
        RECT 370.730 1996.090 371.910 1997.270 ;
        RECT 369.130 1994.490 370.310 1995.670 ;
        RECT 370.730 1994.490 371.910 1995.670 ;
        RECT 369.130 1816.090 370.310 1817.270 ;
        RECT 370.730 1816.090 371.910 1817.270 ;
        RECT 369.130 1814.490 370.310 1815.670 ;
        RECT 370.730 1814.490 371.910 1815.670 ;
        RECT 369.130 1636.090 370.310 1637.270 ;
        RECT 370.730 1636.090 371.910 1637.270 ;
        RECT 369.130 1634.490 370.310 1635.670 ;
        RECT 370.730 1634.490 371.910 1635.670 ;
        RECT 369.130 1456.090 370.310 1457.270 ;
        RECT 370.730 1456.090 371.910 1457.270 ;
        RECT 369.130 1454.490 370.310 1455.670 ;
        RECT 370.730 1454.490 371.910 1455.670 ;
        RECT 369.130 1276.090 370.310 1277.270 ;
        RECT 370.730 1276.090 371.910 1277.270 ;
        RECT 369.130 1274.490 370.310 1275.670 ;
        RECT 370.730 1274.490 371.910 1275.670 ;
        RECT 369.130 1096.090 370.310 1097.270 ;
        RECT 370.730 1096.090 371.910 1097.270 ;
        RECT 369.130 1094.490 370.310 1095.670 ;
        RECT 370.730 1094.490 371.910 1095.670 ;
        RECT 549.130 3523.010 550.310 3524.190 ;
        RECT 550.730 3523.010 551.910 3524.190 ;
        RECT 549.130 3521.410 550.310 3522.590 ;
        RECT 550.730 3521.410 551.910 3522.590 ;
        RECT 549.130 3436.090 550.310 3437.270 ;
        RECT 550.730 3436.090 551.910 3437.270 ;
        RECT 549.130 3434.490 550.310 3435.670 ;
        RECT 550.730 3434.490 551.910 3435.670 ;
        RECT 549.130 3256.090 550.310 3257.270 ;
        RECT 550.730 3256.090 551.910 3257.270 ;
        RECT 549.130 3254.490 550.310 3255.670 ;
        RECT 550.730 3254.490 551.910 3255.670 ;
        RECT 549.130 3076.090 550.310 3077.270 ;
        RECT 550.730 3076.090 551.910 3077.270 ;
        RECT 549.130 3074.490 550.310 3075.670 ;
        RECT 550.730 3074.490 551.910 3075.670 ;
        RECT 549.130 2896.090 550.310 2897.270 ;
        RECT 550.730 2896.090 551.910 2897.270 ;
        RECT 549.130 2894.490 550.310 2895.670 ;
        RECT 550.730 2894.490 551.910 2895.670 ;
        RECT 549.130 2716.090 550.310 2717.270 ;
        RECT 550.730 2716.090 551.910 2717.270 ;
        RECT 549.130 2714.490 550.310 2715.670 ;
        RECT 550.730 2714.490 551.910 2715.670 ;
        RECT 549.130 2536.090 550.310 2537.270 ;
        RECT 550.730 2536.090 551.910 2537.270 ;
        RECT 549.130 2534.490 550.310 2535.670 ;
        RECT 550.730 2534.490 551.910 2535.670 ;
        RECT 549.130 2356.090 550.310 2357.270 ;
        RECT 550.730 2356.090 551.910 2357.270 ;
        RECT 549.130 2354.490 550.310 2355.670 ;
        RECT 550.730 2354.490 551.910 2355.670 ;
        RECT 549.130 2176.090 550.310 2177.270 ;
        RECT 550.730 2176.090 551.910 2177.270 ;
        RECT 549.130 2174.490 550.310 2175.670 ;
        RECT 550.730 2174.490 551.910 2175.670 ;
        RECT 549.130 1996.090 550.310 1997.270 ;
        RECT 550.730 1996.090 551.910 1997.270 ;
        RECT 549.130 1994.490 550.310 1995.670 ;
        RECT 550.730 1994.490 551.910 1995.670 ;
        RECT 549.130 1816.090 550.310 1817.270 ;
        RECT 550.730 1816.090 551.910 1817.270 ;
        RECT 549.130 1814.490 550.310 1815.670 ;
        RECT 550.730 1814.490 551.910 1815.670 ;
        RECT 549.130 1636.090 550.310 1637.270 ;
        RECT 550.730 1636.090 551.910 1637.270 ;
        RECT 549.130 1634.490 550.310 1635.670 ;
        RECT 550.730 1634.490 551.910 1635.670 ;
        RECT 549.130 1456.090 550.310 1457.270 ;
        RECT 550.730 1456.090 551.910 1457.270 ;
        RECT 549.130 1454.490 550.310 1455.670 ;
        RECT 550.730 1454.490 551.910 1455.670 ;
        RECT 549.130 1276.090 550.310 1277.270 ;
        RECT 550.730 1276.090 551.910 1277.270 ;
        RECT 549.130 1274.490 550.310 1275.670 ;
        RECT 550.730 1274.490 551.910 1275.670 ;
        RECT 549.130 1096.090 550.310 1097.270 ;
        RECT 550.730 1096.090 551.910 1097.270 ;
        RECT 549.130 1094.490 550.310 1095.670 ;
        RECT 550.730 1094.490 551.910 1095.670 ;
        RECT 729.130 3523.010 730.310 3524.190 ;
        RECT 730.730 3523.010 731.910 3524.190 ;
        RECT 729.130 3521.410 730.310 3522.590 ;
        RECT 730.730 3521.410 731.910 3522.590 ;
        RECT 729.130 3436.090 730.310 3437.270 ;
        RECT 730.730 3436.090 731.910 3437.270 ;
        RECT 729.130 3434.490 730.310 3435.670 ;
        RECT 730.730 3434.490 731.910 3435.670 ;
        RECT 729.130 3256.090 730.310 3257.270 ;
        RECT 730.730 3256.090 731.910 3257.270 ;
        RECT 729.130 3254.490 730.310 3255.670 ;
        RECT 730.730 3254.490 731.910 3255.670 ;
        RECT 729.130 3076.090 730.310 3077.270 ;
        RECT 730.730 3076.090 731.910 3077.270 ;
        RECT 729.130 3074.490 730.310 3075.670 ;
        RECT 730.730 3074.490 731.910 3075.670 ;
        RECT 729.130 2896.090 730.310 2897.270 ;
        RECT 730.730 2896.090 731.910 2897.270 ;
        RECT 729.130 2894.490 730.310 2895.670 ;
        RECT 730.730 2894.490 731.910 2895.670 ;
        RECT 729.130 2716.090 730.310 2717.270 ;
        RECT 730.730 2716.090 731.910 2717.270 ;
        RECT 729.130 2714.490 730.310 2715.670 ;
        RECT 730.730 2714.490 731.910 2715.670 ;
        RECT 729.130 2536.090 730.310 2537.270 ;
        RECT 730.730 2536.090 731.910 2537.270 ;
        RECT 729.130 2534.490 730.310 2535.670 ;
        RECT 730.730 2534.490 731.910 2535.670 ;
        RECT 729.130 2356.090 730.310 2357.270 ;
        RECT 730.730 2356.090 731.910 2357.270 ;
        RECT 729.130 2354.490 730.310 2355.670 ;
        RECT 730.730 2354.490 731.910 2355.670 ;
        RECT 729.130 2176.090 730.310 2177.270 ;
        RECT 730.730 2176.090 731.910 2177.270 ;
        RECT 729.130 2174.490 730.310 2175.670 ;
        RECT 730.730 2174.490 731.910 2175.670 ;
        RECT 729.130 1996.090 730.310 1997.270 ;
        RECT 730.730 1996.090 731.910 1997.270 ;
        RECT 729.130 1994.490 730.310 1995.670 ;
        RECT 730.730 1994.490 731.910 1995.670 ;
        RECT 729.130 1816.090 730.310 1817.270 ;
        RECT 730.730 1816.090 731.910 1817.270 ;
        RECT 729.130 1814.490 730.310 1815.670 ;
        RECT 730.730 1814.490 731.910 1815.670 ;
        RECT 729.130 1636.090 730.310 1637.270 ;
        RECT 730.730 1636.090 731.910 1637.270 ;
        RECT 729.130 1634.490 730.310 1635.670 ;
        RECT 730.730 1634.490 731.910 1635.670 ;
        RECT 729.130 1456.090 730.310 1457.270 ;
        RECT 730.730 1456.090 731.910 1457.270 ;
        RECT 729.130 1454.490 730.310 1455.670 ;
        RECT 730.730 1454.490 731.910 1455.670 ;
        RECT 729.130 1276.090 730.310 1277.270 ;
        RECT 730.730 1276.090 731.910 1277.270 ;
        RECT 729.130 1274.490 730.310 1275.670 ;
        RECT 730.730 1274.490 731.910 1275.670 ;
        RECT 729.130 1096.090 730.310 1097.270 ;
        RECT 730.730 1096.090 731.910 1097.270 ;
        RECT 729.130 1094.490 730.310 1095.670 ;
        RECT 730.730 1094.490 731.910 1095.670 ;
        RECT 909.130 3523.010 910.310 3524.190 ;
        RECT 910.730 3523.010 911.910 3524.190 ;
        RECT 909.130 3521.410 910.310 3522.590 ;
        RECT 910.730 3521.410 911.910 3522.590 ;
        RECT 909.130 3436.090 910.310 3437.270 ;
        RECT 910.730 3436.090 911.910 3437.270 ;
        RECT 909.130 3434.490 910.310 3435.670 ;
        RECT 910.730 3434.490 911.910 3435.670 ;
        RECT 909.130 3256.090 910.310 3257.270 ;
        RECT 910.730 3256.090 911.910 3257.270 ;
        RECT 909.130 3254.490 910.310 3255.670 ;
        RECT 910.730 3254.490 911.910 3255.670 ;
        RECT 909.130 3076.090 910.310 3077.270 ;
        RECT 910.730 3076.090 911.910 3077.270 ;
        RECT 909.130 3074.490 910.310 3075.670 ;
        RECT 910.730 3074.490 911.910 3075.670 ;
        RECT 909.130 2896.090 910.310 2897.270 ;
        RECT 910.730 2896.090 911.910 2897.270 ;
        RECT 909.130 2894.490 910.310 2895.670 ;
        RECT 910.730 2894.490 911.910 2895.670 ;
        RECT 909.130 2716.090 910.310 2717.270 ;
        RECT 910.730 2716.090 911.910 2717.270 ;
        RECT 909.130 2714.490 910.310 2715.670 ;
        RECT 910.730 2714.490 911.910 2715.670 ;
        RECT 909.130 2536.090 910.310 2537.270 ;
        RECT 910.730 2536.090 911.910 2537.270 ;
        RECT 909.130 2534.490 910.310 2535.670 ;
        RECT 910.730 2534.490 911.910 2535.670 ;
        RECT 909.130 2356.090 910.310 2357.270 ;
        RECT 910.730 2356.090 911.910 2357.270 ;
        RECT 909.130 2354.490 910.310 2355.670 ;
        RECT 910.730 2354.490 911.910 2355.670 ;
        RECT 909.130 2176.090 910.310 2177.270 ;
        RECT 910.730 2176.090 911.910 2177.270 ;
        RECT 909.130 2174.490 910.310 2175.670 ;
        RECT 910.730 2174.490 911.910 2175.670 ;
        RECT 909.130 1996.090 910.310 1997.270 ;
        RECT 910.730 1996.090 911.910 1997.270 ;
        RECT 909.130 1994.490 910.310 1995.670 ;
        RECT 910.730 1994.490 911.910 1995.670 ;
        RECT 909.130 1816.090 910.310 1817.270 ;
        RECT 910.730 1816.090 911.910 1817.270 ;
        RECT 909.130 1814.490 910.310 1815.670 ;
        RECT 910.730 1814.490 911.910 1815.670 ;
        RECT 909.130 1636.090 910.310 1637.270 ;
        RECT 910.730 1636.090 911.910 1637.270 ;
        RECT 909.130 1634.490 910.310 1635.670 ;
        RECT 910.730 1634.490 911.910 1635.670 ;
        RECT 909.130 1456.090 910.310 1457.270 ;
        RECT 910.730 1456.090 911.910 1457.270 ;
        RECT 909.130 1454.490 910.310 1455.670 ;
        RECT 910.730 1454.490 911.910 1455.670 ;
        RECT 909.130 1276.090 910.310 1277.270 ;
        RECT 910.730 1276.090 911.910 1277.270 ;
        RECT 909.130 1274.490 910.310 1275.670 ;
        RECT 910.730 1274.490 911.910 1275.670 ;
        RECT 909.130 1096.090 910.310 1097.270 ;
        RECT 910.730 1096.090 911.910 1097.270 ;
        RECT 909.130 1094.490 910.310 1095.670 ;
        RECT 910.730 1094.490 911.910 1095.670 ;
        RECT 1089.130 3523.010 1090.310 3524.190 ;
        RECT 1090.730 3523.010 1091.910 3524.190 ;
        RECT 1089.130 3521.410 1090.310 3522.590 ;
        RECT 1090.730 3521.410 1091.910 3522.590 ;
        RECT 1089.130 3436.090 1090.310 3437.270 ;
        RECT 1090.730 3436.090 1091.910 3437.270 ;
        RECT 1089.130 3434.490 1090.310 3435.670 ;
        RECT 1090.730 3434.490 1091.910 3435.670 ;
        RECT 1089.130 3256.090 1090.310 3257.270 ;
        RECT 1090.730 3256.090 1091.910 3257.270 ;
        RECT 1089.130 3254.490 1090.310 3255.670 ;
        RECT 1090.730 3254.490 1091.910 3255.670 ;
        RECT 1089.130 3076.090 1090.310 3077.270 ;
        RECT 1090.730 3076.090 1091.910 3077.270 ;
        RECT 1089.130 3074.490 1090.310 3075.670 ;
        RECT 1090.730 3074.490 1091.910 3075.670 ;
        RECT 1089.130 2896.090 1090.310 2897.270 ;
        RECT 1090.730 2896.090 1091.910 2897.270 ;
        RECT 1089.130 2894.490 1090.310 2895.670 ;
        RECT 1090.730 2894.490 1091.910 2895.670 ;
        RECT 1089.130 2716.090 1090.310 2717.270 ;
        RECT 1090.730 2716.090 1091.910 2717.270 ;
        RECT 1089.130 2714.490 1090.310 2715.670 ;
        RECT 1090.730 2714.490 1091.910 2715.670 ;
        RECT 1089.130 2536.090 1090.310 2537.270 ;
        RECT 1090.730 2536.090 1091.910 2537.270 ;
        RECT 1089.130 2534.490 1090.310 2535.670 ;
        RECT 1090.730 2534.490 1091.910 2535.670 ;
        RECT 1089.130 2356.090 1090.310 2357.270 ;
        RECT 1090.730 2356.090 1091.910 2357.270 ;
        RECT 1089.130 2354.490 1090.310 2355.670 ;
        RECT 1090.730 2354.490 1091.910 2355.670 ;
        RECT 1089.130 2176.090 1090.310 2177.270 ;
        RECT 1090.730 2176.090 1091.910 2177.270 ;
        RECT 1089.130 2174.490 1090.310 2175.670 ;
        RECT 1090.730 2174.490 1091.910 2175.670 ;
        RECT 1089.130 1996.090 1090.310 1997.270 ;
        RECT 1090.730 1996.090 1091.910 1997.270 ;
        RECT 1089.130 1994.490 1090.310 1995.670 ;
        RECT 1090.730 1994.490 1091.910 1995.670 ;
        RECT 1089.130 1816.090 1090.310 1817.270 ;
        RECT 1090.730 1816.090 1091.910 1817.270 ;
        RECT 1089.130 1814.490 1090.310 1815.670 ;
        RECT 1090.730 1814.490 1091.910 1815.670 ;
        RECT 1089.130 1636.090 1090.310 1637.270 ;
        RECT 1090.730 1636.090 1091.910 1637.270 ;
        RECT 1089.130 1634.490 1090.310 1635.670 ;
        RECT 1090.730 1634.490 1091.910 1635.670 ;
        RECT 1089.130 1456.090 1090.310 1457.270 ;
        RECT 1090.730 1456.090 1091.910 1457.270 ;
        RECT 1089.130 1454.490 1090.310 1455.670 ;
        RECT 1090.730 1454.490 1091.910 1455.670 ;
        RECT 1089.130 1276.090 1090.310 1277.270 ;
        RECT 1090.730 1276.090 1091.910 1277.270 ;
        RECT 1089.130 1274.490 1090.310 1275.670 ;
        RECT 1090.730 1274.490 1091.910 1275.670 ;
        RECT 1089.130 1096.090 1090.310 1097.270 ;
        RECT 1090.730 1096.090 1091.910 1097.270 ;
        RECT 1089.130 1094.490 1090.310 1095.670 ;
        RECT 1090.730 1094.490 1091.910 1095.670 ;
        RECT 1269.130 3523.010 1270.310 3524.190 ;
        RECT 1270.730 3523.010 1271.910 3524.190 ;
        RECT 1269.130 3521.410 1270.310 3522.590 ;
        RECT 1270.730 3521.410 1271.910 3522.590 ;
        RECT 1269.130 3436.090 1270.310 3437.270 ;
        RECT 1270.730 3436.090 1271.910 3437.270 ;
        RECT 1269.130 3434.490 1270.310 3435.670 ;
        RECT 1270.730 3434.490 1271.910 3435.670 ;
        RECT 1269.130 3256.090 1270.310 3257.270 ;
        RECT 1270.730 3256.090 1271.910 3257.270 ;
        RECT 1269.130 3254.490 1270.310 3255.670 ;
        RECT 1270.730 3254.490 1271.910 3255.670 ;
        RECT 1269.130 3076.090 1270.310 3077.270 ;
        RECT 1270.730 3076.090 1271.910 3077.270 ;
        RECT 1269.130 3074.490 1270.310 3075.670 ;
        RECT 1270.730 3074.490 1271.910 3075.670 ;
        RECT 1269.130 2896.090 1270.310 2897.270 ;
        RECT 1270.730 2896.090 1271.910 2897.270 ;
        RECT 1269.130 2894.490 1270.310 2895.670 ;
        RECT 1270.730 2894.490 1271.910 2895.670 ;
        RECT 1269.130 2716.090 1270.310 2717.270 ;
        RECT 1270.730 2716.090 1271.910 2717.270 ;
        RECT 1269.130 2714.490 1270.310 2715.670 ;
        RECT 1270.730 2714.490 1271.910 2715.670 ;
        RECT 1269.130 2536.090 1270.310 2537.270 ;
        RECT 1270.730 2536.090 1271.910 2537.270 ;
        RECT 1269.130 2534.490 1270.310 2535.670 ;
        RECT 1270.730 2534.490 1271.910 2535.670 ;
        RECT 1269.130 2356.090 1270.310 2357.270 ;
        RECT 1270.730 2356.090 1271.910 2357.270 ;
        RECT 1269.130 2354.490 1270.310 2355.670 ;
        RECT 1270.730 2354.490 1271.910 2355.670 ;
        RECT 1269.130 2176.090 1270.310 2177.270 ;
        RECT 1270.730 2176.090 1271.910 2177.270 ;
        RECT 1269.130 2174.490 1270.310 2175.670 ;
        RECT 1270.730 2174.490 1271.910 2175.670 ;
        RECT 1269.130 1996.090 1270.310 1997.270 ;
        RECT 1270.730 1996.090 1271.910 1997.270 ;
        RECT 1269.130 1994.490 1270.310 1995.670 ;
        RECT 1270.730 1994.490 1271.910 1995.670 ;
        RECT 1269.130 1816.090 1270.310 1817.270 ;
        RECT 1270.730 1816.090 1271.910 1817.270 ;
        RECT 1269.130 1814.490 1270.310 1815.670 ;
        RECT 1270.730 1814.490 1271.910 1815.670 ;
        RECT 1269.130 1636.090 1270.310 1637.270 ;
        RECT 1270.730 1636.090 1271.910 1637.270 ;
        RECT 1269.130 1634.490 1270.310 1635.670 ;
        RECT 1270.730 1634.490 1271.910 1635.670 ;
        RECT 1269.130 1456.090 1270.310 1457.270 ;
        RECT 1270.730 1456.090 1271.910 1457.270 ;
        RECT 1269.130 1454.490 1270.310 1455.670 ;
        RECT 1270.730 1454.490 1271.910 1455.670 ;
        RECT 1269.130 1276.090 1270.310 1277.270 ;
        RECT 1270.730 1276.090 1271.910 1277.270 ;
        RECT 1269.130 1274.490 1270.310 1275.670 ;
        RECT 1270.730 1274.490 1271.910 1275.670 ;
        RECT 1269.130 1096.090 1270.310 1097.270 ;
        RECT 1270.730 1096.090 1271.910 1097.270 ;
        RECT 1269.130 1094.490 1270.310 1095.670 ;
        RECT 1270.730 1094.490 1271.910 1095.670 ;
        RECT 9.130 916.090 10.310 917.270 ;
        RECT 10.730 916.090 11.910 917.270 ;
        RECT 9.130 914.490 10.310 915.670 ;
        RECT 10.730 914.490 11.910 915.670 ;
        RECT 9.130 736.090 10.310 737.270 ;
        RECT 10.730 736.090 11.910 737.270 ;
        RECT 9.130 734.490 10.310 735.670 ;
        RECT 10.730 734.490 11.910 735.670 ;
        RECT 9.130 556.090 10.310 557.270 ;
        RECT 10.730 556.090 11.910 557.270 ;
        RECT 9.130 554.490 10.310 555.670 ;
        RECT 10.730 554.490 11.910 555.670 ;
        RECT 221.250 916.090 222.430 917.270 ;
        RECT 221.250 914.490 222.430 915.670 ;
        RECT 221.250 736.090 222.430 737.270 ;
        RECT 221.250 734.490 222.430 735.670 ;
        RECT 221.250 556.090 222.430 557.270 ;
        RECT 221.250 554.490 222.430 555.670 ;
        RECT 374.850 916.090 376.030 917.270 ;
        RECT 374.850 914.490 376.030 915.670 ;
        RECT 374.850 736.090 376.030 737.270 ;
        RECT 374.850 734.490 376.030 735.670 ;
        RECT 374.850 556.090 376.030 557.270 ;
        RECT 374.850 554.490 376.030 555.670 ;
        RECT 528.450 916.090 529.630 917.270 ;
        RECT 528.450 914.490 529.630 915.670 ;
        RECT 528.450 736.090 529.630 737.270 ;
        RECT 528.450 734.490 529.630 735.670 ;
        RECT 528.450 556.090 529.630 557.270 ;
        RECT 528.450 554.490 529.630 555.670 ;
        RECT 682.050 916.090 683.230 917.270 ;
        RECT 682.050 914.490 683.230 915.670 ;
        RECT 682.050 736.090 683.230 737.270 ;
        RECT 682.050 734.490 683.230 735.670 ;
        RECT 682.050 556.090 683.230 557.270 ;
        RECT 682.050 554.490 683.230 555.670 ;
        RECT 835.650 916.090 836.830 917.270 ;
        RECT 835.650 914.490 836.830 915.670 ;
        RECT 835.650 736.090 836.830 737.270 ;
        RECT 835.650 734.490 836.830 735.670 ;
        RECT 835.650 556.090 836.830 557.270 ;
        RECT 835.650 554.490 836.830 555.670 ;
        RECT 989.250 916.090 990.430 917.270 ;
        RECT 989.250 914.490 990.430 915.670 ;
        RECT 989.250 736.090 990.430 737.270 ;
        RECT 989.250 734.490 990.430 735.670 ;
        RECT 989.250 556.090 990.430 557.270 ;
        RECT 989.250 554.490 990.430 555.670 ;
        RECT 1269.130 916.090 1270.310 917.270 ;
        RECT 1270.730 916.090 1271.910 917.270 ;
        RECT 1269.130 914.490 1270.310 915.670 ;
        RECT 1270.730 914.490 1271.910 915.670 ;
        RECT 1269.130 736.090 1270.310 737.270 ;
        RECT 1270.730 736.090 1271.910 737.270 ;
        RECT 1269.130 734.490 1270.310 735.670 ;
        RECT 1270.730 734.490 1271.910 735.670 ;
        RECT 1269.130 556.090 1270.310 557.270 ;
        RECT 1270.730 556.090 1271.910 557.270 ;
        RECT 1269.130 554.490 1270.310 555.670 ;
        RECT 1270.730 554.490 1271.910 555.670 ;
        RECT 9.130 376.090 10.310 377.270 ;
        RECT 10.730 376.090 11.910 377.270 ;
        RECT 9.130 374.490 10.310 375.670 ;
        RECT 10.730 374.490 11.910 375.670 ;
        RECT 9.130 196.090 10.310 197.270 ;
        RECT 10.730 196.090 11.910 197.270 ;
        RECT 9.130 194.490 10.310 195.670 ;
        RECT 10.730 194.490 11.910 195.670 ;
        RECT 9.130 16.090 10.310 17.270 ;
        RECT 10.730 16.090 11.910 17.270 ;
        RECT 9.130 14.490 10.310 15.670 ;
        RECT 10.730 14.490 11.910 15.670 ;
        RECT 9.130 -2.910 10.310 -1.730 ;
        RECT 10.730 -2.910 11.910 -1.730 ;
        RECT 9.130 -4.510 10.310 -3.330 ;
        RECT 10.730 -4.510 11.910 -3.330 ;
        RECT 189.130 376.090 190.310 377.270 ;
        RECT 190.730 376.090 191.910 377.270 ;
        RECT 189.130 374.490 190.310 375.670 ;
        RECT 190.730 374.490 191.910 375.670 ;
        RECT 189.130 196.090 190.310 197.270 ;
        RECT 190.730 196.090 191.910 197.270 ;
        RECT 189.130 194.490 190.310 195.670 ;
        RECT 190.730 194.490 191.910 195.670 ;
        RECT 189.130 16.090 190.310 17.270 ;
        RECT 190.730 16.090 191.910 17.270 ;
        RECT 189.130 14.490 190.310 15.670 ;
        RECT 190.730 14.490 191.910 15.670 ;
        RECT 189.130 -2.910 190.310 -1.730 ;
        RECT 190.730 -2.910 191.910 -1.730 ;
        RECT 189.130 -4.510 190.310 -3.330 ;
        RECT 190.730 -4.510 191.910 -3.330 ;
        RECT 369.130 376.090 370.310 377.270 ;
        RECT 370.730 376.090 371.910 377.270 ;
        RECT 369.130 374.490 370.310 375.670 ;
        RECT 370.730 374.490 371.910 375.670 ;
        RECT 369.130 196.090 370.310 197.270 ;
        RECT 370.730 196.090 371.910 197.270 ;
        RECT 369.130 194.490 370.310 195.670 ;
        RECT 370.730 194.490 371.910 195.670 ;
        RECT 369.130 16.090 370.310 17.270 ;
        RECT 370.730 16.090 371.910 17.270 ;
        RECT 369.130 14.490 370.310 15.670 ;
        RECT 370.730 14.490 371.910 15.670 ;
        RECT 369.130 -2.910 370.310 -1.730 ;
        RECT 370.730 -2.910 371.910 -1.730 ;
        RECT 369.130 -4.510 370.310 -3.330 ;
        RECT 370.730 -4.510 371.910 -3.330 ;
        RECT 549.130 376.090 550.310 377.270 ;
        RECT 550.730 376.090 551.910 377.270 ;
        RECT 549.130 374.490 550.310 375.670 ;
        RECT 550.730 374.490 551.910 375.670 ;
        RECT 549.130 196.090 550.310 197.270 ;
        RECT 550.730 196.090 551.910 197.270 ;
        RECT 549.130 194.490 550.310 195.670 ;
        RECT 550.730 194.490 551.910 195.670 ;
        RECT 549.130 16.090 550.310 17.270 ;
        RECT 550.730 16.090 551.910 17.270 ;
        RECT 549.130 14.490 550.310 15.670 ;
        RECT 550.730 14.490 551.910 15.670 ;
        RECT 549.130 -2.910 550.310 -1.730 ;
        RECT 550.730 -2.910 551.910 -1.730 ;
        RECT 549.130 -4.510 550.310 -3.330 ;
        RECT 550.730 -4.510 551.910 -3.330 ;
        RECT 729.130 376.090 730.310 377.270 ;
        RECT 730.730 376.090 731.910 377.270 ;
        RECT 729.130 374.490 730.310 375.670 ;
        RECT 730.730 374.490 731.910 375.670 ;
        RECT 729.130 196.090 730.310 197.270 ;
        RECT 730.730 196.090 731.910 197.270 ;
        RECT 729.130 194.490 730.310 195.670 ;
        RECT 730.730 194.490 731.910 195.670 ;
        RECT 729.130 16.090 730.310 17.270 ;
        RECT 730.730 16.090 731.910 17.270 ;
        RECT 729.130 14.490 730.310 15.670 ;
        RECT 730.730 14.490 731.910 15.670 ;
        RECT 729.130 -2.910 730.310 -1.730 ;
        RECT 730.730 -2.910 731.910 -1.730 ;
        RECT 729.130 -4.510 730.310 -3.330 ;
        RECT 730.730 -4.510 731.910 -3.330 ;
        RECT 909.130 376.090 910.310 377.270 ;
        RECT 910.730 376.090 911.910 377.270 ;
        RECT 909.130 374.490 910.310 375.670 ;
        RECT 910.730 374.490 911.910 375.670 ;
        RECT 909.130 196.090 910.310 197.270 ;
        RECT 910.730 196.090 911.910 197.270 ;
        RECT 909.130 194.490 910.310 195.670 ;
        RECT 910.730 194.490 911.910 195.670 ;
        RECT 909.130 16.090 910.310 17.270 ;
        RECT 910.730 16.090 911.910 17.270 ;
        RECT 909.130 14.490 910.310 15.670 ;
        RECT 910.730 14.490 911.910 15.670 ;
        RECT 909.130 -2.910 910.310 -1.730 ;
        RECT 910.730 -2.910 911.910 -1.730 ;
        RECT 909.130 -4.510 910.310 -3.330 ;
        RECT 910.730 -4.510 911.910 -3.330 ;
        RECT 1089.130 376.090 1090.310 377.270 ;
        RECT 1090.730 376.090 1091.910 377.270 ;
        RECT 1089.130 374.490 1090.310 375.670 ;
        RECT 1090.730 374.490 1091.910 375.670 ;
        RECT 1089.130 196.090 1090.310 197.270 ;
        RECT 1090.730 196.090 1091.910 197.270 ;
        RECT 1089.130 194.490 1090.310 195.670 ;
        RECT 1090.730 194.490 1091.910 195.670 ;
        RECT 1089.130 16.090 1090.310 17.270 ;
        RECT 1090.730 16.090 1091.910 17.270 ;
        RECT 1089.130 14.490 1090.310 15.670 ;
        RECT 1090.730 14.490 1091.910 15.670 ;
        RECT 1089.130 -2.910 1090.310 -1.730 ;
        RECT 1090.730 -2.910 1091.910 -1.730 ;
        RECT 1089.130 -4.510 1090.310 -3.330 ;
        RECT 1090.730 -4.510 1091.910 -3.330 ;
        RECT 1269.130 376.090 1270.310 377.270 ;
        RECT 1270.730 376.090 1271.910 377.270 ;
        RECT 1269.130 374.490 1270.310 375.670 ;
        RECT 1270.730 374.490 1271.910 375.670 ;
        RECT 1269.130 196.090 1270.310 197.270 ;
        RECT 1270.730 196.090 1271.910 197.270 ;
        RECT 1269.130 194.490 1270.310 195.670 ;
        RECT 1270.730 194.490 1271.910 195.670 ;
        RECT 1269.130 16.090 1270.310 17.270 ;
        RECT 1270.730 16.090 1271.910 17.270 ;
        RECT 1269.130 14.490 1270.310 15.670 ;
        RECT 1270.730 14.490 1271.910 15.670 ;
        RECT 1269.130 -2.910 1270.310 -1.730 ;
        RECT 1270.730 -2.910 1271.910 -1.730 ;
        RECT 1269.130 -4.510 1270.310 -3.330 ;
        RECT 1270.730 -4.510 1271.910 -3.330 ;
        RECT 1449.130 3523.010 1450.310 3524.190 ;
        RECT 1450.730 3523.010 1451.910 3524.190 ;
        RECT 1449.130 3521.410 1450.310 3522.590 ;
        RECT 1450.730 3521.410 1451.910 3522.590 ;
        RECT 1449.130 3436.090 1450.310 3437.270 ;
        RECT 1450.730 3436.090 1451.910 3437.270 ;
        RECT 1449.130 3434.490 1450.310 3435.670 ;
        RECT 1450.730 3434.490 1451.910 3435.670 ;
        RECT 1449.130 3256.090 1450.310 3257.270 ;
        RECT 1450.730 3256.090 1451.910 3257.270 ;
        RECT 1449.130 3254.490 1450.310 3255.670 ;
        RECT 1450.730 3254.490 1451.910 3255.670 ;
        RECT 1449.130 3076.090 1450.310 3077.270 ;
        RECT 1450.730 3076.090 1451.910 3077.270 ;
        RECT 1449.130 3074.490 1450.310 3075.670 ;
        RECT 1450.730 3074.490 1451.910 3075.670 ;
        RECT 1449.130 2896.090 1450.310 2897.270 ;
        RECT 1450.730 2896.090 1451.910 2897.270 ;
        RECT 1449.130 2894.490 1450.310 2895.670 ;
        RECT 1450.730 2894.490 1451.910 2895.670 ;
        RECT 1449.130 2716.090 1450.310 2717.270 ;
        RECT 1450.730 2716.090 1451.910 2717.270 ;
        RECT 1449.130 2714.490 1450.310 2715.670 ;
        RECT 1450.730 2714.490 1451.910 2715.670 ;
        RECT 1449.130 2536.090 1450.310 2537.270 ;
        RECT 1450.730 2536.090 1451.910 2537.270 ;
        RECT 1449.130 2534.490 1450.310 2535.670 ;
        RECT 1450.730 2534.490 1451.910 2535.670 ;
        RECT 1449.130 2356.090 1450.310 2357.270 ;
        RECT 1450.730 2356.090 1451.910 2357.270 ;
        RECT 1449.130 2354.490 1450.310 2355.670 ;
        RECT 1450.730 2354.490 1451.910 2355.670 ;
        RECT 1449.130 2176.090 1450.310 2177.270 ;
        RECT 1450.730 2176.090 1451.910 2177.270 ;
        RECT 1449.130 2174.490 1450.310 2175.670 ;
        RECT 1450.730 2174.490 1451.910 2175.670 ;
        RECT 1449.130 1996.090 1450.310 1997.270 ;
        RECT 1450.730 1996.090 1451.910 1997.270 ;
        RECT 1449.130 1994.490 1450.310 1995.670 ;
        RECT 1450.730 1994.490 1451.910 1995.670 ;
        RECT 1449.130 1816.090 1450.310 1817.270 ;
        RECT 1450.730 1816.090 1451.910 1817.270 ;
        RECT 1449.130 1814.490 1450.310 1815.670 ;
        RECT 1450.730 1814.490 1451.910 1815.670 ;
        RECT 1449.130 1636.090 1450.310 1637.270 ;
        RECT 1450.730 1636.090 1451.910 1637.270 ;
        RECT 1449.130 1634.490 1450.310 1635.670 ;
        RECT 1450.730 1634.490 1451.910 1635.670 ;
        RECT 1449.130 1456.090 1450.310 1457.270 ;
        RECT 1450.730 1456.090 1451.910 1457.270 ;
        RECT 1449.130 1454.490 1450.310 1455.670 ;
        RECT 1450.730 1454.490 1451.910 1455.670 ;
        RECT 1449.130 1276.090 1450.310 1277.270 ;
        RECT 1450.730 1276.090 1451.910 1277.270 ;
        RECT 1449.130 1274.490 1450.310 1275.670 ;
        RECT 1450.730 1274.490 1451.910 1275.670 ;
        RECT 1449.130 1096.090 1450.310 1097.270 ;
        RECT 1450.730 1096.090 1451.910 1097.270 ;
        RECT 1449.130 1094.490 1450.310 1095.670 ;
        RECT 1450.730 1094.490 1451.910 1095.670 ;
        RECT 1449.130 916.090 1450.310 917.270 ;
        RECT 1450.730 916.090 1451.910 917.270 ;
        RECT 1449.130 914.490 1450.310 915.670 ;
        RECT 1450.730 914.490 1451.910 915.670 ;
        RECT 1449.130 736.090 1450.310 737.270 ;
        RECT 1450.730 736.090 1451.910 737.270 ;
        RECT 1449.130 734.490 1450.310 735.670 ;
        RECT 1450.730 734.490 1451.910 735.670 ;
        RECT 1449.130 556.090 1450.310 557.270 ;
        RECT 1450.730 556.090 1451.910 557.270 ;
        RECT 1449.130 554.490 1450.310 555.670 ;
        RECT 1450.730 554.490 1451.910 555.670 ;
        RECT 1449.130 376.090 1450.310 377.270 ;
        RECT 1450.730 376.090 1451.910 377.270 ;
        RECT 1449.130 374.490 1450.310 375.670 ;
        RECT 1450.730 374.490 1451.910 375.670 ;
        RECT 1449.130 196.090 1450.310 197.270 ;
        RECT 1450.730 196.090 1451.910 197.270 ;
        RECT 1449.130 194.490 1450.310 195.670 ;
        RECT 1450.730 194.490 1451.910 195.670 ;
        RECT 1449.130 16.090 1450.310 17.270 ;
        RECT 1450.730 16.090 1451.910 17.270 ;
        RECT 1449.130 14.490 1450.310 15.670 ;
        RECT 1450.730 14.490 1451.910 15.670 ;
        RECT 1449.130 -2.910 1450.310 -1.730 ;
        RECT 1450.730 -2.910 1451.910 -1.730 ;
        RECT 1449.130 -4.510 1450.310 -3.330 ;
        RECT 1450.730 -4.510 1451.910 -3.330 ;
        RECT 1629.130 3523.010 1630.310 3524.190 ;
        RECT 1630.730 3523.010 1631.910 3524.190 ;
        RECT 1629.130 3521.410 1630.310 3522.590 ;
        RECT 1630.730 3521.410 1631.910 3522.590 ;
        RECT 1629.130 3436.090 1630.310 3437.270 ;
        RECT 1630.730 3436.090 1631.910 3437.270 ;
        RECT 1629.130 3434.490 1630.310 3435.670 ;
        RECT 1630.730 3434.490 1631.910 3435.670 ;
        RECT 1629.130 3256.090 1630.310 3257.270 ;
        RECT 1630.730 3256.090 1631.910 3257.270 ;
        RECT 1629.130 3254.490 1630.310 3255.670 ;
        RECT 1630.730 3254.490 1631.910 3255.670 ;
        RECT 1629.130 3076.090 1630.310 3077.270 ;
        RECT 1630.730 3076.090 1631.910 3077.270 ;
        RECT 1629.130 3074.490 1630.310 3075.670 ;
        RECT 1630.730 3074.490 1631.910 3075.670 ;
        RECT 1629.130 2896.090 1630.310 2897.270 ;
        RECT 1630.730 2896.090 1631.910 2897.270 ;
        RECT 1629.130 2894.490 1630.310 2895.670 ;
        RECT 1630.730 2894.490 1631.910 2895.670 ;
        RECT 1629.130 2716.090 1630.310 2717.270 ;
        RECT 1630.730 2716.090 1631.910 2717.270 ;
        RECT 1629.130 2714.490 1630.310 2715.670 ;
        RECT 1630.730 2714.490 1631.910 2715.670 ;
        RECT 1629.130 2536.090 1630.310 2537.270 ;
        RECT 1630.730 2536.090 1631.910 2537.270 ;
        RECT 1629.130 2534.490 1630.310 2535.670 ;
        RECT 1630.730 2534.490 1631.910 2535.670 ;
        RECT 1629.130 2356.090 1630.310 2357.270 ;
        RECT 1630.730 2356.090 1631.910 2357.270 ;
        RECT 1629.130 2354.490 1630.310 2355.670 ;
        RECT 1630.730 2354.490 1631.910 2355.670 ;
        RECT 1629.130 2176.090 1630.310 2177.270 ;
        RECT 1630.730 2176.090 1631.910 2177.270 ;
        RECT 1629.130 2174.490 1630.310 2175.670 ;
        RECT 1630.730 2174.490 1631.910 2175.670 ;
        RECT 1629.130 1996.090 1630.310 1997.270 ;
        RECT 1630.730 1996.090 1631.910 1997.270 ;
        RECT 1629.130 1994.490 1630.310 1995.670 ;
        RECT 1630.730 1994.490 1631.910 1995.670 ;
        RECT 1629.130 1816.090 1630.310 1817.270 ;
        RECT 1630.730 1816.090 1631.910 1817.270 ;
        RECT 1629.130 1814.490 1630.310 1815.670 ;
        RECT 1630.730 1814.490 1631.910 1815.670 ;
        RECT 1629.130 1636.090 1630.310 1637.270 ;
        RECT 1630.730 1636.090 1631.910 1637.270 ;
        RECT 1629.130 1634.490 1630.310 1635.670 ;
        RECT 1630.730 1634.490 1631.910 1635.670 ;
        RECT 1629.130 1456.090 1630.310 1457.270 ;
        RECT 1630.730 1456.090 1631.910 1457.270 ;
        RECT 1629.130 1454.490 1630.310 1455.670 ;
        RECT 1630.730 1454.490 1631.910 1455.670 ;
        RECT 1629.130 1276.090 1630.310 1277.270 ;
        RECT 1630.730 1276.090 1631.910 1277.270 ;
        RECT 1629.130 1274.490 1630.310 1275.670 ;
        RECT 1630.730 1274.490 1631.910 1275.670 ;
        RECT 1629.130 1096.090 1630.310 1097.270 ;
        RECT 1630.730 1096.090 1631.910 1097.270 ;
        RECT 1629.130 1094.490 1630.310 1095.670 ;
        RECT 1630.730 1094.490 1631.910 1095.670 ;
        RECT 1629.130 916.090 1630.310 917.270 ;
        RECT 1630.730 916.090 1631.910 917.270 ;
        RECT 1629.130 914.490 1630.310 915.670 ;
        RECT 1630.730 914.490 1631.910 915.670 ;
        RECT 1629.130 736.090 1630.310 737.270 ;
        RECT 1630.730 736.090 1631.910 737.270 ;
        RECT 1629.130 734.490 1630.310 735.670 ;
        RECT 1630.730 734.490 1631.910 735.670 ;
        RECT 1629.130 556.090 1630.310 557.270 ;
        RECT 1630.730 556.090 1631.910 557.270 ;
        RECT 1629.130 554.490 1630.310 555.670 ;
        RECT 1630.730 554.490 1631.910 555.670 ;
        RECT 1629.130 376.090 1630.310 377.270 ;
        RECT 1630.730 376.090 1631.910 377.270 ;
        RECT 1629.130 374.490 1630.310 375.670 ;
        RECT 1630.730 374.490 1631.910 375.670 ;
        RECT 1629.130 196.090 1630.310 197.270 ;
        RECT 1630.730 196.090 1631.910 197.270 ;
        RECT 1629.130 194.490 1630.310 195.670 ;
        RECT 1630.730 194.490 1631.910 195.670 ;
        RECT 1629.130 16.090 1630.310 17.270 ;
        RECT 1630.730 16.090 1631.910 17.270 ;
        RECT 1629.130 14.490 1630.310 15.670 ;
        RECT 1630.730 14.490 1631.910 15.670 ;
        RECT 1629.130 -2.910 1630.310 -1.730 ;
        RECT 1630.730 -2.910 1631.910 -1.730 ;
        RECT 1629.130 -4.510 1630.310 -3.330 ;
        RECT 1630.730 -4.510 1631.910 -3.330 ;
        RECT 1809.130 3523.010 1810.310 3524.190 ;
        RECT 1810.730 3523.010 1811.910 3524.190 ;
        RECT 1809.130 3521.410 1810.310 3522.590 ;
        RECT 1810.730 3521.410 1811.910 3522.590 ;
        RECT 1809.130 3436.090 1810.310 3437.270 ;
        RECT 1810.730 3436.090 1811.910 3437.270 ;
        RECT 1809.130 3434.490 1810.310 3435.670 ;
        RECT 1810.730 3434.490 1811.910 3435.670 ;
        RECT 1809.130 3256.090 1810.310 3257.270 ;
        RECT 1810.730 3256.090 1811.910 3257.270 ;
        RECT 1809.130 3254.490 1810.310 3255.670 ;
        RECT 1810.730 3254.490 1811.910 3255.670 ;
        RECT 1809.130 3076.090 1810.310 3077.270 ;
        RECT 1810.730 3076.090 1811.910 3077.270 ;
        RECT 1809.130 3074.490 1810.310 3075.670 ;
        RECT 1810.730 3074.490 1811.910 3075.670 ;
        RECT 1809.130 2896.090 1810.310 2897.270 ;
        RECT 1810.730 2896.090 1811.910 2897.270 ;
        RECT 1809.130 2894.490 1810.310 2895.670 ;
        RECT 1810.730 2894.490 1811.910 2895.670 ;
        RECT 1809.130 2716.090 1810.310 2717.270 ;
        RECT 1810.730 2716.090 1811.910 2717.270 ;
        RECT 1809.130 2714.490 1810.310 2715.670 ;
        RECT 1810.730 2714.490 1811.910 2715.670 ;
        RECT 1809.130 2536.090 1810.310 2537.270 ;
        RECT 1810.730 2536.090 1811.910 2537.270 ;
        RECT 1809.130 2534.490 1810.310 2535.670 ;
        RECT 1810.730 2534.490 1811.910 2535.670 ;
        RECT 1809.130 2356.090 1810.310 2357.270 ;
        RECT 1810.730 2356.090 1811.910 2357.270 ;
        RECT 1809.130 2354.490 1810.310 2355.670 ;
        RECT 1810.730 2354.490 1811.910 2355.670 ;
        RECT 1809.130 2176.090 1810.310 2177.270 ;
        RECT 1810.730 2176.090 1811.910 2177.270 ;
        RECT 1809.130 2174.490 1810.310 2175.670 ;
        RECT 1810.730 2174.490 1811.910 2175.670 ;
        RECT 1809.130 1996.090 1810.310 1997.270 ;
        RECT 1810.730 1996.090 1811.910 1997.270 ;
        RECT 1809.130 1994.490 1810.310 1995.670 ;
        RECT 1810.730 1994.490 1811.910 1995.670 ;
        RECT 1809.130 1816.090 1810.310 1817.270 ;
        RECT 1810.730 1816.090 1811.910 1817.270 ;
        RECT 1809.130 1814.490 1810.310 1815.670 ;
        RECT 1810.730 1814.490 1811.910 1815.670 ;
        RECT 1809.130 1636.090 1810.310 1637.270 ;
        RECT 1810.730 1636.090 1811.910 1637.270 ;
        RECT 1809.130 1634.490 1810.310 1635.670 ;
        RECT 1810.730 1634.490 1811.910 1635.670 ;
        RECT 1809.130 1456.090 1810.310 1457.270 ;
        RECT 1810.730 1456.090 1811.910 1457.270 ;
        RECT 1809.130 1454.490 1810.310 1455.670 ;
        RECT 1810.730 1454.490 1811.910 1455.670 ;
        RECT 1809.130 1276.090 1810.310 1277.270 ;
        RECT 1810.730 1276.090 1811.910 1277.270 ;
        RECT 1809.130 1274.490 1810.310 1275.670 ;
        RECT 1810.730 1274.490 1811.910 1275.670 ;
        RECT 1809.130 1096.090 1810.310 1097.270 ;
        RECT 1810.730 1096.090 1811.910 1097.270 ;
        RECT 1809.130 1094.490 1810.310 1095.670 ;
        RECT 1810.730 1094.490 1811.910 1095.670 ;
        RECT 1809.130 916.090 1810.310 917.270 ;
        RECT 1810.730 916.090 1811.910 917.270 ;
        RECT 1809.130 914.490 1810.310 915.670 ;
        RECT 1810.730 914.490 1811.910 915.670 ;
        RECT 1809.130 736.090 1810.310 737.270 ;
        RECT 1810.730 736.090 1811.910 737.270 ;
        RECT 1809.130 734.490 1810.310 735.670 ;
        RECT 1810.730 734.490 1811.910 735.670 ;
        RECT 1809.130 556.090 1810.310 557.270 ;
        RECT 1810.730 556.090 1811.910 557.270 ;
        RECT 1809.130 554.490 1810.310 555.670 ;
        RECT 1810.730 554.490 1811.910 555.670 ;
        RECT 1809.130 376.090 1810.310 377.270 ;
        RECT 1810.730 376.090 1811.910 377.270 ;
        RECT 1809.130 374.490 1810.310 375.670 ;
        RECT 1810.730 374.490 1811.910 375.670 ;
        RECT 1809.130 196.090 1810.310 197.270 ;
        RECT 1810.730 196.090 1811.910 197.270 ;
        RECT 1809.130 194.490 1810.310 195.670 ;
        RECT 1810.730 194.490 1811.910 195.670 ;
        RECT 1809.130 16.090 1810.310 17.270 ;
        RECT 1810.730 16.090 1811.910 17.270 ;
        RECT 1809.130 14.490 1810.310 15.670 ;
        RECT 1810.730 14.490 1811.910 15.670 ;
        RECT 1809.130 -2.910 1810.310 -1.730 ;
        RECT 1810.730 -2.910 1811.910 -1.730 ;
        RECT 1809.130 -4.510 1810.310 -3.330 ;
        RECT 1810.730 -4.510 1811.910 -3.330 ;
        RECT 1989.130 3523.010 1990.310 3524.190 ;
        RECT 1990.730 3523.010 1991.910 3524.190 ;
        RECT 1989.130 3521.410 1990.310 3522.590 ;
        RECT 1990.730 3521.410 1991.910 3522.590 ;
        RECT 1989.130 3436.090 1990.310 3437.270 ;
        RECT 1990.730 3436.090 1991.910 3437.270 ;
        RECT 1989.130 3434.490 1990.310 3435.670 ;
        RECT 1990.730 3434.490 1991.910 3435.670 ;
        RECT 1989.130 3256.090 1990.310 3257.270 ;
        RECT 1990.730 3256.090 1991.910 3257.270 ;
        RECT 1989.130 3254.490 1990.310 3255.670 ;
        RECT 1990.730 3254.490 1991.910 3255.670 ;
        RECT 1989.130 3076.090 1990.310 3077.270 ;
        RECT 1990.730 3076.090 1991.910 3077.270 ;
        RECT 1989.130 3074.490 1990.310 3075.670 ;
        RECT 1990.730 3074.490 1991.910 3075.670 ;
        RECT 1989.130 2896.090 1990.310 2897.270 ;
        RECT 1990.730 2896.090 1991.910 2897.270 ;
        RECT 1989.130 2894.490 1990.310 2895.670 ;
        RECT 1990.730 2894.490 1991.910 2895.670 ;
        RECT 1989.130 2716.090 1990.310 2717.270 ;
        RECT 1990.730 2716.090 1991.910 2717.270 ;
        RECT 1989.130 2714.490 1990.310 2715.670 ;
        RECT 1990.730 2714.490 1991.910 2715.670 ;
        RECT 1989.130 2536.090 1990.310 2537.270 ;
        RECT 1990.730 2536.090 1991.910 2537.270 ;
        RECT 1989.130 2534.490 1990.310 2535.670 ;
        RECT 1990.730 2534.490 1991.910 2535.670 ;
        RECT 1989.130 2356.090 1990.310 2357.270 ;
        RECT 1990.730 2356.090 1991.910 2357.270 ;
        RECT 1989.130 2354.490 1990.310 2355.670 ;
        RECT 1990.730 2354.490 1991.910 2355.670 ;
        RECT 1989.130 2176.090 1990.310 2177.270 ;
        RECT 1990.730 2176.090 1991.910 2177.270 ;
        RECT 1989.130 2174.490 1990.310 2175.670 ;
        RECT 1990.730 2174.490 1991.910 2175.670 ;
        RECT 1989.130 1996.090 1990.310 1997.270 ;
        RECT 1990.730 1996.090 1991.910 1997.270 ;
        RECT 1989.130 1994.490 1990.310 1995.670 ;
        RECT 1990.730 1994.490 1991.910 1995.670 ;
        RECT 1989.130 1816.090 1990.310 1817.270 ;
        RECT 1990.730 1816.090 1991.910 1817.270 ;
        RECT 1989.130 1814.490 1990.310 1815.670 ;
        RECT 1990.730 1814.490 1991.910 1815.670 ;
        RECT 1989.130 1636.090 1990.310 1637.270 ;
        RECT 1990.730 1636.090 1991.910 1637.270 ;
        RECT 1989.130 1634.490 1990.310 1635.670 ;
        RECT 1990.730 1634.490 1991.910 1635.670 ;
        RECT 1989.130 1456.090 1990.310 1457.270 ;
        RECT 1990.730 1456.090 1991.910 1457.270 ;
        RECT 1989.130 1454.490 1990.310 1455.670 ;
        RECT 1990.730 1454.490 1991.910 1455.670 ;
        RECT 1989.130 1276.090 1990.310 1277.270 ;
        RECT 1990.730 1276.090 1991.910 1277.270 ;
        RECT 1989.130 1274.490 1990.310 1275.670 ;
        RECT 1990.730 1274.490 1991.910 1275.670 ;
        RECT 1989.130 1096.090 1990.310 1097.270 ;
        RECT 1990.730 1096.090 1991.910 1097.270 ;
        RECT 1989.130 1094.490 1990.310 1095.670 ;
        RECT 1990.730 1094.490 1991.910 1095.670 ;
        RECT 1989.130 916.090 1990.310 917.270 ;
        RECT 1990.730 916.090 1991.910 917.270 ;
        RECT 1989.130 914.490 1990.310 915.670 ;
        RECT 1990.730 914.490 1991.910 915.670 ;
        RECT 1989.130 736.090 1990.310 737.270 ;
        RECT 1990.730 736.090 1991.910 737.270 ;
        RECT 1989.130 734.490 1990.310 735.670 ;
        RECT 1990.730 734.490 1991.910 735.670 ;
        RECT 1989.130 556.090 1990.310 557.270 ;
        RECT 1990.730 556.090 1991.910 557.270 ;
        RECT 1989.130 554.490 1990.310 555.670 ;
        RECT 1990.730 554.490 1991.910 555.670 ;
        RECT 1989.130 376.090 1990.310 377.270 ;
        RECT 1990.730 376.090 1991.910 377.270 ;
        RECT 1989.130 374.490 1990.310 375.670 ;
        RECT 1990.730 374.490 1991.910 375.670 ;
        RECT 1989.130 196.090 1990.310 197.270 ;
        RECT 1990.730 196.090 1991.910 197.270 ;
        RECT 1989.130 194.490 1990.310 195.670 ;
        RECT 1990.730 194.490 1991.910 195.670 ;
        RECT 1989.130 16.090 1990.310 17.270 ;
        RECT 1990.730 16.090 1991.910 17.270 ;
        RECT 1989.130 14.490 1990.310 15.670 ;
        RECT 1990.730 14.490 1991.910 15.670 ;
        RECT 1989.130 -2.910 1990.310 -1.730 ;
        RECT 1990.730 -2.910 1991.910 -1.730 ;
        RECT 1989.130 -4.510 1990.310 -3.330 ;
        RECT 1990.730 -4.510 1991.910 -3.330 ;
        RECT 2169.130 3523.010 2170.310 3524.190 ;
        RECT 2170.730 3523.010 2171.910 3524.190 ;
        RECT 2169.130 3521.410 2170.310 3522.590 ;
        RECT 2170.730 3521.410 2171.910 3522.590 ;
        RECT 2169.130 3436.090 2170.310 3437.270 ;
        RECT 2170.730 3436.090 2171.910 3437.270 ;
        RECT 2169.130 3434.490 2170.310 3435.670 ;
        RECT 2170.730 3434.490 2171.910 3435.670 ;
        RECT 2169.130 3256.090 2170.310 3257.270 ;
        RECT 2170.730 3256.090 2171.910 3257.270 ;
        RECT 2169.130 3254.490 2170.310 3255.670 ;
        RECT 2170.730 3254.490 2171.910 3255.670 ;
        RECT 2169.130 3076.090 2170.310 3077.270 ;
        RECT 2170.730 3076.090 2171.910 3077.270 ;
        RECT 2169.130 3074.490 2170.310 3075.670 ;
        RECT 2170.730 3074.490 2171.910 3075.670 ;
        RECT 2169.130 2896.090 2170.310 2897.270 ;
        RECT 2170.730 2896.090 2171.910 2897.270 ;
        RECT 2169.130 2894.490 2170.310 2895.670 ;
        RECT 2170.730 2894.490 2171.910 2895.670 ;
        RECT 2169.130 2716.090 2170.310 2717.270 ;
        RECT 2170.730 2716.090 2171.910 2717.270 ;
        RECT 2169.130 2714.490 2170.310 2715.670 ;
        RECT 2170.730 2714.490 2171.910 2715.670 ;
        RECT 2169.130 2536.090 2170.310 2537.270 ;
        RECT 2170.730 2536.090 2171.910 2537.270 ;
        RECT 2169.130 2534.490 2170.310 2535.670 ;
        RECT 2170.730 2534.490 2171.910 2535.670 ;
        RECT 2169.130 2356.090 2170.310 2357.270 ;
        RECT 2170.730 2356.090 2171.910 2357.270 ;
        RECT 2169.130 2354.490 2170.310 2355.670 ;
        RECT 2170.730 2354.490 2171.910 2355.670 ;
        RECT 2169.130 2176.090 2170.310 2177.270 ;
        RECT 2170.730 2176.090 2171.910 2177.270 ;
        RECT 2169.130 2174.490 2170.310 2175.670 ;
        RECT 2170.730 2174.490 2171.910 2175.670 ;
        RECT 2169.130 1996.090 2170.310 1997.270 ;
        RECT 2170.730 1996.090 2171.910 1997.270 ;
        RECT 2169.130 1994.490 2170.310 1995.670 ;
        RECT 2170.730 1994.490 2171.910 1995.670 ;
        RECT 2169.130 1816.090 2170.310 1817.270 ;
        RECT 2170.730 1816.090 2171.910 1817.270 ;
        RECT 2169.130 1814.490 2170.310 1815.670 ;
        RECT 2170.730 1814.490 2171.910 1815.670 ;
        RECT 2169.130 1636.090 2170.310 1637.270 ;
        RECT 2170.730 1636.090 2171.910 1637.270 ;
        RECT 2169.130 1634.490 2170.310 1635.670 ;
        RECT 2170.730 1634.490 2171.910 1635.670 ;
        RECT 2169.130 1456.090 2170.310 1457.270 ;
        RECT 2170.730 1456.090 2171.910 1457.270 ;
        RECT 2169.130 1454.490 2170.310 1455.670 ;
        RECT 2170.730 1454.490 2171.910 1455.670 ;
        RECT 2169.130 1276.090 2170.310 1277.270 ;
        RECT 2170.730 1276.090 2171.910 1277.270 ;
        RECT 2169.130 1274.490 2170.310 1275.670 ;
        RECT 2170.730 1274.490 2171.910 1275.670 ;
        RECT 2169.130 1096.090 2170.310 1097.270 ;
        RECT 2170.730 1096.090 2171.910 1097.270 ;
        RECT 2169.130 1094.490 2170.310 1095.670 ;
        RECT 2170.730 1094.490 2171.910 1095.670 ;
        RECT 2169.130 916.090 2170.310 917.270 ;
        RECT 2170.730 916.090 2171.910 917.270 ;
        RECT 2169.130 914.490 2170.310 915.670 ;
        RECT 2170.730 914.490 2171.910 915.670 ;
        RECT 2169.130 736.090 2170.310 737.270 ;
        RECT 2170.730 736.090 2171.910 737.270 ;
        RECT 2169.130 734.490 2170.310 735.670 ;
        RECT 2170.730 734.490 2171.910 735.670 ;
        RECT 2169.130 556.090 2170.310 557.270 ;
        RECT 2170.730 556.090 2171.910 557.270 ;
        RECT 2169.130 554.490 2170.310 555.670 ;
        RECT 2170.730 554.490 2171.910 555.670 ;
        RECT 2169.130 376.090 2170.310 377.270 ;
        RECT 2170.730 376.090 2171.910 377.270 ;
        RECT 2169.130 374.490 2170.310 375.670 ;
        RECT 2170.730 374.490 2171.910 375.670 ;
        RECT 2169.130 196.090 2170.310 197.270 ;
        RECT 2170.730 196.090 2171.910 197.270 ;
        RECT 2169.130 194.490 2170.310 195.670 ;
        RECT 2170.730 194.490 2171.910 195.670 ;
        RECT 2169.130 16.090 2170.310 17.270 ;
        RECT 2170.730 16.090 2171.910 17.270 ;
        RECT 2169.130 14.490 2170.310 15.670 ;
        RECT 2170.730 14.490 2171.910 15.670 ;
        RECT 2169.130 -2.910 2170.310 -1.730 ;
        RECT 2170.730 -2.910 2171.910 -1.730 ;
        RECT 2169.130 -4.510 2170.310 -3.330 ;
        RECT 2170.730 -4.510 2171.910 -3.330 ;
        RECT 2349.130 3523.010 2350.310 3524.190 ;
        RECT 2350.730 3523.010 2351.910 3524.190 ;
        RECT 2349.130 3521.410 2350.310 3522.590 ;
        RECT 2350.730 3521.410 2351.910 3522.590 ;
        RECT 2349.130 3436.090 2350.310 3437.270 ;
        RECT 2350.730 3436.090 2351.910 3437.270 ;
        RECT 2349.130 3434.490 2350.310 3435.670 ;
        RECT 2350.730 3434.490 2351.910 3435.670 ;
        RECT 2349.130 3256.090 2350.310 3257.270 ;
        RECT 2350.730 3256.090 2351.910 3257.270 ;
        RECT 2349.130 3254.490 2350.310 3255.670 ;
        RECT 2350.730 3254.490 2351.910 3255.670 ;
        RECT 2349.130 3076.090 2350.310 3077.270 ;
        RECT 2350.730 3076.090 2351.910 3077.270 ;
        RECT 2349.130 3074.490 2350.310 3075.670 ;
        RECT 2350.730 3074.490 2351.910 3075.670 ;
        RECT 2349.130 2896.090 2350.310 2897.270 ;
        RECT 2350.730 2896.090 2351.910 2897.270 ;
        RECT 2349.130 2894.490 2350.310 2895.670 ;
        RECT 2350.730 2894.490 2351.910 2895.670 ;
        RECT 2349.130 2716.090 2350.310 2717.270 ;
        RECT 2350.730 2716.090 2351.910 2717.270 ;
        RECT 2349.130 2714.490 2350.310 2715.670 ;
        RECT 2350.730 2714.490 2351.910 2715.670 ;
        RECT 2349.130 2536.090 2350.310 2537.270 ;
        RECT 2350.730 2536.090 2351.910 2537.270 ;
        RECT 2349.130 2534.490 2350.310 2535.670 ;
        RECT 2350.730 2534.490 2351.910 2535.670 ;
        RECT 2349.130 2356.090 2350.310 2357.270 ;
        RECT 2350.730 2356.090 2351.910 2357.270 ;
        RECT 2349.130 2354.490 2350.310 2355.670 ;
        RECT 2350.730 2354.490 2351.910 2355.670 ;
        RECT 2349.130 2176.090 2350.310 2177.270 ;
        RECT 2350.730 2176.090 2351.910 2177.270 ;
        RECT 2349.130 2174.490 2350.310 2175.670 ;
        RECT 2350.730 2174.490 2351.910 2175.670 ;
        RECT 2349.130 1996.090 2350.310 1997.270 ;
        RECT 2350.730 1996.090 2351.910 1997.270 ;
        RECT 2349.130 1994.490 2350.310 1995.670 ;
        RECT 2350.730 1994.490 2351.910 1995.670 ;
        RECT 2349.130 1816.090 2350.310 1817.270 ;
        RECT 2350.730 1816.090 2351.910 1817.270 ;
        RECT 2349.130 1814.490 2350.310 1815.670 ;
        RECT 2350.730 1814.490 2351.910 1815.670 ;
        RECT 2349.130 1636.090 2350.310 1637.270 ;
        RECT 2350.730 1636.090 2351.910 1637.270 ;
        RECT 2349.130 1634.490 2350.310 1635.670 ;
        RECT 2350.730 1634.490 2351.910 1635.670 ;
        RECT 2349.130 1456.090 2350.310 1457.270 ;
        RECT 2350.730 1456.090 2351.910 1457.270 ;
        RECT 2349.130 1454.490 2350.310 1455.670 ;
        RECT 2350.730 1454.490 2351.910 1455.670 ;
        RECT 2349.130 1276.090 2350.310 1277.270 ;
        RECT 2350.730 1276.090 2351.910 1277.270 ;
        RECT 2349.130 1274.490 2350.310 1275.670 ;
        RECT 2350.730 1274.490 2351.910 1275.670 ;
        RECT 2349.130 1096.090 2350.310 1097.270 ;
        RECT 2350.730 1096.090 2351.910 1097.270 ;
        RECT 2349.130 1094.490 2350.310 1095.670 ;
        RECT 2350.730 1094.490 2351.910 1095.670 ;
        RECT 2349.130 916.090 2350.310 917.270 ;
        RECT 2350.730 916.090 2351.910 917.270 ;
        RECT 2349.130 914.490 2350.310 915.670 ;
        RECT 2350.730 914.490 2351.910 915.670 ;
        RECT 2349.130 736.090 2350.310 737.270 ;
        RECT 2350.730 736.090 2351.910 737.270 ;
        RECT 2349.130 734.490 2350.310 735.670 ;
        RECT 2350.730 734.490 2351.910 735.670 ;
        RECT 2349.130 556.090 2350.310 557.270 ;
        RECT 2350.730 556.090 2351.910 557.270 ;
        RECT 2349.130 554.490 2350.310 555.670 ;
        RECT 2350.730 554.490 2351.910 555.670 ;
        RECT 2349.130 376.090 2350.310 377.270 ;
        RECT 2350.730 376.090 2351.910 377.270 ;
        RECT 2349.130 374.490 2350.310 375.670 ;
        RECT 2350.730 374.490 2351.910 375.670 ;
        RECT 2349.130 196.090 2350.310 197.270 ;
        RECT 2350.730 196.090 2351.910 197.270 ;
        RECT 2349.130 194.490 2350.310 195.670 ;
        RECT 2350.730 194.490 2351.910 195.670 ;
        RECT 2349.130 16.090 2350.310 17.270 ;
        RECT 2350.730 16.090 2351.910 17.270 ;
        RECT 2349.130 14.490 2350.310 15.670 ;
        RECT 2350.730 14.490 2351.910 15.670 ;
        RECT 2349.130 -2.910 2350.310 -1.730 ;
        RECT 2350.730 -2.910 2351.910 -1.730 ;
        RECT 2349.130 -4.510 2350.310 -3.330 ;
        RECT 2350.730 -4.510 2351.910 -3.330 ;
        RECT 2529.130 3523.010 2530.310 3524.190 ;
        RECT 2530.730 3523.010 2531.910 3524.190 ;
        RECT 2529.130 3521.410 2530.310 3522.590 ;
        RECT 2530.730 3521.410 2531.910 3522.590 ;
        RECT 2529.130 3436.090 2530.310 3437.270 ;
        RECT 2530.730 3436.090 2531.910 3437.270 ;
        RECT 2529.130 3434.490 2530.310 3435.670 ;
        RECT 2530.730 3434.490 2531.910 3435.670 ;
        RECT 2529.130 3256.090 2530.310 3257.270 ;
        RECT 2530.730 3256.090 2531.910 3257.270 ;
        RECT 2529.130 3254.490 2530.310 3255.670 ;
        RECT 2530.730 3254.490 2531.910 3255.670 ;
        RECT 2529.130 3076.090 2530.310 3077.270 ;
        RECT 2530.730 3076.090 2531.910 3077.270 ;
        RECT 2529.130 3074.490 2530.310 3075.670 ;
        RECT 2530.730 3074.490 2531.910 3075.670 ;
        RECT 2529.130 2896.090 2530.310 2897.270 ;
        RECT 2530.730 2896.090 2531.910 2897.270 ;
        RECT 2529.130 2894.490 2530.310 2895.670 ;
        RECT 2530.730 2894.490 2531.910 2895.670 ;
        RECT 2529.130 2716.090 2530.310 2717.270 ;
        RECT 2530.730 2716.090 2531.910 2717.270 ;
        RECT 2529.130 2714.490 2530.310 2715.670 ;
        RECT 2530.730 2714.490 2531.910 2715.670 ;
        RECT 2529.130 2536.090 2530.310 2537.270 ;
        RECT 2530.730 2536.090 2531.910 2537.270 ;
        RECT 2529.130 2534.490 2530.310 2535.670 ;
        RECT 2530.730 2534.490 2531.910 2535.670 ;
        RECT 2529.130 2356.090 2530.310 2357.270 ;
        RECT 2530.730 2356.090 2531.910 2357.270 ;
        RECT 2529.130 2354.490 2530.310 2355.670 ;
        RECT 2530.730 2354.490 2531.910 2355.670 ;
        RECT 2529.130 2176.090 2530.310 2177.270 ;
        RECT 2530.730 2176.090 2531.910 2177.270 ;
        RECT 2529.130 2174.490 2530.310 2175.670 ;
        RECT 2530.730 2174.490 2531.910 2175.670 ;
        RECT 2529.130 1996.090 2530.310 1997.270 ;
        RECT 2530.730 1996.090 2531.910 1997.270 ;
        RECT 2529.130 1994.490 2530.310 1995.670 ;
        RECT 2530.730 1994.490 2531.910 1995.670 ;
        RECT 2529.130 1816.090 2530.310 1817.270 ;
        RECT 2530.730 1816.090 2531.910 1817.270 ;
        RECT 2529.130 1814.490 2530.310 1815.670 ;
        RECT 2530.730 1814.490 2531.910 1815.670 ;
        RECT 2529.130 1636.090 2530.310 1637.270 ;
        RECT 2530.730 1636.090 2531.910 1637.270 ;
        RECT 2529.130 1634.490 2530.310 1635.670 ;
        RECT 2530.730 1634.490 2531.910 1635.670 ;
        RECT 2529.130 1456.090 2530.310 1457.270 ;
        RECT 2530.730 1456.090 2531.910 1457.270 ;
        RECT 2529.130 1454.490 2530.310 1455.670 ;
        RECT 2530.730 1454.490 2531.910 1455.670 ;
        RECT 2529.130 1276.090 2530.310 1277.270 ;
        RECT 2530.730 1276.090 2531.910 1277.270 ;
        RECT 2529.130 1274.490 2530.310 1275.670 ;
        RECT 2530.730 1274.490 2531.910 1275.670 ;
        RECT 2529.130 1096.090 2530.310 1097.270 ;
        RECT 2530.730 1096.090 2531.910 1097.270 ;
        RECT 2529.130 1094.490 2530.310 1095.670 ;
        RECT 2530.730 1094.490 2531.910 1095.670 ;
        RECT 2529.130 916.090 2530.310 917.270 ;
        RECT 2530.730 916.090 2531.910 917.270 ;
        RECT 2529.130 914.490 2530.310 915.670 ;
        RECT 2530.730 914.490 2531.910 915.670 ;
        RECT 2529.130 736.090 2530.310 737.270 ;
        RECT 2530.730 736.090 2531.910 737.270 ;
        RECT 2529.130 734.490 2530.310 735.670 ;
        RECT 2530.730 734.490 2531.910 735.670 ;
        RECT 2529.130 556.090 2530.310 557.270 ;
        RECT 2530.730 556.090 2531.910 557.270 ;
        RECT 2529.130 554.490 2530.310 555.670 ;
        RECT 2530.730 554.490 2531.910 555.670 ;
        RECT 2529.130 376.090 2530.310 377.270 ;
        RECT 2530.730 376.090 2531.910 377.270 ;
        RECT 2529.130 374.490 2530.310 375.670 ;
        RECT 2530.730 374.490 2531.910 375.670 ;
        RECT 2529.130 196.090 2530.310 197.270 ;
        RECT 2530.730 196.090 2531.910 197.270 ;
        RECT 2529.130 194.490 2530.310 195.670 ;
        RECT 2530.730 194.490 2531.910 195.670 ;
        RECT 2529.130 16.090 2530.310 17.270 ;
        RECT 2530.730 16.090 2531.910 17.270 ;
        RECT 2529.130 14.490 2530.310 15.670 ;
        RECT 2530.730 14.490 2531.910 15.670 ;
        RECT 2529.130 -2.910 2530.310 -1.730 ;
        RECT 2530.730 -2.910 2531.910 -1.730 ;
        RECT 2529.130 -4.510 2530.310 -3.330 ;
        RECT 2530.730 -4.510 2531.910 -3.330 ;
        RECT 2709.130 3523.010 2710.310 3524.190 ;
        RECT 2710.730 3523.010 2711.910 3524.190 ;
        RECT 2709.130 3521.410 2710.310 3522.590 ;
        RECT 2710.730 3521.410 2711.910 3522.590 ;
        RECT 2709.130 3436.090 2710.310 3437.270 ;
        RECT 2710.730 3436.090 2711.910 3437.270 ;
        RECT 2709.130 3434.490 2710.310 3435.670 ;
        RECT 2710.730 3434.490 2711.910 3435.670 ;
        RECT 2709.130 3256.090 2710.310 3257.270 ;
        RECT 2710.730 3256.090 2711.910 3257.270 ;
        RECT 2709.130 3254.490 2710.310 3255.670 ;
        RECT 2710.730 3254.490 2711.910 3255.670 ;
        RECT 2709.130 3076.090 2710.310 3077.270 ;
        RECT 2710.730 3076.090 2711.910 3077.270 ;
        RECT 2709.130 3074.490 2710.310 3075.670 ;
        RECT 2710.730 3074.490 2711.910 3075.670 ;
        RECT 2709.130 2896.090 2710.310 2897.270 ;
        RECT 2710.730 2896.090 2711.910 2897.270 ;
        RECT 2709.130 2894.490 2710.310 2895.670 ;
        RECT 2710.730 2894.490 2711.910 2895.670 ;
        RECT 2709.130 2716.090 2710.310 2717.270 ;
        RECT 2710.730 2716.090 2711.910 2717.270 ;
        RECT 2709.130 2714.490 2710.310 2715.670 ;
        RECT 2710.730 2714.490 2711.910 2715.670 ;
        RECT 2709.130 2536.090 2710.310 2537.270 ;
        RECT 2710.730 2536.090 2711.910 2537.270 ;
        RECT 2709.130 2534.490 2710.310 2535.670 ;
        RECT 2710.730 2534.490 2711.910 2535.670 ;
        RECT 2709.130 2356.090 2710.310 2357.270 ;
        RECT 2710.730 2356.090 2711.910 2357.270 ;
        RECT 2709.130 2354.490 2710.310 2355.670 ;
        RECT 2710.730 2354.490 2711.910 2355.670 ;
        RECT 2709.130 2176.090 2710.310 2177.270 ;
        RECT 2710.730 2176.090 2711.910 2177.270 ;
        RECT 2709.130 2174.490 2710.310 2175.670 ;
        RECT 2710.730 2174.490 2711.910 2175.670 ;
        RECT 2709.130 1996.090 2710.310 1997.270 ;
        RECT 2710.730 1996.090 2711.910 1997.270 ;
        RECT 2709.130 1994.490 2710.310 1995.670 ;
        RECT 2710.730 1994.490 2711.910 1995.670 ;
        RECT 2709.130 1816.090 2710.310 1817.270 ;
        RECT 2710.730 1816.090 2711.910 1817.270 ;
        RECT 2709.130 1814.490 2710.310 1815.670 ;
        RECT 2710.730 1814.490 2711.910 1815.670 ;
        RECT 2709.130 1636.090 2710.310 1637.270 ;
        RECT 2710.730 1636.090 2711.910 1637.270 ;
        RECT 2709.130 1634.490 2710.310 1635.670 ;
        RECT 2710.730 1634.490 2711.910 1635.670 ;
        RECT 2709.130 1456.090 2710.310 1457.270 ;
        RECT 2710.730 1456.090 2711.910 1457.270 ;
        RECT 2709.130 1454.490 2710.310 1455.670 ;
        RECT 2710.730 1454.490 2711.910 1455.670 ;
        RECT 2709.130 1276.090 2710.310 1277.270 ;
        RECT 2710.730 1276.090 2711.910 1277.270 ;
        RECT 2709.130 1274.490 2710.310 1275.670 ;
        RECT 2710.730 1274.490 2711.910 1275.670 ;
        RECT 2709.130 1096.090 2710.310 1097.270 ;
        RECT 2710.730 1096.090 2711.910 1097.270 ;
        RECT 2709.130 1094.490 2710.310 1095.670 ;
        RECT 2710.730 1094.490 2711.910 1095.670 ;
        RECT 2709.130 916.090 2710.310 917.270 ;
        RECT 2710.730 916.090 2711.910 917.270 ;
        RECT 2709.130 914.490 2710.310 915.670 ;
        RECT 2710.730 914.490 2711.910 915.670 ;
        RECT 2709.130 736.090 2710.310 737.270 ;
        RECT 2710.730 736.090 2711.910 737.270 ;
        RECT 2709.130 734.490 2710.310 735.670 ;
        RECT 2710.730 734.490 2711.910 735.670 ;
        RECT 2709.130 556.090 2710.310 557.270 ;
        RECT 2710.730 556.090 2711.910 557.270 ;
        RECT 2709.130 554.490 2710.310 555.670 ;
        RECT 2710.730 554.490 2711.910 555.670 ;
        RECT 2709.130 376.090 2710.310 377.270 ;
        RECT 2710.730 376.090 2711.910 377.270 ;
        RECT 2709.130 374.490 2710.310 375.670 ;
        RECT 2710.730 374.490 2711.910 375.670 ;
        RECT 2709.130 196.090 2710.310 197.270 ;
        RECT 2710.730 196.090 2711.910 197.270 ;
        RECT 2709.130 194.490 2710.310 195.670 ;
        RECT 2710.730 194.490 2711.910 195.670 ;
        RECT 2709.130 16.090 2710.310 17.270 ;
        RECT 2710.730 16.090 2711.910 17.270 ;
        RECT 2709.130 14.490 2710.310 15.670 ;
        RECT 2710.730 14.490 2711.910 15.670 ;
        RECT 2709.130 -2.910 2710.310 -1.730 ;
        RECT 2710.730 -2.910 2711.910 -1.730 ;
        RECT 2709.130 -4.510 2710.310 -3.330 ;
        RECT 2710.730 -4.510 2711.910 -3.330 ;
        RECT 2889.130 3523.010 2890.310 3524.190 ;
        RECT 2890.730 3523.010 2891.910 3524.190 ;
        RECT 2889.130 3521.410 2890.310 3522.590 ;
        RECT 2890.730 3521.410 2891.910 3522.590 ;
        RECT 2889.130 3436.090 2890.310 3437.270 ;
        RECT 2890.730 3436.090 2891.910 3437.270 ;
        RECT 2889.130 3434.490 2890.310 3435.670 ;
        RECT 2890.730 3434.490 2891.910 3435.670 ;
        RECT 2889.130 3256.090 2890.310 3257.270 ;
        RECT 2890.730 3256.090 2891.910 3257.270 ;
        RECT 2889.130 3254.490 2890.310 3255.670 ;
        RECT 2890.730 3254.490 2891.910 3255.670 ;
        RECT 2889.130 3076.090 2890.310 3077.270 ;
        RECT 2890.730 3076.090 2891.910 3077.270 ;
        RECT 2889.130 3074.490 2890.310 3075.670 ;
        RECT 2890.730 3074.490 2891.910 3075.670 ;
        RECT 2889.130 2896.090 2890.310 2897.270 ;
        RECT 2890.730 2896.090 2891.910 2897.270 ;
        RECT 2889.130 2894.490 2890.310 2895.670 ;
        RECT 2890.730 2894.490 2891.910 2895.670 ;
        RECT 2889.130 2716.090 2890.310 2717.270 ;
        RECT 2890.730 2716.090 2891.910 2717.270 ;
        RECT 2889.130 2714.490 2890.310 2715.670 ;
        RECT 2890.730 2714.490 2891.910 2715.670 ;
        RECT 2889.130 2536.090 2890.310 2537.270 ;
        RECT 2890.730 2536.090 2891.910 2537.270 ;
        RECT 2889.130 2534.490 2890.310 2535.670 ;
        RECT 2890.730 2534.490 2891.910 2535.670 ;
        RECT 2889.130 2356.090 2890.310 2357.270 ;
        RECT 2890.730 2356.090 2891.910 2357.270 ;
        RECT 2889.130 2354.490 2890.310 2355.670 ;
        RECT 2890.730 2354.490 2891.910 2355.670 ;
        RECT 2889.130 2176.090 2890.310 2177.270 ;
        RECT 2890.730 2176.090 2891.910 2177.270 ;
        RECT 2889.130 2174.490 2890.310 2175.670 ;
        RECT 2890.730 2174.490 2891.910 2175.670 ;
        RECT 2889.130 1996.090 2890.310 1997.270 ;
        RECT 2890.730 1996.090 2891.910 1997.270 ;
        RECT 2889.130 1994.490 2890.310 1995.670 ;
        RECT 2890.730 1994.490 2891.910 1995.670 ;
        RECT 2889.130 1816.090 2890.310 1817.270 ;
        RECT 2890.730 1816.090 2891.910 1817.270 ;
        RECT 2889.130 1814.490 2890.310 1815.670 ;
        RECT 2890.730 1814.490 2891.910 1815.670 ;
        RECT 2889.130 1636.090 2890.310 1637.270 ;
        RECT 2890.730 1636.090 2891.910 1637.270 ;
        RECT 2889.130 1634.490 2890.310 1635.670 ;
        RECT 2890.730 1634.490 2891.910 1635.670 ;
        RECT 2889.130 1456.090 2890.310 1457.270 ;
        RECT 2890.730 1456.090 2891.910 1457.270 ;
        RECT 2889.130 1454.490 2890.310 1455.670 ;
        RECT 2890.730 1454.490 2891.910 1455.670 ;
        RECT 2889.130 1276.090 2890.310 1277.270 ;
        RECT 2890.730 1276.090 2891.910 1277.270 ;
        RECT 2889.130 1274.490 2890.310 1275.670 ;
        RECT 2890.730 1274.490 2891.910 1275.670 ;
        RECT 2889.130 1096.090 2890.310 1097.270 ;
        RECT 2890.730 1096.090 2891.910 1097.270 ;
        RECT 2889.130 1094.490 2890.310 1095.670 ;
        RECT 2890.730 1094.490 2891.910 1095.670 ;
        RECT 2889.130 916.090 2890.310 917.270 ;
        RECT 2890.730 916.090 2891.910 917.270 ;
        RECT 2889.130 914.490 2890.310 915.670 ;
        RECT 2890.730 914.490 2891.910 915.670 ;
        RECT 2889.130 736.090 2890.310 737.270 ;
        RECT 2890.730 736.090 2891.910 737.270 ;
        RECT 2889.130 734.490 2890.310 735.670 ;
        RECT 2890.730 734.490 2891.910 735.670 ;
        RECT 2889.130 556.090 2890.310 557.270 ;
        RECT 2890.730 556.090 2891.910 557.270 ;
        RECT 2889.130 554.490 2890.310 555.670 ;
        RECT 2890.730 554.490 2891.910 555.670 ;
        RECT 2889.130 376.090 2890.310 377.270 ;
        RECT 2890.730 376.090 2891.910 377.270 ;
        RECT 2889.130 374.490 2890.310 375.670 ;
        RECT 2890.730 374.490 2891.910 375.670 ;
        RECT 2889.130 196.090 2890.310 197.270 ;
        RECT 2890.730 196.090 2891.910 197.270 ;
        RECT 2889.130 194.490 2890.310 195.670 ;
        RECT 2890.730 194.490 2891.910 195.670 ;
        RECT 2889.130 16.090 2890.310 17.270 ;
        RECT 2890.730 16.090 2891.910 17.270 ;
        RECT 2889.130 14.490 2890.310 15.670 ;
        RECT 2890.730 14.490 2891.910 15.670 ;
        RECT 2889.130 -2.910 2890.310 -1.730 ;
        RECT 2890.730 -2.910 2891.910 -1.730 ;
        RECT 2889.130 -4.510 2890.310 -3.330 ;
        RECT 2890.730 -4.510 2891.910 -3.330 ;
        RECT 2926.710 3523.010 2927.890 3524.190 ;
        RECT 2928.310 3523.010 2929.490 3524.190 ;
        RECT 2926.710 3521.410 2927.890 3522.590 ;
        RECT 2928.310 3521.410 2929.490 3522.590 ;
        RECT 2926.710 3436.090 2927.890 3437.270 ;
        RECT 2928.310 3436.090 2929.490 3437.270 ;
        RECT 2926.710 3434.490 2927.890 3435.670 ;
        RECT 2928.310 3434.490 2929.490 3435.670 ;
        RECT 2926.710 3256.090 2927.890 3257.270 ;
        RECT 2928.310 3256.090 2929.490 3257.270 ;
        RECT 2926.710 3254.490 2927.890 3255.670 ;
        RECT 2928.310 3254.490 2929.490 3255.670 ;
        RECT 2926.710 3076.090 2927.890 3077.270 ;
        RECT 2928.310 3076.090 2929.490 3077.270 ;
        RECT 2926.710 3074.490 2927.890 3075.670 ;
        RECT 2928.310 3074.490 2929.490 3075.670 ;
        RECT 2926.710 2896.090 2927.890 2897.270 ;
        RECT 2928.310 2896.090 2929.490 2897.270 ;
        RECT 2926.710 2894.490 2927.890 2895.670 ;
        RECT 2928.310 2894.490 2929.490 2895.670 ;
        RECT 2926.710 2716.090 2927.890 2717.270 ;
        RECT 2928.310 2716.090 2929.490 2717.270 ;
        RECT 2926.710 2714.490 2927.890 2715.670 ;
        RECT 2928.310 2714.490 2929.490 2715.670 ;
        RECT 2926.710 2536.090 2927.890 2537.270 ;
        RECT 2928.310 2536.090 2929.490 2537.270 ;
        RECT 2926.710 2534.490 2927.890 2535.670 ;
        RECT 2928.310 2534.490 2929.490 2535.670 ;
        RECT 2926.710 2356.090 2927.890 2357.270 ;
        RECT 2928.310 2356.090 2929.490 2357.270 ;
        RECT 2926.710 2354.490 2927.890 2355.670 ;
        RECT 2928.310 2354.490 2929.490 2355.670 ;
        RECT 2926.710 2176.090 2927.890 2177.270 ;
        RECT 2928.310 2176.090 2929.490 2177.270 ;
        RECT 2926.710 2174.490 2927.890 2175.670 ;
        RECT 2928.310 2174.490 2929.490 2175.670 ;
        RECT 2926.710 1996.090 2927.890 1997.270 ;
        RECT 2928.310 1996.090 2929.490 1997.270 ;
        RECT 2926.710 1994.490 2927.890 1995.670 ;
        RECT 2928.310 1994.490 2929.490 1995.670 ;
        RECT 2926.710 1816.090 2927.890 1817.270 ;
        RECT 2928.310 1816.090 2929.490 1817.270 ;
        RECT 2926.710 1814.490 2927.890 1815.670 ;
        RECT 2928.310 1814.490 2929.490 1815.670 ;
        RECT 2926.710 1636.090 2927.890 1637.270 ;
        RECT 2928.310 1636.090 2929.490 1637.270 ;
        RECT 2926.710 1634.490 2927.890 1635.670 ;
        RECT 2928.310 1634.490 2929.490 1635.670 ;
        RECT 2926.710 1456.090 2927.890 1457.270 ;
        RECT 2928.310 1456.090 2929.490 1457.270 ;
        RECT 2926.710 1454.490 2927.890 1455.670 ;
        RECT 2928.310 1454.490 2929.490 1455.670 ;
        RECT 2926.710 1276.090 2927.890 1277.270 ;
        RECT 2928.310 1276.090 2929.490 1277.270 ;
        RECT 2926.710 1274.490 2927.890 1275.670 ;
        RECT 2928.310 1274.490 2929.490 1275.670 ;
        RECT 2926.710 1096.090 2927.890 1097.270 ;
        RECT 2928.310 1096.090 2929.490 1097.270 ;
        RECT 2926.710 1094.490 2927.890 1095.670 ;
        RECT 2928.310 1094.490 2929.490 1095.670 ;
        RECT 2926.710 916.090 2927.890 917.270 ;
        RECT 2928.310 916.090 2929.490 917.270 ;
        RECT 2926.710 914.490 2927.890 915.670 ;
        RECT 2928.310 914.490 2929.490 915.670 ;
        RECT 2926.710 736.090 2927.890 737.270 ;
        RECT 2928.310 736.090 2929.490 737.270 ;
        RECT 2926.710 734.490 2927.890 735.670 ;
        RECT 2928.310 734.490 2929.490 735.670 ;
        RECT 2926.710 556.090 2927.890 557.270 ;
        RECT 2928.310 556.090 2929.490 557.270 ;
        RECT 2926.710 554.490 2927.890 555.670 ;
        RECT 2928.310 554.490 2929.490 555.670 ;
        RECT 2926.710 376.090 2927.890 377.270 ;
        RECT 2928.310 376.090 2929.490 377.270 ;
        RECT 2926.710 374.490 2927.890 375.670 ;
        RECT 2928.310 374.490 2929.490 375.670 ;
        RECT 2926.710 196.090 2927.890 197.270 ;
        RECT 2928.310 196.090 2929.490 197.270 ;
        RECT 2926.710 194.490 2927.890 195.670 ;
        RECT 2928.310 194.490 2929.490 195.670 ;
        RECT 2926.710 16.090 2927.890 17.270 ;
        RECT 2928.310 16.090 2929.490 17.270 ;
        RECT 2926.710 14.490 2927.890 15.670 ;
        RECT 2928.310 14.490 2929.490 15.670 ;
        RECT 2926.710 -2.910 2927.890 -1.730 ;
        RECT 2928.310 -2.910 2929.490 -1.730 ;
        RECT 2926.710 -4.510 2927.890 -3.330 ;
        RECT 2928.310 -4.510 2929.490 -3.330 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
        RECT -14.830 914.330 2934.450 917.430 ;
        RECT -14.830 734.330 2934.450 737.430 ;
        RECT -14.830 554.330 2934.450 557.430 ;
        RECT -14.830 374.330 2934.450 377.430 ;
        RECT -14.830 194.330 2934.450 197.430 ;
        RECT -14.830 14.330 2934.450 17.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
        RECT 207.570 1010.000 210.670 3538.750 ;
        RECT 387.570 1010.000 390.670 3538.750 ;
        RECT 567.570 1010.000 570.670 3538.750 ;
        RECT 747.570 1010.000 750.670 3538.750 ;
        RECT 927.570 1010.000 930.670 3538.750 ;
        RECT 1107.570 1010.000 1110.670 3538.750 ;
        RECT 207.570 -19.070 210.670 390.000 ;
        RECT 387.570 -19.070 390.670 390.000 ;
        RECT 567.570 -19.070 570.670 390.000 ;
        RECT 747.570 -19.070 750.670 390.000 ;
        RECT 927.570 -19.070 930.670 390.000 ;
        RECT 1107.570 -19.070 1110.670 390.000 ;
        RECT 1287.570 -19.070 1290.670 3538.750 ;
        RECT 1467.570 -19.070 1470.670 3538.750 ;
        RECT 1647.570 -19.070 1650.670 3538.750 ;
        RECT 1827.570 -19.070 1830.670 3538.750 ;
        RECT 2007.570 -19.070 2010.670 3538.750 ;
        RECT 2187.570 -19.070 2190.670 3538.750 ;
        RECT 2367.570 -19.070 2370.670 3538.750 ;
        RECT 2547.570 -19.070 2550.670 3538.750 ;
        RECT 2727.570 -19.070 2730.670 3538.750 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER via4 ;
        RECT -19.470 3532.610 -18.290 3533.790 ;
        RECT -17.870 3532.610 -16.690 3533.790 ;
        RECT -19.470 3531.010 -18.290 3532.190 ;
        RECT -17.870 3531.010 -16.690 3532.190 ;
        RECT -19.470 3454.690 -18.290 3455.870 ;
        RECT -17.870 3454.690 -16.690 3455.870 ;
        RECT -19.470 3453.090 -18.290 3454.270 ;
        RECT -17.870 3453.090 -16.690 3454.270 ;
        RECT -19.470 3274.690 -18.290 3275.870 ;
        RECT -17.870 3274.690 -16.690 3275.870 ;
        RECT -19.470 3273.090 -18.290 3274.270 ;
        RECT -17.870 3273.090 -16.690 3274.270 ;
        RECT -19.470 3094.690 -18.290 3095.870 ;
        RECT -17.870 3094.690 -16.690 3095.870 ;
        RECT -19.470 3093.090 -18.290 3094.270 ;
        RECT -17.870 3093.090 -16.690 3094.270 ;
        RECT -19.470 2914.690 -18.290 2915.870 ;
        RECT -17.870 2914.690 -16.690 2915.870 ;
        RECT -19.470 2913.090 -18.290 2914.270 ;
        RECT -17.870 2913.090 -16.690 2914.270 ;
        RECT -19.470 2734.690 -18.290 2735.870 ;
        RECT -17.870 2734.690 -16.690 2735.870 ;
        RECT -19.470 2733.090 -18.290 2734.270 ;
        RECT -17.870 2733.090 -16.690 2734.270 ;
        RECT -19.470 2554.690 -18.290 2555.870 ;
        RECT -17.870 2554.690 -16.690 2555.870 ;
        RECT -19.470 2553.090 -18.290 2554.270 ;
        RECT -17.870 2553.090 -16.690 2554.270 ;
        RECT -19.470 2374.690 -18.290 2375.870 ;
        RECT -17.870 2374.690 -16.690 2375.870 ;
        RECT -19.470 2373.090 -18.290 2374.270 ;
        RECT -17.870 2373.090 -16.690 2374.270 ;
        RECT -19.470 2194.690 -18.290 2195.870 ;
        RECT -17.870 2194.690 -16.690 2195.870 ;
        RECT -19.470 2193.090 -18.290 2194.270 ;
        RECT -17.870 2193.090 -16.690 2194.270 ;
        RECT -19.470 2014.690 -18.290 2015.870 ;
        RECT -17.870 2014.690 -16.690 2015.870 ;
        RECT -19.470 2013.090 -18.290 2014.270 ;
        RECT -17.870 2013.090 -16.690 2014.270 ;
        RECT -19.470 1834.690 -18.290 1835.870 ;
        RECT -17.870 1834.690 -16.690 1835.870 ;
        RECT -19.470 1833.090 -18.290 1834.270 ;
        RECT -17.870 1833.090 -16.690 1834.270 ;
        RECT -19.470 1654.690 -18.290 1655.870 ;
        RECT -17.870 1654.690 -16.690 1655.870 ;
        RECT -19.470 1653.090 -18.290 1654.270 ;
        RECT -17.870 1653.090 -16.690 1654.270 ;
        RECT -19.470 1474.690 -18.290 1475.870 ;
        RECT -17.870 1474.690 -16.690 1475.870 ;
        RECT -19.470 1473.090 -18.290 1474.270 ;
        RECT -17.870 1473.090 -16.690 1474.270 ;
        RECT -19.470 1294.690 -18.290 1295.870 ;
        RECT -17.870 1294.690 -16.690 1295.870 ;
        RECT -19.470 1293.090 -18.290 1294.270 ;
        RECT -17.870 1293.090 -16.690 1294.270 ;
        RECT -19.470 1114.690 -18.290 1115.870 ;
        RECT -17.870 1114.690 -16.690 1115.870 ;
        RECT -19.470 1113.090 -18.290 1114.270 ;
        RECT -17.870 1113.090 -16.690 1114.270 ;
        RECT -19.470 934.690 -18.290 935.870 ;
        RECT -17.870 934.690 -16.690 935.870 ;
        RECT -19.470 933.090 -18.290 934.270 ;
        RECT -17.870 933.090 -16.690 934.270 ;
        RECT -19.470 754.690 -18.290 755.870 ;
        RECT -17.870 754.690 -16.690 755.870 ;
        RECT -19.470 753.090 -18.290 754.270 ;
        RECT -17.870 753.090 -16.690 754.270 ;
        RECT -19.470 574.690 -18.290 575.870 ;
        RECT -17.870 574.690 -16.690 575.870 ;
        RECT -19.470 573.090 -18.290 574.270 ;
        RECT -17.870 573.090 -16.690 574.270 ;
        RECT -19.470 394.690 -18.290 395.870 ;
        RECT -17.870 394.690 -16.690 395.870 ;
        RECT -19.470 393.090 -18.290 394.270 ;
        RECT -17.870 393.090 -16.690 394.270 ;
        RECT -19.470 214.690 -18.290 215.870 ;
        RECT -17.870 214.690 -16.690 215.870 ;
        RECT -19.470 213.090 -18.290 214.270 ;
        RECT -17.870 213.090 -16.690 214.270 ;
        RECT -19.470 34.690 -18.290 35.870 ;
        RECT -17.870 34.690 -16.690 35.870 ;
        RECT -19.470 33.090 -18.290 34.270 ;
        RECT -17.870 33.090 -16.690 34.270 ;
        RECT -19.470 -12.510 -18.290 -11.330 ;
        RECT -17.870 -12.510 -16.690 -11.330 ;
        RECT -19.470 -14.110 -18.290 -12.930 ;
        RECT -17.870 -14.110 -16.690 -12.930 ;
        RECT 27.730 3532.610 28.910 3533.790 ;
        RECT 29.330 3532.610 30.510 3533.790 ;
        RECT 27.730 3531.010 28.910 3532.190 ;
        RECT 29.330 3531.010 30.510 3532.190 ;
        RECT 27.730 3454.690 28.910 3455.870 ;
        RECT 29.330 3454.690 30.510 3455.870 ;
        RECT 27.730 3453.090 28.910 3454.270 ;
        RECT 29.330 3453.090 30.510 3454.270 ;
        RECT 27.730 3274.690 28.910 3275.870 ;
        RECT 29.330 3274.690 30.510 3275.870 ;
        RECT 27.730 3273.090 28.910 3274.270 ;
        RECT 29.330 3273.090 30.510 3274.270 ;
        RECT 27.730 3094.690 28.910 3095.870 ;
        RECT 29.330 3094.690 30.510 3095.870 ;
        RECT 27.730 3093.090 28.910 3094.270 ;
        RECT 29.330 3093.090 30.510 3094.270 ;
        RECT 27.730 2914.690 28.910 2915.870 ;
        RECT 29.330 2914.690 30.510 2915.870 ;
        RECT 27.730 2913.090 28.910 2914.270 ;
        RECT 29.330 2913.090 30.510 2914.270 ;
        RECT 27.730 2734.690 28.910 2735.870 ;
        RECT 29.330 2734.690 30.510 2735.870 ;
        RECT 27.730 2733.090 28.910 2734.270 ;
        RECT 29.330 2733.090 30.510 2734.270 ;
        RECT 27.730 2554.690 28.910 2555.870 ;
        RECT 29.330 2554.690 30.510 2555.870 ;
        RECT 27.730 2553.090 28.910 2554.270 ;
        RECT 29.330 2553.090 30.510 2554.270 ;
        RECT 27.730 2374.690 28.910 2375.870 ;
        RECT 29.330 2374.690 30.510 2375.870 ;
        RECT 27.730 2373.090 28.910 2374.270 ;
        RECT 29.330 2373.090 30.510 2374.270 ;
        RECT 27.730 2194.690 28.910 2195.870 ;
        RECT 29.330 2194.690 30.510 2195.870 ;
        RECT 27.730 2193.090 28.910 2194.270 ;
        RECT 29.330 2193.090 30.510 2194.270 ;
        RECT 27.730 2014.690 28.910 2015.870 ;
        RECT 29.330 2014.690 30.510 2015.870 ;
        RECT 27.730 2013.090 28.910 2014.270 ;
        RECT 29.330 2013.090 30.510 2014.270 ;
        RECT 27.730 1834.690 28.910 1835.870 ;
        RECT 29.330 1834.690 30.510 1835.870 ;
        RECT 27.730 1833.090 28.910 1834.270 ;
        RECT 29.330 1833.090 30.510 1834.270 ;
        RECT 27.730 1654.690 28.910 1655.870 ;
        RECT 29.330 1654.690 30.510 1655.870 ;
        RECT 27.730 1653.090 28.910 1654.270 ;
        RECT 29.330 1653.090 30.510 1654.270 ;
        RECT 27.730 1474.690 28.910 1475.870 ;
        RECT 29.330 1474.690 30.510 1475.870 ;
        RECT 27.730 1473.090 28.910 1474.270 ;
        RECT 29.330 1473.090 30.510 1474.270 ;
        RECT 27.730 1294.690 28.910 1295.870 ;
        RECT 29.330 1294.690 30.510 1295.870 ;
        RECT 27.730 1293.090 28.910 1294.270 ;
        RECT 29.330 1293.090 30.510 1294.270 ;
        RECT 27.730 1114.690 28.910 1115.870 ;
        RECT 29.330 1114.690 30.510 1115.870 ;
        RECT 27.730 1113.090 28.910 1114.270 ;
        RECT 29.330 1113.090 30.510 1114.270 ;
        RECT 207.730 3532.610 208.910 3533.790 ;
        RECT 209.330 3532.610 210.510 3533.790 ;
        RECT 207.730 3531.010 208.910 3532.190 ;
        RECT 209.330 3531.010 210.510 3532.190 ;
        RECT 207.730 3454.690 208.910 3455.870 ;
        RECT 209.330 3454.690 210.510 3455.870 ;
        RECT 207.730 3453.090 208.910 3454.270 ;
        RECT 209.330 3453.090 210.510 3454.270 ;
        RECT 207.730 3274.690 208.910 3275.870 ;
        RECT 209.330 3274.690 210.510 3275.870 ;
        RECT 207.730 3273.090 208.910 3274.270 ;
        RECT 209.330 3273.090 210.510 3274.270 ;
        RECT 207.730 3094.690 208.910 3095.870 ;
        RECT 209.330 3094.690 210.510 3095.870 ;
        RECT 207.730 3093.090 208.910 3094.270 ;
        RECT 209.330 3093.090 210.510 3094.270 ;
        RECT 207.730 2914.690 208.910 2915.870 ;
        RECT 209.330 2914.690 210.510 2915.870 ;
        RECT 207.730 2913.090 208.910 2914.270 ;
        RECT 209.330 2913.090 210.510 2914.270 ;
        RECT 207.730 2734.690 208.910 2735.870 ;
        RECT 209.330 2734.690 210.510 2735.870 ;
        RECT 207.730 2733.090 208.910 2734.270 ;
        RECT 209.330 2733.090 210.510 2734.270 ;
        RECT 207.730 2554.690 208.910 2555.870 ;
        RECT 209.330 2554.690 210.510 2555.870 ;
        RECT 207.730 2553.090 208.910 2554.270 ;
        RECT 209.330 2553.090 210.510 2554.270 ;
        RECT 207.730 2374.690 208.910 2375.870 ;
        RECT 209.330 2374.690 210.510 2375.870 ;
        RECT 207.730 2373.090 208.910 2374.270 ;
        RECT 209.330 2373.090 210.510 2374.270 ;
        RECT 207.730 2194.690 208.910 2195.870 ;
        RECT 209.330 2194.690 210.510 2195.870 ;
        RECT 207.730 2193.090 208.910 2194.270 ;
        RECT 209.330 2193.090 210.510 2194.270 ;
        RECT 207.730 2014.690 208.910 2015.870 ;
        RECT 209.330 2014.690 210.510 2015.870 ;
        RECT 207.730 2013.090 208.910 2014.270 ;
        RECT 209.330 2013.090 210.510 2014.270 ;
        RECT 207.730 1834.690 208.910 1835.870 ;
        RECT 209.330 1834.690 210.510 1835.870 ;
        RECT 207.730 1833.090 208.910 1834.270 ;
        RECT 209.330 1833.090 210.510 1834.270 ;
        RECT 207.730 1654.690 208.910 1655.870 ;
        RECT 209.330 1654.690 210.510 1655.870 ;
        RECT 207.730 1653.090 208.910 1654.270 ;
        RECT 209.330 1653.090 210.510 1654.270 ;
        RECT 207.730 1474.690 208.910 1475.870 ;
        RECT 209.330 1474.690 210.510 1475.870 ;
        RECT 207.730 1473.090 208.910 1474.270 ;
        RECT 209.330 1473.090 210.510 1474.270 ;
        RECT 207.730 1294.690 208.910 1295.870 ;
        RECT 209.330 1294.690 210.510 1295.870 ;
        RECT 207.730 1293.090 208.910 1294.270 ;
        RECT 209.330 1293.090 210.510 1294.270 ;
        RECT 207.730 1114.690 208.910 1115.870 ;
        RECT 209.330 1114.690 210.510 1115.870 ;
        RECT 207.730 1113.090 208.910 1114.270 ;
        RECT 209.330 1113.090 210.510 1114.270 ;
        RECT 387.730 3532.610 388.910 3533.790 ;
        RECT 389.330 3532.610 390.510 3533.790 ;
        RECT 387.730 3531.010 388.910 3532.190 ;
        RECT 389.330 3531.010 390.510 3532.190 ;
        RECT 387.730 3454.690 388.910 3455.870 ;
        RECT 389.330 3454.690 390.510 3455.870 ;
        RECT 387.730 3453.090 388.910 3454.270 ;
        RECT 389.330 3453.090 390.510 3454.270 ;
        RECT 387.730 3274.690 388.910 3275.870 ;
        RECT 389.330 3274.690 390.510 3275.870 ;
        RECT 387.730 3273.090 388.910 3274.270 ;
        RECT 389.330 3273.090 390.510 3274.270 ;
        RECT 387.730 3094.690 388.910 3095.870 ;
        RECT 389.330 3094.690 390.510 3095.870 ;
        RECT 387.730 3093.090 388.910 3094.270 ;
        RECT 389.330 3093.090 390.510 3094.270 ;
        RECT 387.730 2914.690 388.910 2915.870 ;
        RECT 389.330 2914.690 390.510 2915.870 ;
        RECT 387.730 2913.090 388.910 2914.270 ;
        RECT 389.330 2913.090 390.510 2914.270 ;
        RECT 387.730 2734.690 388.910 2735.870 ;
        RECT 389.330 2734.690 390.510 2735.870 ;
        RECT 387.730 2733.090 388.910 2734.270 ;
        RECT 389.330 2733.090 390.510 2734.270 ;
        RECT 387.730 2554.690 388.910 2555.870 ;
        RECT 389.330 2554.690 390.510 2555.870 ;
        RECT 387.730 2553.090 388.910 2554.270 ;
        RECT 389.330 2553.090 390.510 2554.270 ;
        RECT 387.730 2374.690 388.910 2375.870 ;
        RECT 389.330 2374.690 390.510 2375.870 ;
        RECT 387.730 2373.090 388.910 2374.270 ;
        RECT 389.330 2373.090 390.510 2374.270 ;
        RECT 387.730 2194.690 388.910 2195.870 ;
        RECT 389.330 2194.690 390.510 2195.870 ;
        RECT 387.730 2193.090 388.910 2194.270 ;
        RECT 389.330 2193.090 390.510 2194.270 ;
        RECT 387.730 2014.690 388.910 2015.870 ;
        RECT 389.330 2014.690 390.510 2015.870 ;
        RECT 387.730 2013.090 388.910 2014.270 ;
        RECT 389.330 2013.090 390.510 2014.270 ;
        RECT 387.730 1834.690 388.910 1835.870 ;
        RECT 389.330 1834.690 390.510 1835.870 ;
        RECT 387.730 1833.090 388.910 1834.270 ;
        RECT 389.330 1833.090 390.510 1834.270 ;
        RECT 387.730 1654.690 388.910 1655.870 ;
        RECT 389.330 1654.690 390.510 1655.870 ;
        RECT 387.730 1653.090 388.910 1654.270 ;
        RECT 389.330 1653.090 390.510 1654.270 ;
        RECT 387.730 1474.690 388.910 1475.870 ;
        RECT 389.330 1474.690 390.510 1475.870 ;
        RECT 387.730 1473.090 388.910 1474.270 ;
        RECT 389.330 1473.090 390.510 1474.270 ;
        RECT 387.730 1294.690 388.910 1295.870 ;
        RECT 389.330 1294.690 390.510 1295.870 ;
        RECT 387.730 1293.090 388.910 1294.270 ;
        RECT 389.330 1293.090 390.510 1294.270 ;
        RECT 387.730 1114.690 388.910 1115.870 ;
        RECT 389.330 1114.690 390.510 1115.870 ;
        RECT 387.730 1113.090 388.910 1114.270 ;
        RECT 389.330 1113.090 390.510 1114.270 ;
        RECT 567.730 3532.610 568.910 3533.790 ;
        RECT 569.330 3532.610 570.510 3533.790 ;
        RECT 567.730 3531.010 568.910 3532.190 ;
        RECT 569.330 3531.010 570.510 3532.190 ;
        RECT 567.730 3454.690 568.910 3455.870 ;
        RECT 569.330 3454.690 570.510 3455.870 ;
        RECT 567.730 3453.090 568.910 3454.270 ;
        RECT 569.330 3453.090 570.510 3454.270 ;
        RECT 567.730 3274.690 568.910 3275.870 ;
        RECT 569.330 3274.690 570.510 3275.870 ;
        RECT 567.730 3273.090 568.910 3274.270 ;
        RECT 569.330 3273.090 570.510 3274.270 ;
        RECT 567.730 3094.690 568.910 3095.870 ;
        RECT 569.330 3094.690 570.510 3095.870 ;
        RECT 567.730 3093.090 568.910 3094.270 ;
        RECT 569.330 3093.090 570.510 3094.270 ;
        RECT 567.730 2914.690 568.910 2915.870 ;
        RECT 569.330 2914.690 570.510 2915.870 ;
        RECT 567.730 2913.090 568.910 2914.270 ;
        RECT 569.330 2913.090 570.510 2914.270 ;
        RECT 567.730 2734.690 568.910 2735.870 ;
        RECT 569.330 2734.690 570.510 2735.870 ;
        RECT 567.730 2733.090 568.910 2734.270 ;
        RECT 569.330 2733.090 570.510 2734.270 ;
        RECT 567.730 2554.690 568.910 2555.870 ;
        RECT 569.330 2554.690 570.510 2555.870 ;
        RECT 567.730 2553.090 568.910 2554.270 ;
        RECT 569.330 2553.090 570.510 2554.270 ;
        RECT 567.730 2374.690 568.910 2375.870 ;
        RECT 569.330 2374.690 570.510 2375.870 ;
        RECT 567.730 2373.090 568.910 2374.270 ;
        RECT 569.330 2373.090 570.510 2374.270 ;
        RECT 567.730 2194.690 568.910 2195.870 ;
        RECT 569.330 2194.690 570.510 2195.870 ;
        RECT 567.730 2193.090 568.910 2194.270 ;
        RECT 569.330 2193.090 570.510 2194.270 ;
        RECT 567.730 2014.690 568.910 2015.870 ;
        RECT 569.330 2014.690 570.510 2015.870 ;
        RECT 567.730 2013.090 568.910 2014.270 ;
        RECT 569.330 2013.090 570.510 2014.270 ;
        RECT 567.730 1834.690 568.910 1835.870 ;
        RECT 569.330 1834.690 570.510 1835.870 ;
        RECT 567.730 1833.090 568.910 1834.270 ;
        RECT 569.330 1833.090 570.510 1834.270 ;
        RECT 567.730 1654.690 568.910 1655.870 ;
        RECT 569.330 1654.690 570.510 1655.870 ;
        RECT 567.730 1653.090 568.910 1654.270 ;
        RECT 569.330 1653.090 570.510 1654.270 ;
        RECT 567.730 1474.690 568.910 1475.870 ;
        RECT 569.330 1474.690 570.510 1475.870 ;
        RECT 567.730 1473.090 568.910 1474.270 ;
        RECT 569.330 1473.090 570.510 1474.270 ;
        RECT 567.730 1294.690 568.910 1295.870 ;
        RECT 569.330 1294.690 570.510 1295.870 ;
        RECT 567.730 1293.090 568.910 1294.270 ;
        RECT 569.330 1293.090 570.510 1294.270 ;
        RECT 567.730 1114.690 568.910 1115.870 ;
        RECT 569.330 1114.690 570.510 1115.870 ;
        RECT 567.730 1113.090 568.910 1114.270 ;
        RECT 569.330 1113.090 570.510 1114.270 ;
        RECT 747.730 3532.610 748.910 3533.790 ;
        RECT 749.330 3532.610 750.510 3533.790 ;
        RECT 747.730 3531.010 748.910 3532.190 ;
        RECT 749.330 3531.010 750.510 3532.190 ;
        RECT 747.730 3454.690 748.910 3455.870 ;
        RECT 749.330 3454.690 750.510 3455.870 ;
        RECT 747.730 3453.090 748.910 3454.270 ;
        RECT 749.330 3453.090 750.510 3454.270 ;
        RECT 747.730 3274.690 748.910 3275.870 ;
        RECT 749.330 3274.690 750.510 3275.870 ;
        RECT 747.730 3273.090 748.910 3274.270 ;
        RECT 749.330 3273.090 750.510 3274.270 ;
        RECT 747.730 3094.690 748.910 3095.870 ;
        RECT 749.330 3094.690 750.510 3095.870 ;
        RECT 747.730 3093.090 748.910 3094.270 ;
        RECT 749.330 3093.090 750.510 3094.270 ;
        RECT 747.730 2914.690 748.910 2915.870 ;
        RECT 749.330 2914.690 750.510 2915.870 ;
        RECT 747.730 2913.090 748.910 2914.270 ;
        RECT 749.330 2913.090 750.510 2914.270 ;
        RECT 747.730 2734.690 748.910 2735.870 ;
        RECT 749.330 2734.690 750.510 2735.870 ;
        RECT 747.730 2733.090 748.910 2734.270 ;
        RECT 749.330 2733.090 750.510 2734.270 ;
        RECT 747.730 2554.690 748.910 2555.870 ;
        RECT 749.330 2554.690 750.510 2555.870 ;
        RECT 747.730 2553.090 748.910 2554.270 ;
        RECT 749.330 2553.090 750.510 2554.270 ;
        RECT 747.730 2374.690 748.910 2375.870 ;
        RECT 749.330 2374.690 750.510 2375.870 ;
        RECT 747.730 2373.090 748.910 2374.270 ;
        RECT 749.330 2373.090 750.510 2374.270 ;
        RECT 747.730 2194.690 748.910 2195.870 ;
        RECT 749.330 2194.690 750.510 2195.870 ;
        RECT 747.730 2193.090 748.910 2194.270 ;
        RECT 749.330 2193.090 750.510 2194.270 ;
        RECT 747.730 2014.690 748.910 2015.870 ;
        RECT 749.330 2014.690 750.510 2015.870 ;
        RECT 747.730 2013.090 748.910 2014.270 ;
        RECT 749.330 2013.090 750.510 2014.270 ;
        RECT 747.730 1834.690 748.910 1835.870 ;
        RECT 749.330 1834.690 750.510 1835.870 ;
        RECT 747.730 1833.090 748.910 1834.270 ;
        RECT 749.330 1833.090 750.510 1834.270 ;
        RECT 747.730 1654.690 748.910 1655.870 ;
        RECT 749.330 1654.690 750.510 1655.870 ;
        RECT 747.730 1653.090 748.910 1654.270 ;
        RECT 749.330 1653.090 750.510 1654.270 ;
        RECT 747.730 1474.690 748.910 1475.870 ;
        RECT 749.330 1474.690 750.510 1475.870 ;
        RECT 747.730 1473.090 748.910 1474.270 ;
        RECT 749.330 1473.090 750.510 1474.270 ;
        RECT 747.730 1294.690 748.910 1295.870 ;
        RECT 749.330 1294.690 750.510 1295.870 ;
        RECT 747.730 1293.090 748.910 1294.270 ;
        RECT 749.330 1293.090 750.510 1294.270 ;
        RECT 747.730 1114.690 748.910 1115.870 ;
        RECT 749.330 1114.690 750.510 1115.870 ;
        RECT 747.730 1113.090 748.910 1114.270 ;
        RECT 749.330 1113.090 750.510 1114.270 ;
        RECT 927.730 3532.610 928.910 3533.790 ;
        RECT 929.330 3532.610 930.510 3533.790 ;
        RECT 927.730 3531.010 928.910 3532.190 ;
        RECT 929.330 3531.010 930.510 3532.190 ;
        RECT 927.730 3454.690 928.910 3455.870 ;
        RECT 929.330 3454.690 930.510 3455.870 ;
        RECT 927.730 3453.090 928.910 3454.270 ;
        RECT 929.330 3453.090 930.510 3454.270 ;
        RECT 927.730 3274.690 928.910 3275.870 ;
        RECT 929.330 3274.690 930.510 3275.870 ;
        RECT 927.730 3273.090 928.910 3274.270 ;
        RECT 929.330 3273.090 930.510 3274.270 ;
        RECT 927.730 3094.690 928.910 3095.870 ;
        RECT 929.330 3094.690 930.510 3095.870 ;
        RECT 927.730 3093.090 928.910 3094.270 ;
        RECT 929.330 3093.090 930.510 3094.270 ;
        RECT 927.730 2914.690 928.910 2915.870 ;
        RECT 929.330 2914.690 930.510 2915.870 ;
        RECT 927.730 2913.090 928.910 2914.270 ;
        RECT 929.330 2913.090 930.510 2914.270 ;
        RECT 927.730 2734.690 928.910 2735.870 ;
        RECT 929.330 2734.690 930.510 2735.870 ;
        RECT 927.730 2733.090 928.910 2734.270 ;
        RECT 929.330 2733.090 930.510 2734.270 ;
        RECT 927.730 2554.690 928.910 2555.870 ;
        RECT 929.330 2554.690 930.510 2555.870 ;
        RECT 927.730 2553.090 928.910 2554.270 ;
        RECT 929.330 2553.090 930.510 2554.270 ;
        RECT 927.730 2374.690 928.910 2375.870 ;
        RECT 929.330 2374.690 930.510 2375.870 ;
        RECT 927.730 2373.090 928.910 2374.270 ;
        RECT 929.330 2373.090 930.510 2374.270 ;
        RECT 927.730 2194.690 928.910 2195.870 ;
        RECT 929.330 2194.690 930.510 2195.870 ;
        RECT 927.730 2193.090 928.910 2194.270 ;
        RECT 929.330 2193.090 930.510 2194.270 ;
        RECT 927.730 2014.690 928.910 2015.870 ;
        RECT 929.330 2014.690 930.510 2015.870 ;
        RECT 927.730 2013.090 928.910 2014.270 ;
        RECT 929.330 2013.090 930.510 2014.270 ;
        RECT 927.730 1834.690 928.910 1835.870 ;
        RECT 929.330 1834.690 930.510 1835.870 ;
        RECT 927.730 1833.090 928.910 1834.270 ;
        RECT 929.330 1833.090 930.510 1834.270 ;
        RECT 927.730 1654.690 928.910 1655.870 ;
        RECT 929.330 1654.690 930.510 1655.870 ;
        RECT 927.730 1653.090 928.910 1654.270 ;
        RECT 929.330 1653.090 930.510 1654.270 ;
        RECT 927.730 1474.690 928.910 1475.870 ;
        RECT 929.330 1474.690 930.510 1475.870 ;
        RECT 927.730 1473.090 928.910 1474.270 ;
        RECT 929.330 1473.090 930.510 1474.270 ;
        RECT 927.730 1294.690 928.910 1295.870 ;
        RECT 929.330 1294.690 930.510 1295.870 ;
        RECT 927.730 1293.090 928.910 1294.270 ;
        RECT 929.330 1293.090 930.510 1294.270 ;
        RECT 927.730 1114.690 928.910 1115.870 ;
        RECT 929.330 1114.690 930.510 1115.870 ;
        RECT 927.730 1113.090 928.910 1114.270 ;
        RECT 929.330 1113.090 930.510 1114.270 ;
        RECT 1107.730 3532.610 1108.910 3533.790 ;
        RECT 1109.330 3532.610 1110.510 3533.790 ;
        RECT 1107.730 3531.010 1108.910 3532.190 ;
        RECT 1109.330 3531.010 1110.510 3532.190 ;
        RECT 1107.730 3454.690 1108.910 3455.870 ;
        RECT 1109.330 3454.690 1110.510 3455.870 ;
        RECT 1107.730 3453.090 1108.910 3454.270 ;
        RECT 1109.330 3453.090 1110.510 3454.270 ;
        RECT 1107.730 3274.690 1108.910 3275.870 ;
        RECT 1109.330 3274.690 1110.510 3275.870 ;
        RECT 1107.730 3273.090 1108.910 3274.270 ;
        RECT 1109.330 3273.090 1110.510 3274.270 ;
        RECT 1107.730 3094.690 1108.910 3095.870 ;
        RECT 1109.330 3094.690 1110.510 3095.870 ;
        RECT 1107.730 3093.090 1108.910 3094.270 ;
        RECT 1109.330 3093.090 1110.510 3094.270 ;
        RECT 1107.730 2914.690 1108.910 2915.870 ;
        RECT 1109.330 2914.690 1110.510 2915.870 ;
        RECT 1107.730 2913.090 1108.910 2914.270 ;
        RECT 1109.330 2913.090 1110.510 2914.270 ;
        RECT 1107.730 2734.690 1108.910 2735.870 ;
        RECT 1109.330 2734.690 1110.510 2735.870 ;
        RECT 1107.730 2733.090 1108.910 2734.270 ;
        RECT 1109.330 2733.090 1110.510 2734.270 ;
        RECT 1107.730 2554.690 1108.910 2555.870 ;
        RECT 1109.330 2554.690 1110.510 2555.870 ;
        RECT 1107.730 2553.090 1108.910 2554.270 ;
        RECT 1109.330 2553.090 1110.510 2554.270 ;
        RECT 1107.730 2374.690 1108.910 2375.870 ;
        RECT 1109.330 2374.690 1110.510 2375.870 ;
        RECT 1107.730 2373.090 1108.910 2374.270 ;
        RECT 1109.330 2373.090 1110.510 2374.270 ;
        RECT 1107.730 2194.690 1108.910 2195.870 ;
        RECT 1109.330 2194.690 1110.510 2195.870 ;
        RECT 1107.730 2193.090 1108.910 2194.270 ;
        RECT 1109.330 2193.090 1110.510 2194.270 ;
        RECT 1107.730 2014.690 1108.910 2015.870 ;
        RECT 1109.330 2014.690 1110.510 2015.870 ;
        RECT 1107.730 2013.090 1108.910 2014.270 ;
        RECT 1109.330 2013.090 1110.510 2014.270 ;
        RECT 1107.730 1834.690 1108.910 1835.870 ;
        RECT 1109.330 1834.690 1110.510 1835.870 ;
        RECT 1107.730 1833.090 1108.910 1834.270 ;
        RECT 1109.330 1833.090 1110.510 1834.270 ;
        RECT 1107.730 1654.690 1108.910 1655.870 ;
        RECT 1109.330 1654.690 1110.510 1655.870 ;
        RECT 1107.730 1653.090 1108.910 1654.270 ;
        RECT 1109.330 1653.090 1110.510 1654.270 ;
        RECT 1107.730 1474.690 1108.910 1475.870 ;
        RECT 1109.330 1474.690 1110.510 1475.870 ;
        RECT 1107.730 1473.090 1108.910 1474.270 ;
        RECT 1109.330 1473.090 1110.510 1474.270 ;
        RECT 1107.730 1294.690 1108.910 1295.870 ;
        RECT 1109.330 1294.690 1110.510 1295.870 ;
        RECT 1107.730 1293.090 1108.910 1294.270 ;
        RECT 1109.330 1293.090 1110.510 1294.270 ;
        RECT 1107.730 1114.690 1108.910 1115.870 ;
        RECT 1109.330 1114.690 1110.510 1115.870 ;
        RECT 1107.730 1113.090 1108.910 1114.270 ;
        RECT 1109.330 1113.090 1110.510 1114.270 ;
        RECT 1287.730 3532.610 1288.910 3533.790 ;
        RECT 1289.330 3532.610 1290.510 3533.790 ;
        RECT 1287.730 3531.010 1288.910 3532.190 ;
        RECT 1289.330 3531.010 1290.510 3532.190 ;
        RECT 1287.730 3454.690 1288.910 3455.870 ;
        RECT 1289.330 3454.690 1290.510 3455.870 ;
        RECT 1287.730 3453.090 1288.910 3454.270 ;
        RECT 1289.330 3453.090 1290.510 3454.270 ;
        RECT 1287.730 3274.690 1288.910 3275.870 ;
        RECT 1289.330 3274.690 1290.510 3275.870 ;
        RECT 1287.730 3273.090 1288.910 3274.270 ;
        RECT 1289.330 3273.090 1290.510 3274.270 ;
        RECT 1287.730 3094.690 1288.910 3095.870 ;
        RECT 1289.330 3094.690 1290.510 3095.870 ;
        RECT 1287.730 3093.090 1288.910 3094.270 ;
        RECT 1289.330 3093.090 1290.510 3094.270 ;
        RECT 1287.730 2914.690 1288.910 2915.870 ;
        RECT 1289.330 2914.690 1290.510 2915.870 ;
        RECT 1287.730 2913.090 1288.910 2914.270 ;
        RECT 1289.330 2913.090 1290.510 2914.270 ;
        RECT 1287.730 2734.690 1288.910 2735.870 ;
        RECT 1289.330 2734.690 1290.510 2735.870 ;
        RECT 1287.730 2733.090 1288.910 2734.270 ;
        RECT 1289.330 2733.090 1290.510 2734.270 ;
        RECT 1287.730 2554.690 1288.910 2555.870 ;
        RECT 1289.330 2554.690 1290.510 2555.870 ;
        RECT 1287.730 2553.090 1288.910 2554.270 ;
        RECT 1289.330 2553.090 1290.510 2554.270 ;
        RECT 1287.730 2374.690 1288.910 2375.870 ;
        RECT 1289.330 2374.690 1290.510 2375.870 ;
        RECT 1287.730 2373.090 1288.910 2374.270 ;
        RECT 1289.330 2373.090 1290.510 2374.270 ;
        RECT 1287.730 2194.690 1288.910 2195.870 ;
        RECT 1289.330 2194.690 1290.510 2195.870 ;
        RECT 1287.730 2193.090 1288.910 2194.270 ;
        RECT 1289.330 2193.090 1290.510 2194.270 ;
        RECT 1287.730 2014.690 1288.910 2015.870 ;
        RECT 1289.330 2014.690 1290.510 2015.870 ;
        RECT 1287.730 2013.090 1288.910 2014.270 ;
        RECT 1289.330 2013.090 1290.510 2014.270 ;
        RECT 1287.730 1834.690 1288.910 1835.870 ;
        RECT 1289.330 1834.690 1290.510 1835.870 ;
        RECT 1287.730 1833.090 1288.910 1834.270 ;
        RECT 1289.330 1833.090 1290.510 1834.270 ;
        RECT 1287.730 1654.690 1288.910 1655.870 ;
        RECT 1289.330 1654.690 1290.510 1655.870 ;
        RECT 1287.730 1653.090 1288.910 1654.270 ;
        RECT 1289.330 1653.090 1290.510 1654.270 ;
        RECT 1287.730 1474.690 1288.910 1475.870 ;
        RECT 1289.330 1474.690 1290.510 1475.870 ;
        RECT 1287.730 1473.090 1288.910 1474.270 ;
        RECT 1289.330 1473.090 1290.510 1474.270 ;
        RECT 1287.730 1294.690 1288.910 1295.870 ;
        RECT 1289.330 1294.690 1290.510 1295.870 ;
        RECT 1287.730 1293.090 1288.910 1294.270 ;
        RECT 1289.330 1293.090 1290.510 1294.270 ;
        RECT 1287.730 1114.690 1288.910 1115.870 ;
        RECT 1289.330 1114.690 1290.510 1115.870 ;
        RECT 1287.730 1113.090 1288.910 1114.270 ;
        RECT 1289.330 1113.090 1290.510 1114.270 ;
        RECT 27.730 934.690 28.910 935.870 ;
        RECT 29.330 934.690 30.510 935.870 ;
        RECT 27.730 933.090 28.910 934.270 ;
        RECT 29.330 933.090 30.510 934.270 ;
        RECT 27.730 754.690 28.910 755.870 ;
        RECT 29.330 754.690 30.510 755.870 ;
        RECT 27.730 753.090 28.910 754.270 ;
        RECT 29.330 753.090 30.510 754.270 ;
        RECT 27.730 574.690 28.910 575.870 ;
        RECT 29.330 574.690 30.510 575.870 ;
        RECT 27.730 573.090 28.910 574.270 ;
        RECT 29.330 573.090 30.510 574.270 ;
        RECT 27.730 394.690 28.910 395.870 ;
        RECT 29.330 394.690 30.510 395.870 ;
        RECT 27.730 393.090 28.910 394.270 ;
        RECT 29.330 393.090 30.510 394.270 ;
        RECT 1287.730 934.690 1288.910 935.870 ;
        RECT 1289.330 934.690 1290.510 935.870 ;
        RECT 1287.730 933.090 1288.910 934.270 ;
        RECT 1289.330 933.090 1290.510 934.270 ;
        RECT 1287.730 754.690 1288.910 755.870 ;
        RECT 1289.330 754.690 1290.510 755.870 ;
        RECT 1287.730 753.090 1288.910 754.270 ;
        RECT 1289.330 753.090 1290.510 754.270 ;
        RECT 1287.730 574.690 1288.910 575.870 ;
        RECT 1289.330 574.690 1290.510 575.870 ;
        RECT 1287.730 573.090 1288.910 574.270 ;
        RECT 1289.330 573.090 1290.510 574.270 ;
        RECT 1287.730 394.690 1288.910 395.870 ;
        RECT 1289.330 394.690 1290.510 395.870 ;
        RECT 1287.730 393.090 1288.910 394.270 ;
        RECT 1289.330 393.090 1290.510 394.270 ;
        RECT 27.730 214.690 28.910 215.870 ;
        RECT 29.330 214.690 30.510 215.870 ;
        RECT 27.730 213.090 28.910 214.270 ;
        RECT 29.330 213.090 30.510 214.270 ;
        RECT 27.730 34.690 28.910 35.870 ;
        RECT 29.330 34.690 30.510 35.870 ;
        RECT 27.730 33.090 28.910 34.270 ;
        RECT 29.330 33.090 30.510 34.270 ;
        RECT 27.730 -12.510 28.910 -11.330 ;
        RECT 29.330 -12.510 30.510 -11.330 ;
        RECT 27.730 -14.110 28.910 -12.930 ;
        RECT 29.330 -14.110 30.510 -12.930 ;
        RECT 207.730 214.690 208.910 215.870 ;
        RECT 209.330 214.690 210.510 215.870 ;
        RECT 207.730 213.090 208.910 214.270 ;
        RECT 209.330 213.090 210.510 214.270 ;
        RECT 207.730 34.690 208.910 35.870 ;
        RECT 209.330 34.690 210.510 35.870 ;
        RECT 207.730 33.090 208.910 34.270 ;
        RECT 209.330 33.090 210.510 34.270 ;
        RECT 207.730 -12.510 208.910 -11.330 ;
        RECT 209.330 -12.510 210.510 -11.330 ;
        RECT 207.730 -14.110 208.910 -12.930 ;
        RECT 209.330 -14.110 210.510 -12.930 ;
        RECT 387.730 214.690 388.910 215.870 ;
        RECT 389.330 214.690 390.510 215.870 ;
        RECT 387.730 213.090 388.910 214.270 ;
        RECT 389.330 213.090 390.510 214.270 ;
        RECT 387.730 34.690 388.910 35.870 ;
        RECT 389.330 34.690 390.510 35.870 ;
        RECT 387.730 33.090 388.910 34.270 ;
        RECT 389.330 33.090 390.510 34.270 ;
        RECT 387.730 -12.510 388.910 -11.330 ;
        RECT 389.330 -12.510 390.510 -11.330 ;
        RECT 387.730 -14.110 388.910 -12.930 ;
        RECT 389.330 -14.110 390.510 -12.930 ;
        RECT 567.730 214.690 568.910 215.870 ;
        RECT 569.330 214.690 570.510 215.870 ;
        RECT 567.730 213.090 568.910 214.270 ;
        RECT 569.330 213.090 570.510 214.270 ;
        RECT 567.730 34.690 568.910 35.870 ;
        RECT 569.330 34.690 570.510 35.870 ;
        RECT 567.730 33.090 568.910 34.270 ;
        RECT 569.330 33.090 570.510 34.270 ;
        RECT 567.730 -12.510 568.910 -11.330 ;
        RECT 569.330 -12.510 570.510 -11.330 ;
        RECT 567.730 -14.110 568.910 -12.930 ;
        RECT 569.330 -14.110 570.510 -12.930 ;
        RECT 747.730 214.690 748.910 215.870 ;
        RECT 749.330 214.690 750.510 215.870 ;
        RECT 747.730 213.090 748.910 214.270 ;
        RECT 749.330 213.090 750.510 214.270 ;
        RECT 747.730 34.690 748.910 35.870 ;
        RECT 749.330 34.690 750.510 35.870 ;
        RECT 747.730 33.090 748.910 34.270 ;
        RECT 749.330 33.090 750.510 34.270 ;
        RECT 747.730 -12.510 748.910 -11.330 ;
        RECT 749.330 -12.510 750.510 -11.330 ;
        RECT 747.730 -14.110 748.910 -12.930 ;
        RECT 749.330 -14.110 750.510 -12.930 ;
        RECT 927.730 214.690 928.910 215.870 ;
        RECT 929.330 214.690 930.510 215.870 ;
        RECT 927.730 213.090 928.910 214.270 ;
        RECT 929.330 213.090 930.510 214.270 ;
        RECT 927.730 34.690 928.910 35.870 ;
        RECT 929.330 34.690 930.510 35.870 ;
        RECT 927.730 33.090 928.910 34.270 ;
        RECT 929.330 33.090 930.510 34.270 ;
        RECT 927.730 -12.510 928.910 -11.330 ;
        RECT 929.330 -12.510 930.510 -11.330 ;
        RECT 927.730 -14.110 928.910 -12.930 ;
        RECT 929.330 -14.110 930.510 -12.930 ;
        RECT 1107.730 214.690 1108.910 215.870 ;
        RECT 1109.330 214.690 1110.510 215.870 ;
        RECT 1107.730 213.090 1108.910 214.270 ;
        RECT 1109.330 213.090 1110.510 214.270 ;
        RECT 1107.730 34.690 1108.910 35.870 ;
        RECT 1109.330 34.690 1110.510 35.870 ;
        RECT 1107.730 33.090 1108.910 34.270 ;
        RECT 1109.330 33.090 1110.510 34.270 ;
        RECT 1107.730 -12.510 1108.910 -11.330 ;
        RECT 1109.330 -12.510 1110.510 -11.330 ;
        RECT 1107.730 -14.110 1108.910 -12.930 ;
        RECT 1109.330 -14.110 1110.510 -12.930 ;
        RECT 1287.730 214.690 1288.910 215.870 ;
        RECT 1289.330 214.690 1290.510 215.870 ;
        RECT 1287.730 213.090 1288.910 214.270 ;
        RECT 1289.330 213.090 1290.510 214.270 ;
        RECT 1287.730 34.690 1288.910 35.870 ;
        RECT 1289.330 34.690 1290.510 35.870 ;
        RECT 1287.730 33.090 1288.910 34.270 ;
        RECT 1289.330 33.090 1290.510 34.270 ;
        RECT 1287.730 -12.510 1288.910 -11.330 ;
        RECT 1289.330 -12.510 1290.510 -11.330 ;
        RECT 1287.730 -14.110 1288.910 -12.930 ;
        RECT 1289.330 -14.110 1290.510 -12.930 ;
        RECT 1467.730 3532.610 1468.910 3533.790 ;
        RECT 1469.330 3532.610 1470.510 3533.790 ;
        RECT 1467.730 3531.010 1468.910 3532.190 ;
        RECT 1469.330 3531.010 1470.510 3532.190 ;
        RECT 1467.730 3454.690 1468.910 3455.870 ;
        RECT 1469.330 3454.690 1470.510 3455.870 ;
        RECT 1467.730 3453.090 1468.910 3454.270 ;
        RECT 1469.330 3453.090 1470.510 3454.270 ;
        RECT 1467.730 3274.690 1468.910 3275.870 ;
        RECT 1469.330 3274.690 1470.510 3275.870 ;
        RECT 1467.730 3273.090 1468.910 3274.270 ;
        RECT 1469.330 3273.090 1470.510 3274.270 ;
        RECT 1467.730 3094.690 1468.910 3095.870 ;
        RECT 1469.330 3094.690 1470.510 3095.870 ;
        RECT 1467.730 3093.090 1468.910 3094.270 ;
        RECT 1469.330 3093.090 1470.510 3094.270 ;
        RECT 1467.730 2914.690 1468.910 2915.870 ;
        RECT 1469.330 2914.690 1470.510 2915.870 ;
        RECT 1467.730 2913.090 1468.910 2914.270 ;
        RECT 1469.330 2913.090 1470.510 2914.270 ;
        RECT 1467.730 2734.690 1468.910 2735.870 ;
        RECT 1469.330 2734.690 1470.510 2735.870 ;
        RECT 1467.730 2733.090 1468.910 2734.270 ;
        RECT 1469.330 2733.090 1470.510 2734.270 ;
        RECT 1467.730 2554.690 1468.910 2555.870 ;
        RECT 1469.330 2554.690 1470.510 2555.870 ;
        RECT 1467.730 2553.090 1468.910 2554.270 ;
        RECT 1469.330 2553.090 1470.510 2554.270 ;
        RECT 1467.730 2374.690 1468.910 2375.870 ;
        RECT 1469.330 2374.690 1470.510 2375.870 ;
        RECT 1467.730 2373.090 1468.910 2374.270 ;
        RECT 1469.330 2373.090 1470.510 2374.270 ;
        RECT 1467.730 2194.690 1468.910 2195.870 ;
        RECT 1469.330 2194.690 1470.510 2195.870 ;
        RECT 1467.730 2193.090 1468.910 2194.270 ;
        RECT 1469.330 2193.090 1470.510 2194.270 ;
        RECT 1467.730 2014.690 1468.910 2015.870 ;
        RECT 1469.330 2014.690 1470.510 2015.870 ;
        RECT 1467.730 2013.090 1468.910 2014.270 ;
        RECT 1469.330 2013.090 1470.510 2014.270 ;
        RECT 1467.730 1834.690 1468.910 1835.870 ;
        RECT 1469.330 1834.690 1470.510 1835.870 ;
        RECT 1467.730 1833.090 1468.910 1834.270 ;
        RECT 1469.330 1833.090 1470.510 1834.270 ;
        RECT 1467.730 1654.690 1468.910 1655.870 ;
        RECT 1469.330 1654.690 1470.510 1655.870 ;
        RECT 1467.730 1653.090 1468.910 1654.270 ;
        RECT 1469.330 1653.090 1470.510 1654.270 ;
        RECT 1467.730 1474.690 1468.910 1475.870 ;
        RECT 1469.330 1474.690 1470.510 1475.870 ;
        RECT 1467.730 1473.090 1468.910 1474.270 ;
        RECT 1469.330 1473.090 1470.510 1474.270 ;
        RECT 1467.730 1294.690 1468.910 1295.870 ;
        RECT 1469.330 1294.690 1470.510 1295.870 ;
        RECT 1467.730 1293.090 1468.910 1294.270 ;
        RECT 1469.330 1293.090 1470.510 1294.270 ;
        RECT 1467.730 1114.690 1468.910 1115.870 ;
        RECT 1469.330 1114.690 1470.510 1115.870 ;
        RECT 1467.730 1113.090 1468.910 1114.270 ;
        RECT 1469.330 1113.090 1470.510 1114.270 ;
        RECT 1467.730 934.690 1468.910 935.870 ;
        RECT 1469.330 934.690 1470.510 935.870 ;
        RECT 1467.730 933.090 1468.910 934.270 ;
        RECT 1469.330 933.090 1470.510 934.270 ;
        RECT 1467.730 754.690 1468.910 755.870 ;
        RECT 1469.330 754.690 1470.510 755.870 ;
        RECT 1467.730 753.090 1468.910 754.270 ;
        RECT 1469.330 753.090 1470.510 754.270 ;
        RECT 1467.730 574.690 1468.910 575.870 ;
        RECT 1469.330 574.690 1470.510 575.870 ;
        RECT 1467.730 573.090 1468.910 574.270 ;
        RECT 1469.330 573.090 1470.510 574.270 ;
        RECT 1467.730 394.690 1468.910 395.870 ;
        RECT 1469.330 394.690 1470.510 395.870 ;
        RECT 1467.730 393.090 1468.910 394.270 ;
        RECT 1469.330 393.090 1470.510 394.270 ;
        RECT 1467.730 214.690 1468.910 215.870 ;
        RECT 1469.330 214.690 1470.510 215.870 ;
        RECT 1467.730 213.090 1468.910 214.270 ;
        RECT 1469.330 213.090 1470.510 214.270 ;
        RECT 1467.730 34.690 1468.910 35.870 ;
        RECT 1469.330 34.690 1470.510 35.870 ;
        RECT 1467.730 33.090 1468.910 34.270 ;
        RECT 1469.330 33.090 1470.510 34.270 ;
        RECT 1467.730 -12.510 1468.910 -11.330 ;
        RECT 1469.330 -12.510 1470.510 -11.330 ;
        RECT 1467.730 -14.110 1468.910 -12.930 ;
        RECT 1469.330 -14.110 1470.510 -12.930 ;
        RECT 1647.730 3532.610 1648.910 3533.790 ;
        RECT 1649.330 3532.610 1650.510 3533.790 ;
        RECT 1647.730 3531.010 1648.910 3532.190 ;
        RECT 1649.330 3531.010 1650.510 3532.190 ;
        RECT 1647.730 3454.690 1648.910 3455.870 ;
        RECT 1649.330 3454.690 1650.510 3455.870 ;
        RECT 1647.730 3453.090 1648.910 3454.270 ;
        RECT 1649.330 3453.090 1650.510 3454.270 ;
        RECT 1647.730 3274.690 1648.910 3275.870 ;
        RECT 1649.330 3274.690 1650.510 3275.870 ;
        RECT 1647.730 3273.090 1648.910 3274.270 ;
        RECT 1649.330 3273.090 1650.510 3274.270 ;
        RECT 1647.730 3094.690 1648.910 3095.870 ;
        RECT 1649.330 3094.690 1650.510 3095.870 ;
        RECT 1647.730 3093.090 1648.910 3094.270 ;
        RECT 1649.330 3093.090 1650.510 3094.270 ;
        RECT 1647.730 2914.690 1648.910 2915.870 ;
        RECT 1649.330 2914.690 1650.510 2915.870 ;
        RECT 1647.730 2913.090 1648.910 2914.270 ;
        RECT 1649.330 2913.090 1650.510 2914.270 ;
        RECT 1647.730 2734.690 1648.910 2735.870 ;
        RECT 1649.330 2734.690 1650.510 2735.870 ;
        RECT 1647.730 2733.090 1648.910 2734.270 ;
        RECT 1649.330 2733.090 1650.510 2734.270 ;
        RECT 1647.730 2554.690 1648.910 2555.870 ;
        RECT 1649.330 2554.690 1650.510 2555.870 ;
        RECT 1647.730 2553.090 1648.910 2554.270 ;
        RECT 1649.330 2553.090 1650.510 2554.270 ;
        RECT 1647.730 2374.690 1648.910 2375.870 ;
        RECT 1649.330 2374.690 1650.510 2375.870 ;
        RECT 1647.730 2373.090 1648.910 2374.270 ;
        RECT 1649.330 2373.090 1650.510 2374.270 ;
        RECT 1647.730 2194.690 1648.910 2195.870 ;
        RECT 1649.330 2194.690 1650.510 2195.870 ;
        RECT 1647.730 2193.090 1648.910 2194.270 ;
        RECT 1649.330 2193.090 1650.510 2194.270 ;
        RECT 1647.730 2014.690 1648.910 2015.870 ;
        RECT 1649.330 2014.690 1650.510 2015.870 ;
        RECT 1647.730 2013.090 1648.910 2014.270 ;
        RECT 1649.330 2013.090 1650.510 2014.270 ;
        RECT 1647.730 1834.690 1648.910 1835.870 ;
        RECT 1649.330 1834.690 1650.510 1835.870 ;
        RECT 1647.730 1833.090 1648.910 1834.270 ;
        RECT 1649.330 1833.090 1650.510 1834.270 ;
        RECT 1647.730 1654.690 1648.910 1655.870 ;
        RECT 1649.330 1654.690 1650.510 1655.870 ;
        RECT 1647.730 1653.090 1648.910 1654.270 ;
        RECT 1649.330 1653.090 1650.510 1654.270 ;
        RECT 1647.730 1474.690 1648.910 1475.870 ;
        RECT 1649.330 1474.690 1650.510 1475.870 ;
        RECT 1647.730 1473.090 1648.910 1474.270 ;
        RECT 1649.330 1473.090 1650.510 1474.270 ;
        RECT 1647.730 1294.690 1648.910 1295.870 ;
        RECT 1649.330 1294.690 1650.510 1295.870 ;
        RECT 1647.730 1293.090 1648.910 1294.270 ;
        RECT 1649.330 1293.090 1650.510 1294.270 ;
        RECT 1647.730 1114.690 1648.910 1115.870 ;
        RECT 1649.330 1114.690 1650.510 1115.870 ;
        RECT 1647.730 1113.090 1648.910 1114.270 ;
        RECT 1649.330 1113.090 1650.510 1114.270 ;
        RECT 1647.730 934.690 1648.910 935.870 ;
        RECT 1649.330 934.690 1650.510 935.870 ;
        RECT 1647.730 933.090 1648.910 934.270 ;
        RECT 1649.330 933.090 1650.510 934.270 ;
        RECT 1647.730 754.690 1648.910 755.870 ;
        RECT 1649.330 754.690 1650.510 755.870 ;
        RECT 1647.730 753.090 1648.910 754.270 ;
        RECT 1649.330 753.090 1650.510 754.270 ;
        RECT 1647.730 574.690 1648.910 575.870 ;
        RECT 1649.330 574.690 1650.510 575.870 ;
        RECT 1647.730 573.090 1648.910 574.270 ;
        RECT 1649.330 573.090 1650.510 574.270 ;
        RECT 1647.730 394.690 1648.910 395.870 ;
        RECT 1649.330 394.690 1650.510 395.870 ;
        RECT 1647.730 393.090 1648.910 394.270 ;
        RECT 1649.330 393.090 1650.510 394.270 ;
        RECT 1647.730 214.690 1648.910 215.870 ;
        RECT 1649.330 214.690 1650.510 215.870 ;
        RECT 1647.730 213.090 1648.910 214.270 ;
        RECT 1649.330 213.090 1650.510 214.270 ;
        RECT 1647.730 34.690 1648.910 35.870 ;
        RECT 1649.330 34.690 1650.510 35.870 ;
        RECT 1647.730 33.090 1648.910 34.270 ;
        RECT 1649.330 33.090 1650.510 34.270 ;
        RECT 1647.730 -12.510 1648.910 -11.330 ;
        RECT 1649.330 -12.510 1650.510 -11.330 ;
        RECT 1647.730 -14.110 1648.910 -12.930 ;
        RECT 1649.330 -14.110 1650.510 -12.930 ;
        RECT 1827.730 3532.610 1828.910 3533.790 ;
        RECT 1829.330 3532.610 1830.510 3533.790 ;
        RECT 1827.730 3531.010 1828.910 3532.190 ;
        RECT 1829.330 3531.010 1830.510 3532.190 ;
        RECT 1827.730 3454.690 1828.910 3455.870 ;
        RECT 1829.330 3454.690 1830.510 3455.870 ;
        RECT 1827.730 3453.090 1828.910 3454.270 ;
        RECT 1829.330 3453.090 1830.510 3454.270 ;
        RECT 1827.730 3274.690 1828.910 3275.870 ;
        RECT 1829.330 3274.690 1830.510 3275.870 ;
        RECT 1827.730 3273.090 1828.910 3274.270 ;
        RECT 1829.330 3273.090 1830.510 3274.270 ;
        RECT 1827.730 3094.690 1828.910 3095.870 ;
        RECT 1829.330 3094.690 1830.510 3095.870 ;
        RECT 1827.730 3093.090 1828.910 3094.270 ;
        RECT 1829.330 3093.090 1830.510 3094.270 ;
        RECT 1827.730 2914.690 1828.910 2915.870 ;
        RECT 1829.330 2914.690 1830.510 2915.870 ;
        RECT 1827.730 2913.090 1828.910 2914.270 ;
        RECT 1829.330 2913.090 1830.510 2914.270 ;
        RECT 1827.730 2734.690 1828.910 2735.870 ;
        RECT 1829.330 2734.690 1830.510 2735.870 ;
        RECT 1827.730 2733.090 1828.910 2734.270 ;
        RECT 1829.330 2733.090 1830.510 2734.270 ;
        RECT 1827.730 2554.690 1828.910 2555.870 ;
        RECT 1829.330 2554.690 1830.510 2555.870 ;
        RECT 1827.730 2553.090 1828.910 2554.270 ;
        RECT 1829.330 2553.090 1830.510 2554.270 ;
        RECT 1827.730 2374.690 1828.910 2375.870 ;
        RECT 1829.330 2374.690 1830.510 2375.870 ;
        RECT 1827.730 2373.090 1828.910 2374.270 ;
        RECT 1829.330 2373.090 1830.510 2374.270 ;
        RECT 1827.730 2194.690 1828.910 2195.870 ;
        RECT 1829.330 2194.690 1830.510 2195.870 ;
        RECT 1827.730 2193.090 1828.910 2194.270 ;
        RECT 1829.330 2193.090 1830.510 2194.270 ;
        RECT 1827.730 2014.690 1828.910 2015.870 ;
        RECT 1829.330 2014.690 1830.510 2015.870 ;
        RECT 1827.730 2013.090 1828.910 2014.270 ;
        RECT 1829.330 2013.090 1830.510 2014.270 ;
        RECT 1827.730 1834.690 1828.910 1835.870 ;
        RECT 1829.330 1834.690 1830.510 1835.870 ;
        RECT 1827.730 1833.090 1828.910 1834.270 ;
        RECT 1829.330 1833.090 1830.510 1834.270 ;
        RECT 1827.730 1654.690 1828.910 1655.870 ;
        RECT 1829.330 1654.690 1830.510 1655.870 ;
        RECT 1827.730 1653.090 1828.910 1654.270 ;
        RECT 1829.330 1653.090 1830.510 1654.270 ;
        RECT 1827.730 1474.690 1828.910 1475.870 ;
        RECT 1829.330 1474.690 1830.510 1475.870 ;
        RECT 1827.730 1473.090 1828.910 1474.270 ;
        RECT 1829.330 1473.090 1830.510 1474.270 ;
        RECT 1827.730 1294.690 1828.910 1295.870 ;
        RECT 1829.330 1294.690 1830.510 1295.870 ;
        RECT 1827.730 1293.090 1828.910 1294.270 ;
        RECT 1829.330 1293.090 1830.510 1294.270 ;
        RECT 1827.730 1114.690 1828.910 1115.870 ;
        RECT 1829.330 1114.690 1830.510 1115.870 ;
        RECT 1827.730 1113.090 1828.910 1114.270 ;
        RECT 1829.330 1113.090 1830.510 1114.270 ;
        RECT 1827.730 934.690 1828.910 935.870 ;
        RECT 1829.330 934.690 1830.510 935.870 ;
        RECT 1827.730 933.090 1828.910 934.270 ;
        RECT 1829.330 933.090 1830.510 934.270 ;
        RECT 1827.730 754.690 1828.910 755.870 ;
        RECT 1829.330 754.690 1830.510 755.870 ;
        RECT 1827.730 753.090 1828.910 754.270 ;
        RECT 1829.330 753.090 1830.510 754.270 ;
        RECT 1827.730 574.690 1828.910 575.870 ;
        RECT 1829.330 574.690 1830.510 575.870 ;
        RECT 1827.730 573.090 1828.910 574.270 ;
        RECT 1829.330 573.090 1830.510 574.270 ;
        RECT 1827.730 394.690 1828.910 395.870 ;
        RECT 1829.330 394.690 1830.510 395.870 ;
        RECT 1827.730 393.090 1828.910 394.270 ;
        RECT 1829.330 393.090 1830.510 394.270 ;
        RECT 1827.730 214.690 1828.910 215.870 ;
        RECT 1829.330 214.690 1830.510 215.870 ;
        RECT 1827.730 213.090 1828.910 214.270 ;
        RECT 1829.330 213.090 1830.510 214.270 ;
        RECT 1827.730 34.690 1828.910 35.870 ;
        RECT 1829.330 34.690 1830.510 35.870 ;
        RECT 1827.730 33.090 1828.910 34.270 ;
        RECT 1829.330 33.090 1830.510 34.270 ;
        RECT 1827.730 -12.510 1828.910 -11.330 ;
        RECT 1829.330 -12.510 1830.510 -11.330 ;
        RECT 1827.730 -14.110 1828.910 -12.930 ;
        RECT 1829.330 -14.110 1830.510 -12.930 ;
        RECT 2007.730 3532.610 2008.910 3533.790 ;
        RECT 2009.330 3532.610 2010.510 3533.790 ;
        RECT 2007.730 3531.010 2008.910 3532.190 ;
        RECT 2009.330 3531.010 2010.510 3532.190 ;
        RECT 2007.730 3454.690 2008.910 3455.870 ;
        RECT 2009.330 3454.690 2010.510 3455.870 ;
        RECT 2007.730 3453.090 2008.910 3454.270 ;
        RECT 2009.330 3453.090 2010.510 3454.270 ;
        RECT 2007.730 3274.690 2008.910 3275.870 ;
        RECT 2009.330 3274.690 2010.510 3275.870 ;
        RECT 2007.730 3273.090 2008.910 3274.270 ;
        RECT 2009.330 3273.090 2010.510 3274.270 ;
        RECT 2007.730 3094.690 2008.910 3095.870 ;
        RECT 2009.330 3094.690 2010.510 3095.870 ;
        RECT 2007.730 3093.090 2008.910 3094.270 ;
        RECT 2009.330 3093.090 2010.510 3094.270 ;
        RECT 2007.730 2914.690 2008.910 2915.870 ;
        RECT 2009.330 2914.690 2010.510 2915.870 ;
        RECT 2007.730 2913.090 2008.910 2914.270 ;
        RECT 2009.330 2913.090 2010.510 2914.270 ;
        RECT 2007.730 2734.690 2008.910 2735.870 ;
        RECT 2009.330 2734.690 2010.510 2735.870 ;
        RECT 2007.730 2733.090 2008.910 2734.270 ;
        RECT 2009.330 2733.090 2010.510 2734.270 ;
        RECT 2007.730 2554.690 2008.910 2555.870 ;
        RECT 2009.330 2554.690 2010.510 2555.870 ;
        RECT 2007.730 2553.090 2008.910 2554.270 ;
        RECT 2009.330 2553.090 2010.510 2554.270 ;
        RECT 2007.730 2374.690 2008.910 2375.870 ;
        RECT 2009.330 2374.690 2010.510 2375.870 ;
        RECT 2007.730 2373.090 2008.910 2374.270 ;
        RECT 2009.330 2373.090 2010.510 2374.270 ;
        RECT 2007.730 2194.690 2008.910 2195.870 ;
        RECT 2009.330 2194.690 2010.510 2195.870 ;
        RECT 2007.730 2193.090 2008.910 2194.270 ;
        RECT 2009.330 2193.090 2010.510 2194.270 ;
        RECT 2007.730 2014.690 2008.910 2015.870 ;
        RECT 2009.330 2014.690 2010.510 2015.870 ;
        RECT 2007.730 2013.090 2008.910 2014.270 ;
        RECT 2009.330 2013.090 2010.510 2014.270 ;
        RECT 2007.730 1834.690 2008.910 1835.870 ;
        RECT 2009.330 1834.690 2010.510 1835.870 ;
        RECT 2007.730 1833.090 2008.910 1834.270 ;
        RECT 2009.330 1833.090 2010.510 1834.270 ;
        RECT 2007.730 1654.690 2008.910 1655.870 ;
        RECT 2009.330 1654.690 2010.510 1655.870 ;
        RECT 2007.730 1653.090 2008.910 1654.270 ;
        RECT 2009.330 1653.090 2010.510 1654.270 ;
        RECT 2007.730 1474.690 2008.910 1475.870 ;
        RECT 2009.330 1474.690 2010.510 1475.870 ;
        RECT 2007.730 1473.090 2008.910 1474.270 ;
        RECT 2009.330 1473.090 2010.510 1474.270 ;
        RECT 2007.730 1294.690 2008.910 1295.870 ;
        RECT 2009.330 1294.690 2010.510 1295.870 ;
        RECT 2007.730 1293.090 2008.910 1294.270 ;
        RECT 2009.330 1293.090 2010.510 1294.270 ;
        RECT 2007.730 1114.690 2008.910 1115.870 ;
        RECT 2009.330 1114.690 2010.510 1115.870 ;
        RECT 2007.730 1113.090 2008.910 1114.270 ;
        RECT 2009.330 1113.090 2010.510 1114.270 ;
        RECT 2007.730 934.690 2008.910 935.870 ;
        RECT 2009.330 934.690 2010.510 935.870 ;
        RECT 2007.730 933.090 2008.910 934.270 ;
        RECT 2009.330 933.090 2010.510 934.270 ;
        RECT 2007.730 754.690 2008.910 755.870 ;
        RECT 2009.330 754.690 2010.510 755.870 ;
        RECT 2007.730 753.090 2008.910 754.270 ;
        RECT 2009.330 753.090 2010.510 754.270 ;
        RECT 2007.730 574.690 2008.910 575.870 ;
        RECT 2009.330 574.690 2010.510 575.870 ;
        RECT 2007.730 573.090 2008.910 574.270 ;
        RECT 2009.330 573.090 2010.510 574.270 ;
        RECT 2007.730 394.690 2008.910 395.870 ;
        RECT 2009.330 394.690 2010.510 395.870 ;
        RECT 2007.730 393.090 2008.910 394.270 ;
        RECT 2009.330 393.090 2010.510 394.270 ;
        RECT 2007.730 214.690 2008.910 215.870 ;
        RECT 2009.330 214.690 2010.510 215.870 ;
        RECT 2007.730 213.090 2008.910 214.270 ;
        RECT 2009.330 213.090 2010.510 214.270 ;
        RECT 2007.730 34.690 2008.910 35.870 ;
        RECT 2009.330 34.690 2010.510 35.870 ;
        RECT 2007.730 33.090 2008.910 34.270 ;
        RECT 2009.330 33.090 2010.510 34.270 ;
        RECT 2007.730 -12.510 2008.910 -11.330 ;
        RECT 2009.330 -12.510 2010.510 -11.330 ;
        RECT 2007.730 -14.110 2008.910 -12.930 ;
        RECT 2009.330 -14.110 2010.510 -12.930 ;
        RECT 2187.730 3532.610 2188.910 3533.790 ;
        RECT 2189.330 3532.610 2190.510 3533.790 ;
        RECT 2187.730 3531.010 2188.910 3532.190 ;
        RECT 2189.330 3531.010 2190.510 3532.190 ;
        RECT 2187.730 3454.690 2188.910 3455.870 ;
        RECT 2189.330 3454.690 2190.510 3455.870 ;
        RECT 2187.730 3453.090 2188.910 3454.270 ;
        RECT 2189.330 3453.090 2190.510 3454.270 ;
        RECT 2187.730 3274.690 2188.910 3275.870 ;
        RECT 2189.330 3274.690 2190.510 3275.870 ;
        RECT 2187.730 3273.090 2188.910 3274.270 ;
        RECT 2189.330 3273.090 2190.510 3274.270 ;
        RECT 2187.730 3094.690 2188.910 3095.870 ;
        RECT 2189.330 3094.690 2190.510 3095.870 ;
        RECT 2187.730 3093.090 2188.910 3094.270 ;
        RECT 2189.330 3093.090 2190.510 3094.270 ;
        RECT 2187.730 2914.690 2188.910 2915.870 ;
        RECT 2189.330 2914.690 2190.510 2915.870 ;
        RECT 2187.730 2913.090 2188.910 2914.270 ;
        RECT 2189.330 2913.090 2190.510 2914.270 ;
        RECT 2187.730 2734.690 2188.910 2735.870 ;
        RECT 2189.330 2734.690 2190.510 2735.870 ;
        RECT 2187.730 2733.090 2188.910 2734.270 ;
        RECT 2189.330 2733.090 2190.510 2734.270 ;
        RECT 2187.730 2554.690 2188.910 2555.870 ;
        RECT 2189.330 2554.690 2190.510 2555.870 ;
        RECT 2187.730 2553.090 2188.910 2554.270 ;
        RECT 2189.330 2553.090 2190.510 2554.270 ;
        RECT 2187.730 2374.690 2188.910 2375.870 ;
        RECT 2189.330 2374.690 2190.510 2375.870 ;
        RECT 2187.730 2373.090 2188.910 2374.270 ;
        RECT 2189.330 2373.090 2190.510 2374.270 ;
        RECT 2187.730 2194.690 2188.910 2195.870 ;
        RECT 2189.330 2194.690 2190.510 2195.870 ;
        RECT 2187.730 2193.090 2188.910 2194.270 ;
        RECT 2189.330 2193.090 2190.510 2194.270 ;
        RECT 2187.730 2014.690 2188.910 2015.870 ;
        RECT 2189.330 2014.690 2190.510 2015.870 ;
        RECT 2187.730 2013.090 2188.910 2014.270 ;
        RECT 2189.330 2013.090 2190.510 2014.270 ;
        RECT 2187.730 1834.690 2188.910 1835.870 ;
        RECT 2189.330 1834.690 2190.510 1835.870 ;
        RECT 2187.730 1833.090 2188.910 1834.270 ;
        RECT 2189.330 1833.090 2190.510 1834.270 ;
        RECT 2187.730 1654.690 2188.910 1655.870 ;
        RECT 2189.330 1654.690 2190.510 1655.870 ;
        RECT 2187.730 1653.090 2188.910 1654.270 ;
        RECT 2189.330 1653.090 2190.510 1654.270 ;
        RECT 2187.730 1474.690 2188.910 1475.870 ;
        RECT 2189.330 1474.690 2190.510 1475.870 ;
        RECT 2187.730 1473.090 2188.910 1474.270 ;
        RECT 2189.330 1473.090 2190.510 1474.270 ;
        RECT 2187.730 1294.690 2188.910 1295.870 ;
        RECT 2189.330 1294.690 2190.510 1295.870 ;
        RECT 2187.730 1293.090 2188.910 1294.270 ;
        RECT 2189.330 1293.090 2190.510 1294.270 ;
        RECT 2187.730 1114.690 2188.910 1115.870 ;
        RECT 2189.330 1114.690 2190.510 1115.870 ;
        RECT 2187.730 1113.090 2188.910 1114.270 ;
        RECT 2189.330 1113.090 2190.510 1114.270 ;
        RECT 2187.730 934.690 2188.910 935.870 ;
        RECT 2189.330 934.690 2190.510 935.870 ;
        RECT 2187.730 933.090 2188.910 934.270 ;
        RECT 2189.330 933.090 2190.510 934.270 ;
        RECT 2187.730 754.690 2188.910 755.870 ;
        RECT 2189.330 754.690 2190.510 755.870 ;
        RECT 2187.730 753.090 2188.910 754.270 ;
        RECT 2189.330 753.090 2190.510 754.270 ;
        RECT 2187.730 574.690 2188.910 575.870 ;
        RECT 2189.330 574.690 2190.510 575.870 ;
        RECT 2187.730 573.090 2188.910 574.270 ;
        RECT 2189.330 573.090 2190.510 574.270 ;
        RECT 2187.730 394.690 2188.910 395.870 ;
        RECT 2189.330 394.690 2190.510 395.870 ;
        RECT 2187.730 393.090 2188.910 394.270 ;
        RECT 2189.330 393.090 2190.510 394.270 ;
        RECT 2187.730 214.690 2188.910 215.870 ;
        RECT 2189.330 214.690 2190.510 215.870 ;
        RECT 2187.730 213.090 2188.910 214.270 ;
        RECT 2189.330 213.090 2190.510 214.270 ;
        RECT 2187.730 34.690 2188.910 35.870 ;
        RECT 2189.330 34.690 2190.510 35.870 ;
        RECT 2187.730 33.090 2188.910 34.270 ;
        RECT 2189.330 33.090 2190.510 34.270 ;
        RECT 2187.730 -12.510 2188.910 -11.330 ;
        RECT 2189.330 -12.510 2190.510 -11.330 ;
        RECT 2187.730 -14.110 2188.910 -12.930 ;
        RECT 2189.330 -14.110 2190.510 -12.930 ;
        RECT 2367.730 3532.610 2368.910 3533.790 ;
        RECT 2369.330 3532.610 2370.510 3533.790 ;
        RECT 2367.730 3531.010 2368.910 3532.190 ;
        RECT 2369.330 3531.010 2370.510 3532.190 ;
        RECT 2367.730 3454.690 2368.910 3455.870 ;
        RECT 2369.330 3454.690 2370.510 3455.870 ;
        RECT 2367.730 3453.090 2368.910 3454.270 ;
        RECT 2369.330 3453.090 2370.510 3454.270 ;
        RECT 2367.730 3274.690 2368.910 3275.870 ;
        RECT 2369.330 3274.690 2370.510 3275.870 ;
        RECT 2367.730 3273.090 2368.910 3274.270 ;
        RECT 2369.330 3273.090 2370.510 3274.270 ;
        RECT 2367.730 3094.690 2368.910 3095.870 ;
        RECT 2369.330 3094.690 2370.510 3095.870 ;
        RECT 2367.730 3093.090 2368.910 3094.270 ;
        RECT 2369.330 3093.090 2370.510 3094.270 ;
        RECT 2367.730 2914.690 2368.910 2915.870 ;
        RECT 2369.330 2914.690 2370.510 2915.870 ;
        RECT 2367.730 2913.090 2368.910 2914.270 ;
        RECT 2369.330 2913.090 2370.510 2914.270 ;
        RECT 2367.730 2734.690 2368.910 2735.870 ;
        RECT 2369.330 2734.690 2370.510 2735.870 ;
        RECT 2367.730 2733.090 2368.910 2734.270 ;
        RECT 2369.330 2733.090 2370.510 2734.270 ;
        RECT 2367.730 2554.690 2368.910 2555.870 ;
        RECT 2369.330 2554.690 2370.510 2555.870 ;
        RECT 2367.730 2553.090 2368.910 2554.270 ;
        RECT 2369.330 2553.090 2370.510 2554.270 ;
        RECT 2367.730 2374.690 2368.910 2375.870 ;
        RECT 2369.330 2374.690 2370.510 2375.870 ;
        RECT 2367.730 2373.090 2368.910 2374.270 ;
        RECT 2369.330 2373.090 2370.510 2374.270 ;
        RECT 2367.730 2194.690 2368.910 2195.870 ;
        RECT 2369.330 2194.690 2370.510 2195.870 ;
        RECT 2367.730 2193.090 2368.910 2194.270 ;
        RECT 2369.330 2193.090 2370.510 2194.270 ;
        RECT 2367.730 2014.690 2368.910 2015.870 ;
        RECT 2369.330 2014.690 2370.510 2015.870 ;
        RECT 2367.730 2013.090 2368.910 2014.270 ;
        RECT 2369.330 2013.090 2370.510 2014.270 ;
        RECT 2367.730 1834.690 2368.910 1835.870 ;
        RECT 2369.330 1834.690 2370.510 1835.870 ;
        RECT 2367.730 1833.090 2368.910 1834.270 ;
        RECT 2369.330 1833.090 2370.510 1834.270 ;
        RECT 2367.730 1654.690 2368.910 1655.870 ;
        RECT 2369.330 1654.690 2370.510 1655.870 ;
        RECT 2367.730 1653.090 2368.910 1654.270 ;
        RECT 2369.330 1653.090 2370.510 1654.270 ;
        RECT 2367.730 1474.690 2368.910 1475.870 ;
        RECT 2369.330 1474.690 2370.510 1475.870 ;
        RECT 2367.730 1473.090 2368.910 1474.270 ;
        RECT 2369.330 1473.090 2370.510 1474.270 ;
        RECT 2367.730 1294.690 2368.910 1295.870 ;
        RECT 2369.330 1294.690 2370.510 1295.870 ;
        RECT 2367.730 1293.090 2368.910 1294.270 ;
        RECT 2369.330 1293.090 2370.510 1294.270 ;
        RECT 2367.730 1114.690 2368.910 1115.870 ;
        RECT 2369.330 1114.690 2370.510 1115.870 ;
        RECT 2367.730 1113.090 2368.910 1114.270 ;
        RECT 2369.330 1113.090 2370.510 1114.270 ;
        RECT 2367.730 934.690 2368.910 935.870 ;
        RECT 2369.330 934.690 2370.510 935.870 ;
        RECT 2367.730 933.090 2368.910 934.270 ;
        RECT 2369.330 933.090 2370.510 934.270 ;
        RECT 2367.730 754.690 2368.910 755.870 ;
        RECT 2369.330 754.690 2370.510 755.870 ;
        RECT 2367.730 753.090 2368.910 754.270 ;
        RECT 2369.330 753.090 2370.510 754.270 ;
        RECT 2367.730 574.690 2368.910 575.870 ;
        RECT 2369.330 574.690 2370.510 575.870 ;
        RECT 2367.730 573.090 2368.910 574.270 ;
        RECT 2369.330 573.090 2370.510 574.270 ;
        RECT 2367.730 394.690 2368.910 395.870 ;
        RECT 2369.330 394.690 2370.510 395.870 ;
        RECT 2367.730 393.090 2368.910 394.270 ;
        RECT 2369.330 393.090 2370.510 394.270 ;
        RECT 2367.730 214.690 2368.910 215.870 ;
        RECT 2369.330 214.690 2370.510 215.870 ;
        RECT 2367.730 213.090 2368.910 214.270 ;
        RECT 2369.330 213.090 2370.510 214.270 ;
        RECT 2367.730 34.690 2368.910 35.870 ;
        RECT 2369.330 34.690 2370.510 35.870 ;
        RECT 2367.730 33.090 2368.910 34.270 ;
        RECT 2369.330 33.090 2370.510 34.270 ;
        RECT 2367.730 -12.510 2368.910 -11.330 ;
        RECT 2369.330 -12.510 2370.510 -11.330 ;
        RECT 2367.730 -14.110 2368.910 -12.930 ;
        RECT 2369.330 -14.110 2370.510 -12.930 ;
        RECT 2547.730 3532.610 2548.910 3533.790 ;
        RECT 2549.330 3532.610 2550.510 3533.790 ;
        RECT 2547.730 3531.010 2548.910 3532.190 ;
        RECT 2549.330 3531.010 2550.510 3532.190 ;
        RECT 2547.730 3454.690 2548.910 3455.870 ;
        RECT 2549.330 3454.690 2550.510 3455.870 ;
        RECT 2547.730 3453.090 2548.910 3454.270 ;
        RECT 2549.330 3453.090 2550.510 3454.270 ;
        RECT 2547.730 3274.690 2548.910 3275.870 ;
        RECT 2549.330 3274.690 2550.510 3275.870 ;
        RECT 2547.730 3273.090 2548.910 3274.270 ;
        RECT 2549.330 3273.090 2550.510 3274.270 ;
        RECT 2547.730 3094.690 2548.910 3095.870 ;
        RECT 2549.330 3094.690 2550.510 3095.870 ;
        RECT 2547.730 3093.090 2548.910 3094.270 ;
        RECT 2549.330 3093.090 2550.510 3094.270 ;
        RECT 2547.730 2914.690 2548.910 2915.870 ;
        RECT 2549.330 2914.690 2550.510 2915.870 ;
        RECT 2547.730 2913.090 2548.910 2914.270 ;
        RECT 2549.330 2913.090 2550.510 2914.270 ;
        RECT 2547.730 2734.690 2548.910 2735.870 ;
        RECT 2549.330 2734.690 2550.510 2735.870 ;
        RECT 2547.730 2733.090 2548.910 2734.270 ;
        RECT 2549.330 2733.090 2550.510 2734.270 ;
        RECT 2547.730 2554.690 2548.910 2555.870 ;
        RECT 2549.330 2554.690 2550.510 2555.870 ;
        RECT 2547.730 2553.090 2548.910 2554.270 ;
        RECT 2549.330 2553.090 2550.510 2554.270 ;
        RECT 2547.730 2374.690 2548.910 2375.870 ;
        RECT 2549.330 2374.690 2550.510 2375.870 ;
        RECT 2547.730 2373.090 2548.910 2374.270 ;
        RECT 2549.330 2373.090 2550.510 2374.270 ;
        RECT 2547.730 2194.690 2548.910 2195.870 ;
        RECT 2549.330 2194.690 2550.510 2195.870 ;
        RECT 2547.730 2193.090 2548.910 2194.270 ;
        RECT 2549.330 2193.090 2550.510 2194.270 ;
        RECT 2547.730 2014.690 2548.910 2015.870 ;
        RECT 2549.330 2014.690 2550.510 2015.870 ;
        RECT 2547.730 2013.090 2548.910 2014.270 ;
        RECT 2549.330 2013.090 2550.510 2014.270 ;
        RECT 2547.730 1834.690 2548.910 1835.870 ;
        RECT 2549.330 1834.690 2550.510 1835.870 ;
        RECT 2547.730 1833.090 2548.910 1834.270 ;
        RECT 2549.330 1833.090 2550.510 1834.270 ;
        RECT 2547.730 1654.690 2548.910 1655.870 ;
        RECT 2549.330 1654.690 2550.510 1655.870 ;
        RECT 2547.730 1653.090 2548.910 1654.270 ;
        RECT 2549.330 1653.090 2550.510 1654.270 ;
        RECT 2547.730 1474.690 2548.910 1475.870 ;
        RECT 2549.330 1474.690 2550.510 1475.870 ;
        RECT 2547.730 1473.090 2548.910 1474.270 ;
        RECT 2549.330 1473.090 2550.510 1474.270 ;
        RECT 2547.730 1294.690 2548.910 1295.870 ;
        RECT 2549.330 1294.690 2550.510 1295.870 ;
        RECT 2547.730 1293.090 2548.910 1294.270 ;
        RECT 2549.330 1293.090 2550.510 1294.270 ;
        RECT 2547.730 1114.690 2548.910 1115.870 ;
        RECT 2549.330 1114.690 2550.510 1115.870 ;
        RECT 2547.730 1113.090 2548.910 1114.270 ;
        RECT 2549.330 1113.090 2550.510 1114.270 ;
        RECT 2547.730 934.690 2548.910 935.870 ;
        RECT 2549.330 934.690 2550.510 935.870 ;
        RECT 2547.730 933.090 2548.910 934.270 ;
        RECT 2549.330 933.090 2550.510 934.270 ;
        RECT 2547.730 754.690 2548.910 755.870 ;
        RECT 2549.330 754.690 2550.510 755.870 ;
        RECT 2547.730 753.090 2548.910 754.270 ;
        RECT 2549.330 753.090 2550.510 754.270 ;
        RECT 2547.730 574.690 2548.910 575.870 ;
        RECT 2549.330 574.690 2550.510 575.870 ;
        RECT 2547.730 573.090 2548.910 574.270 ;
        RECT 2549.330 573.090 2550.510 574.270 ;
        RECT 2547.730 394.690 2548.910 395.870 ;
        RECT 2549.330 394.690 2550.510 395.870 ;
        RECT 2547.730 393.090 2548.910 394.270 ;
        RECT 2549.330 393.090 2550.510 394.270 ;
        RECT 2547.730 214.690 2548.910 215.870 ;
        RECT 2549.330 214.690 2550.510 215.870 ;
        RECT 2547.730 213.090 2548.910 214.270 ;
        RECT 2549.330 213.090 2550.510 214.270 ;
        RECT 2547.730 34.690 2548.910 35.870 ;
        RECT 2549.330 34.690 2550.510 35.870 ;
        RECT 2547.730 33.090 2548.910 34.270 ;
        RECT 2549.330 33.090 2550.510 34.270 ;
        RECT 2547.730 -12.510 2548.910 -11.330 ;
        RECT 2549.330 -12.510 2550.510 -11.330 ;
        RECT 2547.730 -14.110 2548.910 -12.930 ;
        RECT 2549.330 -14.110 2550.510 -12.930 ;
        RECT 2727.730 3532.610 2728.910 3533.790 ;
        RECT 2729.330 3532.610 2730.510 3533.790 ;
        RECT 2727.730 3531.010 2728.910 3532.190 ;
        RECT 2729.330 3531.010 2730.510 3532.190 ;
        RECT 2727.730 3454.690 2728.910 3455.870 ;
        RECT 2729.330 3454.690 2730.510 3455.870 ;
        RECT 2727.730 3453.090 2728.910 3454.270 ;
        RECT 2729.330 3453.090 2730.510 3454.270 ;
        RECT 2727.730 3274.690 2728.910 3275.870 ;
        RECT 2729.330 3274.690 2730.510 3275.870 ;
        RECT 2727.730 3273.090 2728.910 3274.270 ;
        RECT 2729.330 3273.090 2730.510 3274.270 ;
        RECT 2727.730 3094.690 2728.910 3095.870 ;
        RECT 2729.330 3094.690 2730.510 3095.870 ;
        RECT 2727.730 3093.090 2728.910 3094.270 ;
        RECT 2729.330 3093.090 2730.510 3094.270 ;
        RECT 2727.730 2914.690 2728.910 2915.870 ;
        RECT 2729.330 2914.690 2730.510 2915.870 ;
        RECT 2727.730 2913.090 2728.910 2914.270 ;
        RECT 2729.330 2913.090 2730.510 2914.270 ;
        RECT 2727.730 2734.690 2728.910 2735.870 ;
        RECT 2729.330 2734.690 2730.510 2735.870 ;
        RECT 2727.730 2733.090 2728.910 2734.270 ;
        RECT 2729.330 2733.090 2730.510 2734.270 ;
        RECT 2727.730 2554.690 2728.910 2555.870 ;
        RECT 2729.330 2554.690 2730.510 2555.870 ;
        RECT 2727.730 2553.090 2728.910 2554.270 ;
        RECT 2729.330 2553.090 2730.510 2554.270 ;
        RECT 2727.730 2374.690 2728.910 2375.870 ;
        RECT 2729.330 2374.690 2730.510 2375.870 ;
        RECT 2727.730 2373.090 2728.910 2374.270 ;
        RECT 2729.330 2373.090 2730.510 2374.270 ;
        RECT 2727.730 2194.690 2728.910 2195.870 ;
        RECT 2729.330 2194.690 2730.510 2195.870 ;
        RECT 2727.730 2193.090 2728.910 2194.270 ;
        RECT 2729.330 2193.090 2730.510 2194.270 ;
        RECT 2727.730 2014.690 2728.910 2015.870 ;
        RECT 2729.330 2014.690 2730.510 2015.870 ;
        RECT 2727.730 2013.090 2728.910 2014.270 ;
        RECT 2729.330 2013.090 2730.510 2014.270 ;
        RECT 2727.730 1834.690 2728.910 1835.870 ;
        RECT 2729.330 1834.690 2730.510 1835.870 ;
        RECT 2727.730 1833.090 2728.910 1834.270 ;
        RECT 2729.330 1833.090 2730.510 1834.270 ;
        RECT 2727.730 1654.690 2728.910 1655.870 ;
        RECT 2729.330 1654.690 2730.510 1655.870 ;
        RECT 2727.730 1653.090 2728.910 1654.270 ;
        RECT 2729.330 1653.090 2730.510 1654.270 ;
        RECT 2727.730 1474.690 2728.910 1475.870 ;
        RECT 2729.330 1474.690 2730.510 1475.870 ;
        RECT 2727.730 1473.090 2728.910 1474.270 ;
        RECT 2729.330 1473.090 2730.510 1474.270 ;
        RECT 2727.730 1294.690 2728.910 1295.870 ;
        RECT 2729.330 1294.690 2730.510 1295.870 ;
        RECT 2727.730 1293.090 2728.910 1294.270 ;
        RECT 2729.330 1293.090 2730.510 1294.270 ;
        RECT 2727.730 1114.690 2728.910 1115.870 ;
        RECT 2729.330 1114.690 2730.510 1115.870 ;
        RECT 2727.730 1113.090 2728.910 1114.270 ;
        RECT 2729.330 1113.090 2730.510 1114.270 ;
        RECT 2727.730 934.690 2728.910 935.870 ;
        RECT 2729.330 934.690 2730.510 935.870 ;
        RECT 2727.730 933.090 2728.910 934.270 ;
        RECT 2729.330 933.090 2730.510 934.270 ;
        RECT 2727.730 754.690 2728.910 755.870 ;
        RECT 2729.330 754.690 2730.510 755.870 ;
        RECT 2727.730 753.090 2728.910 754.270 ;
        RECT 2729.330 753.090 2730.510 754.270 ;
        RECT 2727.730 574.690 2728.910 575.870 ;
        RECT 2729.330 574.690 2730.510 575.870 ;
        RECT 2727.730 573.090 2728.910 574.270 ;
        RECT 2729.330 573.090 2730.510 574.270 ;
        RECT 2727.730 394.690 2728.910 395.870 ;
        RECT 2729.330 394.690 2730.510 395.870 ;
        RECT 2727.730 393.090 2728.910 394.270 ;
        RECT 2729.330 393.090 2730.510 394.270 ;
        RECT 2727.730 214.690 2728.910 215.870 ;
        RECT 2729.330 214.690 2730.510 215.870 ;
        RECT 2727.730 213.090 2728.910 214.270 ;
        RECT 2729.330 213.090 2730.510 214.270 ;
        RECT 2727.730 34.690 2728.910 35.870 ;
        RECT 2729.330 34.690 2730.510 35.870 ;
        RECT 2727.730 33.090 2728.910 34.270 ;
        RECT 2729.330 33.090 2730.510 34.270 ;
        RECT 2727.730 -12.510 2728.910 -11.330 ;
        RECT 2729.330 -12.510 2730.510 -11.330 ;
        RECT 2727.730 -14.110 2728.910 -12.930 ;
        RECT 2729.330 -14.110 2730.510 -12.930 ;
        RECT 2907.730 3532.610 2908.910 3533.790 ;
        RECT 2909.330 3532.610 2910.510 3533.790 ;
        RECT 2907.730 3531.010 2908.910 3532.190 ;
        RECT 2909.330 3531.010 2910.510 3532.190 ;
        RECT 2907.730 3454.690 2908.910 3455.870 ;
        RECT 2909.330 3454.690 2910.510 3455.870 ;
        RECT 2907.730 3453.090 2908.910 3454.270 ;
        RECT 2909.330 3453.090 2910.510 3454.270 ;
        RECT 2907.730 3274.690 2908.910 3275.870 ;
        RECT 2909.330 3274.690 2910.510 3275.870 ;
        RECT 2907.730 3273.090 2908.910 3274.270 ;
        RECT 2909.330 3273.090 2910.510 3274.270 ;
        RECT 2907.730 3094.690 2908.910 3095.870 ;
        RECT 2909.330 3094.690 2910.510 3095.870 ;
        RECT 2907.730 3093.090 2908.910 3094.270 ;
        RECT 2909.330 3093.090 2910.510 3094.270 ;
        RECT 2907.730 2914.690 2908.910 2915.870 ;
        RECT 2909.330 2914.690 2910.510 2915.870 ;
        RECT 2907.730 2913.090 2908.910 2914.270 ;
        RECT 2909.330 2913.090 2910.510 2914.270 ;
        RECT 2907.730 2734.690 2908.910 2735.870 ;
        RECT 2909.330 2734.690 2910.510 2735.870 ;
        RECT 2907.730 2733.090 2908.910 2734.270 ;
        RECT 2909.330 2733.090 2910.510 2734.270 ;
        RECT 2907.730 2554.690 2908.910 2555.870 ;
        RECT 2909.330 2554.690 2910.510 2555.870 ;
        RECT 2907.730 2553.090 2908.910 2554.270 ;
        RECT 2909.330 2553.090 2910.510 2554.270 ;
        RECT 2907.730 2374.690 2908.910 2375.870 ;
        RECT 2909.330 2374.690 2910.510 2375.870 ;
        RECT 2907.730 2373.090 2908.910 2374.270 ;
        RECT 2909.330 2373.090 2910.510 2374.270 ;
        RECT 2907.730 2194.690 2908.910 2195.870 ;
        RECT 2909.330 2194.690 2910.510 2195.870 ;
        RECT 2907.730 2193.090 2908.910 2194.270 ;
        RECT 2909.330 2193.090 2910.510 2194.270 ;
        RECT 2907.730 2014.690 2908.910 2015.870 ;
        RECT 2909.330 2014.690 2910.510 2015.870 ;
        RECT 2907.730 2013.090 2908.910 2014.270 ;
        RECT 2909.330 2013.090 2910.510 2014.270 ;
        RECT 2907.730 1834.690 2908.910 1835.870 ;
        RECT 2909.330 1834.690 2910.510 1835.870 ;
        RECT 2907.730 1833.090 2908.910 1834.270 ;
        RECT 2909.330 1833.090 2910.510 1834.270 ;
        RECT 2907.730 1654.690 2908.910 1655.870 ;
        RECT 2909.330 1654.690 2910.510 1655.870 ;
        RECT 2907.730 1653.090 2908.910 1654.270 ;
        RECT 2909.330 1653.090 2910.510 1654.270 ;
        RECT 2907.730 1474.690 2908.910 1475.870 ;
        RECT 2909.330 1474.690 2910.510 1475.870 ;
        RECT 2907.730 1473.090 2908.910 1474.270 ;
        RECT 2909.330 1473.090 2910.510 1474.270 ;
        RECT 2907.730 1294.690 2908.910 1295.870 ;
        RECT 2909.330 1294.690 2910.510 1295.870 ;
        RECT 2907.730 1293.090 2908.910 1294.270 ;
        RECT 2909.330 1293.090 2910.510 1294.270 ;
        RECT 2907.730 1114.690 2908.910 1115.870 ;
        RECT 2909.330 1114.690 2910.510 1115.870 ;
        RECT 2907.730 1113.090 2908.910 1114.270 ;
        RECT 2909.330 1113.090 2910.510 1114.270 ;
        RECT 2907.730 934.690 2908.910 935.870 ;
        RECT 2909.330 934.690 2910.510 935.870 ;
        RECT 2907.730 933.090 2908.910 934.270 ;
        RECT 2909.330 933.090 2910.510 934.270 ;
        RECT 2907.730 754.690 2908.910 755.870 ;
        RECT 2909.330 754.690 2910.510 755.870 ;
        RECT 2907.730 753.090 2908.910 754.270 ;
        RECT 2909.330 753.090 2910.510 754.270 ;
        RECT 2907.730 574.690 2908.910 575.870 ;
        RECT 2909.330 574.690 2910.510 575.870 ;
        RECT 2907.730 573.090 2908.910 574.270 ;
        RECT 2909.330 573.090 2910.510 574.270 ;
        RECT 2907.730 394.690 2908.910 395.870 ;
        RECT 2909.330 394.690 2910.510 395.870 ;
        RECT 2907.730 393.090 2908.910 394.270 ;
        RECT 2909.330 393.090 2910.510 394.270 ;
        RECT 2907.730 214.690 2908.910 215.870 ;
        RECT 2909.330 214.690 2910.510 215.870 ;
        RECT 2907.730 213.090 2908.910 214.270 ;
        RECT 2909.330 213.090 2910.510 214.270 ;
        RECT 2907.730 34.690 2908.910 35.870 ;
        RECT 2909.330 34.690 2910.510 35.870 ;
        RECT 2907.730 33.090 2908.910 34.270 ;
        RECT 2909.330 33.090 2910.510 34.270 ;
        RECT 2907.730 -12.510 2908.910 -11.330 ;
        RECT 2909.330 -12.510 2910.510 -11.330 ;
        RECT 2907.730 -14.110 2908.910 -12.930 ;
        RECT 2909.330 -14.110 2910.510 -12.930 ;
        RECT 2936.310 3532.610 2937.490 3533.790 ;
        RECT 2937.910 3532.610 2939.090 3533.790 ;
        RECT 2936.310 3531.010 2937.490 3532.190 ;
        RECT 2937.910 3531.010 2939.090 3532.190 ;
        RECT 2936.310 3454.690 2937.490 3455.870 ;
        RECT 2937.910 3454.690 2939.090 3455.870 ;
        RECT 2936.310 3453.090 2937.490 3454.270 ;
        RECT 2937.910 3453.090 2939.090 3454.270 ;
        RECT 2936.310 3274.690 2937.490 3275.870 ;
        RECT 2937.910 3274.690 2939.090 3275.870 ;
        RECT 2936.310 3273.090 2937.490 3274.270 ;
        RECT 2937.910 3273.090 2939.090 3274.270 ;
        RECT 2936.310 3094.690 2937.490 3095.870 ;
        RECT 2937.910 3094.690 2939.090 3095.870 ;
        RECT 2936.310 3093.090 2937.490 3094.270 ;
        RECT 2937.910 3093.090 2939.090 3094.270 ;
        RECT 2936.310 2914.690 2937.490 2915.870 ;
        RECT 2937.910 2914.690 2939.090 2915.870 ;
        RECT 2936.310 2913.090 2937.490 2914.270 ;
        RECT 2937.910 2913.090 2939.090 2914.270 ;
        RECT 2936.310 2734.690 2937.490 2735.870 ;
        RECT 2937.910 2734.690 2939.090 2735.870 ;
        RECT 2936.310 2733.090 2937.490 2734.270 ;
        RECT 2937.910 2733.090 2939.090 2734.270 ;
        RECT 2936.310 2554.690 2937.490 2555.870 ;
        RECT 2937.910 2554.690 2939.090 2555.870 ;
        RECT 2936.310 2553.090 2937.490 2554.270 ;
        RECT 2937.910 2553.090 2939.090 2554.270 ;
        RECT 2936.310 2374.690 2937.490 2375.870 ;
        RECT 2937.910 2374.690 2939.090 2375.870 ;
        RECT 2936.310 2373.090 2937.490 2374.270 ;
        RECT 2937.910 2373.090 2939.090 2374.270 ;
        RECT 2936.310 2194.690 2937.490 2195.870 ;
        RECT 2937.910 2194.690 2939.090 2195.870 ;
        RECT 2936.310 2193.090 2937.490 2194.270 ;
        RECT 2937.910 2193.090 2939.090 2194.270 ;
        RECT 2936.310 2014.690 2937.490 2015.870 ;
        RECT 2937.910 2014.690 2939.090 2015.870 ;
        RECT 2936.310 2013.090 2937.490 2014.270 ;
        RECT 2937.910 2013.090 2939.090 2014.270 ;
        RECT 2936.310 1834.690 2937.490 1835.870 ;
        RECT 2937.910 1834.690 2939.090 1835.870 ;
        RECT 2936.310 1833.090 2937.490 1834.270 ;
        RECT 2937.910 1833.090 2939.090 1834.270 ;
        RECT 2936.310 1654.690 2937.490 1655.870 ;
        RECT 2937.910 1654.690 2939.090 1655.870 ;
        RECT 2936.310 1653.090 2937.490 1654.270 ;
        RECT 2937.910 1653.090 2939.090 1654.270 ;
        RECT 2936.310 1474.690 2937.490 1475.870 ;
        RECT 2937.910 1474.690 2939.090 1475.870 ;
        RECT 2936.310 1473.090 2937.490 1474.270 ;
        RECT 2937.910 1473.090 2939.090 1474.270 ;
        RECT 2936.310 1294.690 2937.490 1295.870 ;
        RECT 2937.910 1294.690 2939.090 1295.870 ;
        RECT 2936.310 1293.090 2937.490 1294.270 ;
        RECT 2937.910 1293.090 2939.090 1294.270 ;
        RECT 2936.310 1114.690 2937.490 1115.870 ;
        RECT 2937.910 1114.690 2939.090 1115.870 ;
        RECT 2936.310 1113.090 2937.490 1114.270 ;
        RECT 2937.910 1113.090 2939.090 1114.270 ;
        RECT 2936.310 934.690 2937.490 935.870 ;
        RECT 2937.910 934.690 2939.090 935.870 ;
        RECT 2936.310 933.090 2937.490 934.270 ;
        RECT 2937.910 933.090 2939.090 934.270 ;
        RECT 2936.310 754.690 2937.490 755.870 ;
        RECT 2937.910 754.690 2939.090 755.870 ;
        RECT 2936.310 753.090 2937.490 754.270 ;
        RECT 2937.910 753.090 2939.090 754.270 ;
        RECT 2936.310 574.690 2937.490 575.870 ;
        RECT 2937.910 574.690 2939.090 575.870 ;
        RECT 2936.310 573.090 2937.490 574.270 ;
        RECT 2937.910 573.090 2939.090 574.270 ;
        RECT 2936.310 394.690 2937.490 395.870 ;
        RECT 2937.910 394.690 2939.090 395.870 ;
        RECT 2936.310 393.090 2937.490 394.270 ;
        RECT 2937.910 393.090 2939.090 394.270 ;
        RECT 2936.310 214.690 2937.490 215.870 ;
        RECT 2937.910 214.690 2939.090 215.870 ;
        RECT 2936.310 213.090 2937.490 214.270 ;
        RECT 2937.910 213.090 2939.090 214.270 ;
        RECT 2936.310 34.690 2937.490 35.870 ;
        RECT 2937.910 34.690 2939.090 35.870 ;
        RECT 2936.310 33.090 2937.490 34.270 ;
        RECT 2937.910 33.090 2939.090 34.270 ;
        RECT 2936.310 -12.510 2937.490 -11.330 ;
        RECT 2937.910 -12.510 2939.090 -11.330 ;
        RECT 2936.310 -14.110 2937.490 -12.930 ;
        RECT 2937.910 -14.110 2939.090 -12.930 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
        RECT -24.430 932.930 2944.050 936.030 ;
        RECT -24.430 752.930 2944.050 756.030 ;
        RECT -24.430 572.930 2944.050 576.030 ;
        RECT -24.430 392.930 2944.050 396.030 ;
        RECT -24.430 212.930 2944.050 216.030 ;
        RECT -24.430 32.930 2944.050 36.030 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
        RECT 226.170 1010.000 229.270 3548.350 ;
        RECT 406.170 1010.000 409.270 3548.350 ;
        RECT 586.170 1010.000 589.270 3548.350 ;
        RECT 766.170 1010.000 769.270 3548.350 ;
        RECT 946.170 1010.000 949.270 3548.350 ;
        RECT 226.170 -28.670 229.270 390.000 ;
        RECT 406.170 -28.670 409.270 390.000 ;
        RECT 586.170 -28.670 589.270 390.000 ;
        RECT 766.170 -28.670 769.270 390.000 ;
        RECT 946.170 -28.670 949.270 390.000 ;
        RECT 1126.170 -28.670 1129.270 3548.350 ;
        RECT 1306.170 -28.670 1309.270 3548.350 ;
        RECT 1486.170 -28.670 1489.270 3548.350 ;
        RECT 1666.170 -28.670 1669.270 3548.350 ;
        RECT 1846.170 -28.670 1849.270 3548.350 ;
        RECT 2026.170 -28.670 2029.270 3548.350 ;
        RECT 2206.170 -28.670 2209.270 3548.350 ;
        RECT 2386.170 -28.670 2389.270 3548.350 ;
        RECT 2566.170 -28.670 2569.270 3548.350 ;
        RECT 2746.170 -28.670 2749.270 3548.350 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER via4 ;
        RECT -29.070 3542.210 -27.890 3543.390 ;
        RECT -27.470 3542.210 -26.290 3543.390 ;
        RECT -29.070 3540.610 -27.890 3541.790 ;
        RECT -27.470 3540.610 -26.290 3541.790 ;
        RECT -29.070 3473.290 -27.890 3474.470 ;
        RECT -27.470 3473.290 -26.290 3474.470 ;
        RECT -29.070 3471.690 -27.890 3472.870 ;
        RECT -27.470 3471.690 -26.290 3472.870 ;
        RECT -29.070 3293.290 -27.890 3294.470 ;
        RECT -27.470 3293.290 -26.290 3294.470 ;
        RECT -29.070 3291.690 -27.890 3292.870 ;
        RECT -27.470 3291.690 -26.290 3292.870 ;
        RECT -29.070 3113.290 -27.890 3114.470 ;
        RECT -27.470 3113.290 -26.290 3114.470 ;
        RECT -29.070 3111.690 -27.890 3112.870 ;
        RECT -27.470 3111.690 -26.290 3112.870 ;
        RECT -29.070 2933.290 -27.890 2934.470 ;
        RECT -27.470 2933.290 -26.290 2934.470 ;
        RECT -29.070 2931.690 -27.890 2932.870 ;
        RECT -27.470 2931.690 -26.290 2932.870 ;
        RECT -29.070 2753.290 -27.890 2754.470 ;
        RECT -27.470 2753.290 -26.290 2754.470 ;
        RECT -29.070 2751.690 -27.890 2752.870 ;
        RECT -27.470 2751.690 -26.290 2752.870 ;
        RECT -29.070 2573.290 -27.890 2574.470 ;
        RECT -27.470 2573.290 -26.290 2574.470 ;
        RECT -29.070 2571.690 -27.890 2572.870 ;
        RECT -27.470 2571.690 -26.290 2572.870 ;
        RECT -29.070 2393.290 -27.890 2394.470 ;
        RECT -27.470 2393.290 -26.290 2394.470 ;
        RECT -29.070 2391.690 -27.890 2392.870 ;
        RECT -27.470 2391.690 -26.290 2392.870 ;
        RECT -29.070 2213.290 -27.890 2214.470 ;
        RECT -27.470 2213.290 -26.290 2214.470 ;
        RECT -29.070 2211.690 -27.890 2212.870 ;
        RECT -27.470 2211.690 -26.290 2212.870 ;
        RECT -29.070 2033.290 -27.890 2034.470 ;
        RECT -27.470 2033.290 -26.290 2034.470 ;
        RECT -29.070 2031.690 -27.890 2032.870 ;
        RECT -27.470 2031.690 -26.290 2032.870 ;
        RECT -29.070 1853.290 -27.890 1854.470 ;
        RECT -27.470 1853.290 -26.290 1854.470 ;
        RECT -29.070 1851.690 -27.890 1852.870 ;
        RECT -27.470 1851.690 -26.290 1852.870 ;
        RECT -29.070 1673.290 -27.890 1674.470 ;
        RECT -27.470 1673.290 -26.290 1674.470 ;
        RECT -29.070 1671.690 -27.890 1672.870 ;
        RECT -27.470 1671.690 -26.290 1672.870 ;
        RECT -29.070 1493.290 -27.890 1494.470 ;
        RECT -27.470 1493.290 -26.290 1494.470 ;
        RECT -29.070 1491.690 -27.890 1492.870 ;
        RECT -27.470 1491.690 -26.290 1492.870 ;
        RECT -29.070 1313.290 -27.890 1314.470 ;
        RECT -27.470 1313.290 -26.290 1314.470 ;
        RECT -29.070 1311.690 -27.890 1312.870 ;
        RECT -27.470 1311.690 -26.290 1312.870 ;
        RECT -29.070 1133.290 -27.890 1134.470 ;
        RECT -27.470 1133.290 -26.290 1134.470 ;
        RECT -29.070 1131.690 -27.890 1132.870 ;
        RECT -27.470 1131.690 -26.290 1132.870 ;
        RECT -29.070 953.290 -27.890 954.470 ;
        RECT -27.470 953.290 -26.290 954.470 ;
        RECT -29.070 951.690 -27.890 952.870 ;
        RECT -27.470 951.690 -26.290 952.870 ;
        RECT -29.070 773.290 -27.890 774.470 ;
        RECT -27.470 773.290 -26.290 774.470 ;
        RECT -29.070 771.690 -27.890 772.870 ;
        RECT -27.470 771.690 -26.290 772.870 ;
        RECT -29.070 593.290 -27.890 594.470 ;
        RECT -27.470 593.290 -26.290 594.470 ;
        RECT -29.070 591.690 -27.890 592.870 ;
        RECT -27.470 591.690 -26.290 592.870 ;
        RECT -29.070 413.290 -27.890 414.470 ;
        RECT -27.470 413.290 -26.290 414.470 ;
        RECT -29.070 411.690 -27.890 412.870 ;
        RECT -27.470 411.690 -26.290 412.870 ;
        RECT -29.070 233.290 -27.890 234.470 ;
        RECT -27.470 233.290 -26.290 234.470 ;
        RECT -29.070 231.690 -27.890 232.870 ;
        RECT -27.470 231.690 -26.290 232.870 ;
        RECT -29.070 53.290 -27.890 54.470 ;
        RECT -27.470 53.290 -26.290 54.470 ;
        RECT -29.070 51.690 -27.890 52.870 ;
        RECT -27.470 51.690 -26.290 52.870 ;
        RECT -29.070 -22.110 -27.890 -20.930 ;
        RECT -27.470 -22.110 -26.290 -20.930 ;
        RECT -29.070 -23.710 -27.890 -22.530 ;
        RECT -27.470 -23.710 -26.290 -22.530 ;
        RECT 46.330 3542.210 47.510 3543.390 ;
        RECT 47.930 3542.210 49.110 3543.390 ;
        RECT 46.330 3540.610 47.510 3541.790 ;
        RECT 47.930 3540.610 49.110 3541.790 ;
        RECT 46.330 3473.290 47.510 3474.470 ;
        RECT 47.930 3473.290 49.110 3474.470 ;
        RECT 46.330 3471.690 47.510 3472.870 ;
        RECT 47.930 3471.690 49.110 3472.870 ;
        RECT 46.330 3293.290 47.510 3294.470 ;
        RECT 47.930 3293.290 49.110 3294.470 ;
        RECT 46.330 3291.690 47.510 3292.870 ;
        RECT 47.930 3291.690 49.110 3292.870 ;
        RECT 46.330 3113.290 47.510 3114.470 ;
        RECT 47.930 3113.290 49.110 3114.470 ;
        RECT 46.330 3111.690 47.510 3112.870 ;
        RECT 47.930 3111.690 49.110 3112.870 ;
        RECT 46.330 2933.290 47.510 2934.470 ;
        RECT 47.930 2933.290 49.110 2934.470 ;
        RECT 46.330 2931.690 47.510 2932.870 ;
        RECT 47.930 2931.690 49.110 2932.870 ;
        RECT 46.330 2753.290 47.510 2754.470 ;
        RECT 47.930 2753.290 49.110 2754.470 ;
        RECT 46.330 2751.690 47.510 2752.870 ;
        RECT 47.930 2751.690 49.110 2752.870 ;
        RECT 46.330 2573.290 47.510 2574.470 ;
        RECT 47.930 2573.290 49.110 2574.470 ;
        RECT 46.330 2571.690 47.510 2572.870 ;
        RECT 47.930 2571.690 49.110 2572.870 ;
        RECT 46.330 2393.290 47.510 2394.470 ;
        RECT 47.930 2393.290 49.110 2394.470 ;
        RECT 46.330 2391.690 47.510 2392.870 ;
        RECT 47.930 2391.690 49.110 2392.870 ;
        RECT 46.330 2213.290 47.510 2214.470 ;
        RECT 47.930 2213.290 49.110 2214.470 ;
        RECT 46.330 2211.690 47.510 2212.870 ;
        RECT 47.930 2211.690 49.110 2212.870 ;
        RECT 46.330 2033.290 47.510 2034.470 ;
        RECT 47.930 2033.290 49.110 2034.470 ;
        RECT 46.330 2031.690 47.510 2032.870 ;
        RECT 47.930 2031.690 49.110 2032.870 ;
        RECT 46.330 1853.290 47.510 1854.470 ;
        RECT 47.930 1853.290 49.110 1854.470 ;
        RECT 46.330 1851.690 47.510 1852.870 ;
        RECT 47.930 1851.690 49.110 1852.870 ;
        RECT 46.330 1673.290 47.510 1674.470 ;
        RECT 47.930 1673.290 49.110 1674.470 ;
        RECT 46.330 1671.690 47.510 1672.870 ;
        RECT 47.930 1671.690 49.110 1672.870 ;
        RECT 46.330 1493.290 47.510 1494.470 ;
        RECT 47.930 1493.290 49.110 1494.470 ;
        RECT 46.330 1491.690 47.510 1492.870 ;
        RECT 47.930 1491.690 49.110 1492.870 ;
        RECT 46.330 1313.290 47.510 1314.470 ;
        RECT 47.930 1313.290 49.110 1314.470 ;
        RECT 46.330 1311.690 47.510 1312.870 ;
        RECT 47.930 1311.690 49.110 1312.870 ;
        RECT 46.330 1133.290 47.510 1134.470 ;
        RECT 47.930 1133.290 49.110 1134.470 ;
        RECT 46.330 1131.690 47.510 1132.870 ;
        RECT 47.930 1131.690 49.110 1132.870 ;
        RECT 226.330 3542.210 227.510 3543.390 ;
        RECT 227.930 3542.210 229.110 3543.390 ;
        RECT 226.330 3540.610 227.510 3541.790 ;
        RECT 227.930 3540.610 229.110 3541.790 ;
        RECT 226.330 3473.290 227.510 3474.470 ;
        RECT 227.930 3473.290 229.110 3474.470 ;
        RECT 226.330 3471.690 227.510 3472.870 ;
        RECT 227.930 3471.690 229.110 3472.870 ;
        RECT 226.330 3293.290 227.510 3294.470 ;
        RECT 227.930 3293.290 229.110 3294.470 ;
        RECT 226.330 3291.690 227.510 3292.870 ;
        RECT 227.930 3291.690 229.110 3292.870 ;
        RECT 226.330 3113.290 227.510 3114.470 ;
        RECT 227.930 3113.290 229.110 3114.470 ;
        RECT 226.330 3111.690 227.510 3112.870 ;
        RECT 227.930 3111.690 229.110 3112.870 ;
        RECT 226.330 2933.290 227.510 2934.470 ;
        RECT 227.930 2933.290 229.110 2934.470 ;
        RECT 226.330 2931.690 227.510 2932.870 ;
        RECT 227.930 2931.690 229.110 2932.870 ;
        RECT 226.330 2753.290 227.510 2754.470 ;
        RECT 227.930 2753.290 229.110 2754.470 ;
        RECT 226.330 2751.690 227.510 2752.870 ;
        RECT 227.930 2751.690 229.110 2752.870 ;
        RECT 226.330 2573.290 227.510 2574.470 ;
        RECT 227.930 2573.290 229.110 2574.470 ;
        RECT 226.330 2571.690 227.510 2572.870 ;
        RECT 227.930 2571.690 229.110 2572.870 ;
        RECT 226.330 2393.290 227.510 2394.470 ;
        RECT 227.930 2393.290 229.110 2394.470 ;
        RECT 226.330 2391.690 227.510 2392.870 ;
        RECT 227.930 2391.690 229.110 2392.870 ;
        RECT 226.330 2213.290 227.510 2214.470 ;
        RECT 227.930 2213.290 229.110 2214.470 ;
        RECT 226.330 2211.690 227.510 2212.870 ;
        RECT 227.930 2211.690 229.110 2212.870 ;
        RECT 226.330 2033.290 227.510 2034.470 ;
        RECT 227.930 2033.290 229.110 2034.470 ;
        RECT 226.330 2031.690 227.510 2032.870 ;
        RECT 227.930 2031.690 229.110 2032.870 ;
        RECT 226.330 1853.290 227.510 1854.470 ;
        RECT 227.930 1853.290 229.110 1854.470 ;
        RECT 226.330 1851.690 227.510 1852.870 ;
        RECT 227.930 1851.690 229.110 1852.870 ;
        RECT 226.330 1673.290 227.510 1674.470 ;
        RECT 227.930 1673.290 229.110 1674.470 ;
        RECT 226.330 1671.690 227.510 1672.870 ;
        RECT 227.930 1671.690 229.110 1672.870 ;
        RECT 226.330 1493.290 227.510 1494.470 ;
        RECT 227.930 1493.290 229.110 1494.470 ;
        RECT 226.330 1491.690 227.510 1492.870 ;
        RECT 227.930 1491.690 229.110 1492.870 ;
        RECT 226.330 1313.290 227.510 1314.470 ;
        RECT 227.930 1313.290 229.110 1314.470 ;
        RECT 226.330 1311.690 227.510 1312.870 ;
        RECT 227.930 1311.690 229.110 1312.870 ;
        RECT 226.330 1133.290 227.510 1134.470 ;
        RECT 227.930 1133.290 229.110 1134.470 ;
        RECT 226.330 1131.690 227.510 1132.870 ;
        RECT 227.930 1131.690 229.110 1132.870 ;
        RECT 406.330 3542.210 407.510 3543.390 ;
        RECT 407.930 3542.210 409.110 3543.390 ;
        RECT 406.330 3540.610 407.510 3541.790 ;
        RECT 407.930 3540.610 409.110 3541.790 ;
        RECT 406.330 3473.290 407.510 3474.470 ;
        RECT 407.930 3473.290 409.110 3474.470 ;
        RECT 406.330 3471.690 407.510 3472.870 ;
        RECT 407.930 3471.690 409.110 3472.870 ;
        RECT 406.330 3293.290 407.510 3294.470 ;
        RECT 407.930 3293.290 409.110 3294.470 ;
        RECT 406.330 3291.690 407.510 3292.870 ;
        RECT 407.930 3291.690 409.110 3292.870 ;
        RECT 406.330 3113.290 407.510 3114.470 ;
        RECT 407.930 3113.290 409.110 3114.470 ;
        RECT 406.330 3111.690 407.510 3112.870 ;
        RECT 407.930 3111.690 409.110 3112.870 ;
        RECT 406.330 2933.290 407.510 2934.470 ;
        RECT 407.930 2933.290 409.110 2934.470 ;
        RECT 406.330 2931.690 407.510 2932.870 ;
        RECT 407.930 2931.690 409.110 2932.870 ;
        RECT 406.330 2753.290 407.510 2754.470 ;
        RECT 407.930 2753.290 409.110 2754.470 ;
        RECT 406.330 2751.690 407.510 2752.870 ;
        RECT 407.930 2751.690 409.110 2752.870 ;
        RECT 406.330 2573.290 407.510 2574.470 ;
        RECT 407.930 2573.290 409.110 2574.470 ;
        RECT 406.330 2571.690 407.510 2572.870 ;
        RECT 407.930 2571.690 409.110 2572.870 ;
        RECT 406.330 2393.290 407.510 2394.470 ;
        RECT 407.930 2393.290 409.110 2394.470 ;
        RECT 406.330 2391.690 407.510 2392.870 ;
        RECT 407.930 2391.690 409.110 2392.870 ;
        RECT 406.330 2213.290 407.510 2214.470 ;
        RECT 407.930 2213.290 409.110 2214.470 ;
        RECT 406.330 2211.690 407.510 2212.870 ;
        RECT 407.930 2211.690 409.110 2212.870 ;
        RECT 406.330 2033.290 407.510 2034.470 ;
        RECT 407.930 2033.290 409.110 2034.470 ;
        RECT 406.330 2031.690 407.510 2032.870 ;
        RECT 407.930 2031.690 409.110 2032.870 ;
        RECT 406.330 1853.290 407.510 1854.470 ;
        RECT 407.930 1853.290 409.110 1854.470 ;
        RECT 406.330 1851.690 407.510 1852.870 ;
        RECT 407.930 1851.690 409.110 1852.870 ;
        RECT 406.330 1673.290 407.510 1674.470 ;
        RECT 407.930 1673.290 409.110 1674.470 ;
        RECT 406.330 1671.690 407.510 1672.870 ;
        RECT 407.930 1671.690 409.110 1672.870 ;
        RECT 406.330 1493.290 407.510 1494.470 ;
        RECT 407.930 1493.290 409.110 1494.470 ;
        RECT 406.330 1491.690 407.510 1492.870 ;
        RECT 407.930 1491.690 409.110 1492.870 ;
        RECT 406.330 1313.290 407.510 1314.470 ;
        RECT 407.930 1313.290 409.110 1314.470 ;
        RECT 406.330 1311.690 407.510 1312.870 ;
        RECT 407.930 1311.690 409.110 1312.870 ;
        RECT 406.330 1133.290 407.510 1134.470 ;
        RECT 407.930 1133.290 409.110 1134.470 ;
        RECT 406.330 1131.690 407.510 1132.870 ;
        RECT 407.930 1131.690 409.110 1132.870 ;
        RECT 586.330 3542.210 587.510 3543.390 ;
        RECT 587.930 3542.210 589.110 3543.390 ;
        RECT 586.330 3540.610 587.510 3541.790 ;
        RECT 587.930 3540.610 589.110 3541.790 ;
        RECT 586.330 3473.290 587.510 3474.470 ;
        RECT 587.930 3473.290 589.110 3474.470 ;
        RECT 586.330 3471.690 587.510 3472.870 ;
        RECT 587.930 3471.690 589.110 3472.870 ;
        RECT 586.330 3293.290 587.510 3294.470 ;
        RECT 587.930 3293.290 589.110 3294.470 ;
        RECT 586.330 3291.690 587.510 3292.870 ;
        RECT 587.930 3291.690 589.110 3292.870 ;
        RECT 586.330 3113.290 587.510 3114.470 ;
        RECT 587.930 3113.290 589.110 3114.470 ;
        RECT 586.330 3111.690 587.510 3112.870 ;
        RECT 587.930 3111.690 589.110 3112.870 ;
        RECT 586.330 2933.290 587.510 2934.470 ;
        RECT 587.930 2933.290 589.110 2934.470 ;
        RECT 586.330 2931.690 587.510 2932.870 ;
        RECT 587.930 2931.690 589.110 2932.870 ;
        RECT 586.330 2753.290 587.510 2754.470 ;
        RECT 587.930 2753.290 589.110 2754.470 ;
        RECT 586.330 2751.690 587.510 2752.870 ;
        RECT 587.930 2751.690 589.110 2752.870 ;
        RECT 586.330 2573.290 587.510 2574.470 ;
        RECT 587.930 2573.290 589.110 2574.470 ;
        RECT 586.330 2571.690 587.510 2572.870 ;
        RECT 587.930 2571.690 589.110 2572.870 ;
        RECT 586.330 2393.290 587.510 2394.470 ;
        RECT 587.930 2393.290 589.110 2394.470 ;
        RECT 586.330 2391.690 587.510 2392.870 ;
        RECT 587.930 2391.690 589.110 2392.870 ;
        RECT 586.330 2213.290 587.510 2214.470 ;
        RECT 587.930 2213.290 589.110 2214.470 ;
        RECT 586.330 2211.690 587.510 2212.870 ;
        RECT 587.930 2211.690 589.110 2212.870 ;
        RECT 586.330 2033.290 587.510 2034.470 ;
        RECT 587.930 2033.290 589.110 2034.470 ;
        RECT 586.330 2031.690 587.510 2032.870 ;
        RECT 587.930 2031.690 589.110 2032.870 ;
        RECT 586.330 1853.290 587.510 1854.470 ;
        RECT 587.930 1853.290 589.110 1854.470 ;
        RECT 586.330 1851.690 587.510 1852.870 ;
        RECT 587.930 1851.690 589.110 1852.870 ;
        RECT 586.330 1673.290 587.510 1674.470 ;
        RECT 587.930 1673.290 589.110 1674.470 ;
        RECT 586.330 1671.690 587.510 1672.870 ;
        RECT 587.930 1671.690 589.110 1672.870 ;
        RECT 586.330 1493.290 587.510 1494.470 ;
        RECT 587.930 1493.290 589.110 1494.470 ;
        RECT 586.330 1491.690 587.510 1492.870 ;
        RECT 587.930 1491.690 589.110 1492.870 ;
        RECT 586.330 1313.290 587.510 1314.470 ;
        RECT 587.930 1313.290 589.110 1314.470 ;
        RECT 586.330 1311.690 587.510 1312.870 ;
        RECT 587.930 1311.690 589.110 1312.870 ;
        RECT 586.330 1133.290 587.510 1134.470 ;
        RECT 587.930 1133.290 589.110 1134.470 ;
        RECT 586.330 1131.690 587.510 1132.870 ;
        RECT 587.930 1131.690 589.110 1132.870 ;
        RECT 766.330 3542.210 767.510 3543.390 ;
        RECT 767.930 3542.210 769.110 3543.390 ;
        RECT 766.330 3540.610 767.510 3541.790 ;
        RECT 767.930 3540.610 769.110 3541.790 ;
        RECT 766.330 3473.290 767.510 3474.470 ;
        RECT 767.930 3473.290 769.110 3474.470 ;
        RECT 766.330 3471.690 767.510 3472.870 ;
        RECT 767.930 3471.690 769.110 3472.870 ;
        RECT 766.330 3293.290 767.510 3294.470 ;
        RECT 767.930 3293.290 769.110 3294.470 ;
        RECT 766.330 3291.690 767.510 3292.870 ;
        RECT 767.930 3291.690 769.110 3292.870 ;
        RECT 766.330 3113.290 767.510 3114.470 ;
        RECT 767.930 3113.290 769.110 3114.470 ;
        RECT 766.330 3111.690 767.510 3112.870 ;
        RECT 767.930 3111.690 769.110 3112.870 ;
        RECT 766.330 2933.290 767.510 2934.470 ;
        RECT 767.930 2933.290 769.110 2934.470 ;
        RECT 766.330 2931.690 767.510 2932.870 ;
        RECT 767.930 2931.690 769.110 2932.870 ;
        RECT 766.330 2753.290 767.510 2754.470 ;
        RECT 767.930 2753.290 769.110 2754.470 ;
        RECT 766.330 2751.690 767.510 2752.870 ;
        RECT 767.930 2751.690 769.110 2752.870 ;
        RECT 766.330 2573.290 767.510 2574.470 ;
        RECT 767.930 2573.290 769.110 2574.470 ;
        RECT 766.330 2571.690 767.510 2572.870 ;
        RECT 767.930 2571.690 769.110 2572.870 ;
        RECT 766.330 2393.290 767.510 2394.470 ;
        RECT 767.930 2393.290 769.110 2394.470 ;
        RECT 766.330 2391.690 767.510 2392.870 ;
        RECT 767.930 2391.690 769.110 2392.870 ;
        RECT 766.330 2213.290 767.510 2214.470 ;
        RECT 767.930 2213.290 769.110 2214.470 ;
        RECT 766.330 2211.690 767.510 2212.870 ;
        RECT 767.930 2211.690 769.110 2212.870 ;
        RECT 766.330 2033.290 767.510 2034.470 ;
        RECT 767.930 2033.290 769.110 2034.470 ;
        RECT 766.330 2031.690 767.510 2032.870 ;
        RECT 767.930 2031.690 769.110 2032.870 ;
        RECT 766.330 1853.290 767.510 1854.470 ;
        RECT 767.930 1853.290 769.110 1854.470 ;
        RECT 766.330 1851.690 767.510 1852.870 ;
        RECT 767.930 1851.690 769.110 1852.870 ;
        RECT 766.330 1673.290 767.510 1674.470 ;
        RECT 767.930 1673.290 769.110 1674.470 ;
        RECT 766.330 1671.690 767.510 1672.870 ;
        RECT 767.930 1671.690 769.110 1672.870 ;
        RECT 766.330 1493.290 767.510 1494.470 ;
        RECT 767.930 1493.290 769.110 1494.470 ;
        RECT 766.330 1491.690 767.510 1492.870 ;
        RECT 767.930 1491.690 769.110 1492.870 ;
        RECT 766.330 1313.290 767.510 1314.470 ;
        RECT 767.930 1313.290 769.110 1314.470 ;
        RECT 766.330 1311.690 767.510 1312.870 ;
        RECT 767.930 1311.690 769.110 1312.870 ;
        RECT 766.330 1133.290 767.510 1134.470 ;
        RECT 767.930 1133.290 769.110 1134.470 ;
        RECT 766.330 1131.690 767.510 1132.870 ;
        RECT 767.930 1131.690 769.110 1132.870 ;
        RECT 946.330 3542.210 947.510 3543.390 ;
        RECT 947.930 3542.210 949.110 3543.390 ;
        RECT 946.330 3540.610 947.510 3541.790 ;
        RECT 947.930 3540.610 949.110 3541.790 ;
        RECT 946.330 3473.290 947.510 3474.470 ;
        RECT 947.930 3473.290 949.110 3474.470 ;
        RECT 946.330 3471.690 947.510 3472.870 ;
        RECT 947.930 3471.690 949.110 3472.870 ;
        RECT 946.330 3293.290 947.510 3294.470 ;
        RECT 947.930 3293.290 949.110 3294.470 ;
        RECT 946.330 3291.690 947.510 3292.870 ;
        RECT 947.930 3291.690 949.110 3292.870 ;
        RECT 946.330 3113.290 947.510 3114.470 ;
        RECT 947.930 3113.290 949.110 3114.470 ;
        RECT 946.330 3111.690 947.510 3112.870 ;
        RECT 947.930 3111.690 949.110 3112.870 ;
        RECT 946.330 2933.290 947.510 2934.470 ;
        RECT 947.930 2933.290 949.110 2934.470 ;
        RECT 946.330 2931.690 947.510 2932.870 ;
        RECT 947.930 2931.690 949.110 2932.870 ;
        RECT 946.330 2753.290 947.510 2754.470 ;
        RECT 947.930 2753.290 949.110 2754.470 ;
        RECT 946.330 2751.690 947.510 2752.870 ;
        RECT 947.930 2751.690 949.110 2752.870 ;
        RECT 946.330 2573.290 947.510 2574.470 ;
        RECT 947.930 2573.290 949.110 2574.470 ;
        RECT 946.330 2571.690 947.510 2572.870 ;
        RECT 947.930 2571.690 949.110 2572.870 ;
        RECT 946.330 2393.290 947.510 2394.470 ;
        RECT 947.930 2393.290 949.110 2394.470 ;
        RECT 946.330 2391.690 947.510 2392.870 ;
        RECT 947.930 2391.690 949.110 2392.870 ;
        RECT 946.330 2213.290 947.510 2214.470 ;
        RECT 947.930 2213.290 949.110 2214.470 ;
        RECT 946.330 2211.690 947.510 2212.870 ;
        RECT 947.930 2211.690 949.110 2212.870 ;
        RECT 946.330 2033.290 947.510 2034.470 ;
        RECT 947.930 2033.290 949.110 2034.470 ;
        RECT 946.330 2031.690 947.510 2032.870 ;
        RECT 947.930 2031.690 949.110 2032.870 ;
        RECT 946.330 1853.290 947.510 1854.470 ;
        RECT 947.930 1853.290 949.110 1854.470 ;
        RECT 946.330 1851.690 947.510 1852.870 ;
        RECT 947.930 1851.690 949.110 1852.870 ;
        RECT 946.330 1673.290 947.510 1674.470 ;
        RECT 947.930 1673.290 949.110 1674.470 ;
        RECT 946.330 1671.690 947.510 1672.870 ;
        RECT 947.930 1671.690 949.110 1672.870 ;
        RECT 946.330 1493.290 947.510 1494.470 ;
        RECT 947.930 1493.290 949.110 1494.470 ;
        RECT 946.330 1491.690 947.510 1492.870 ;
        RECT 947.930 1491.690 949.110 1492.870 ;
        RECT 946.330 1313.290 947.510 1314.470 ;
        RECT 947.930 1313.290 949.110 1314.470 ;
        RECT 946.330 1311.690 947.510 1312.870 ;
        RECT 947.930 1311.690 949.110 1312.870 ;
        RECT 946.330 1133.290 947.510 1134.470 ;
        RECT 947.930 1133.290 949.110 1134.470 ;
        RECT 946.330 1131.690 947.510 1132.870 ;
        RECT 947.930 1131.690 949.110 1132.870 ;
        RECT 1126.330 3542.210 1127.510 3543.390 ;
        RECT 1127.930 3542.210 1129.110 3543.390 ;
        RECT 1126.330 3540.610 1127.510 3541.790 ;
        RECT 1127.930 3540.610 1129.110 3541.790 ;
        RECT 1126.330 3473.290 1127.510 3474.470 ;
        RECT 1127.930 3473.290 1129.110 3474.470 ;
        RECT 1126.330 3471.690 1127.510 3472.870 ;
        RECT 1127.930 3471.690 1129.110 3472.870 ;
        RECT 1126.330 3293.290 1127.510 3294.470 ;
        RECT 1127.930 3293.290 1129.110 3294.470 ;
        RECT 1126.330 3291.690 1127.510 3292.870 ;
        RECT 1127.930 3291.690 1129.110 3292.870 ;
        RECT 1126.330 3113.290 1127.510 3114.470 ;
        RECT 1127.930 3113.290 1129.110 3114.470 ;
        RECT 1126.330 3111.690 1127.510 3112.870 ;
        RECT 1127.930 3111.690 1129.110 3112.870 ;
        RECT 1126.330 2933.290 1127.510 2934.470 ;
        RECT 1127.930 2933.290 1129.110 2934.470 ;
        RECT 1126.330 2931.690 1127.510 2932.870 ;
        RECT 1127.930 2931.690 1129.110 2932.870 ;
        RECT 1126.330 2753.290 1127.510 2754.470 ;
        RECT 1127.930 2753.290 1129.110 2754.470 ;
        RECT 1126.330 2751.690 1127.510 2752.870 ;
        RECT 1127.930 2751.690 1129.110 2752.870 ;
        RECT 1126.330 2573.290 1127.510 2574.470 ;
        RECT 1127.930 2573.290 1129.110 2574.470 ;
        RECT 1126.330 2571.690 1127.510 2572.870 ;
        RECT 1127.930 2571.690 1129.110 2572.870 ;
        RECT 1126.330 2393.290 1127.510 2394.470 ;
        RECT 1127.930 2393.290 1129.110 2394.470 ;
        RECT 1126.330 2391.690 1127.510 2392.870 ;
        RECT 1127.930 2391.690 1129.110 2392.870 ;
        RECT 1126.330 2213.290 1127.510 2214.470 ;
        RECT 1127.930 2213.290 1129.110 2214.470 ;
        RECT 1126.330 2211.690 1127.510 2212.870 ;
        RECT 1127.930 2211.690 1129.110 2212.870 ;
        RECT 1126.330 2033.290 1127.510 2034.470 ;
        RECT 1127.930 2033.290 1129.110 2034.470 ;
        RECT 1126.330 2031.690 1127.510 2032.870 ;
        RECT 1127.930 2031.690 1129.110 2032.870 ;
        RECT 1126.330 1853.290 1127.510 1854.470 ;
        RECT 1127.930 1853.290 1129.110 1854.470 ;
        RECT 1126.330 1851.690 1127.510 1852.870 ;
        RECT 1127.930 1851.690 1129.110 1852.870 ;
        RECT 1126.330 1673.290 1127.510 1674.470 ;
        RECT 1127.930 1673.290 1129.110 1674.470 ;
        RECT 1126.330 1671.690 1127.510 1672.870 ;
        RECT 1127.930 1671.690 1129.110 1672.870 ;
        RECT 1126.330 1493.290 1127.510 1494.470 ;
        RECT 1127.930 1493.290 1129.110 1494.470 ;
        RECT 1126.330 1491.690 1127.510 1492.870 ;
        RECT 1127.930 1491.690 1129.110 1492.870 ;
        RECT 1126.330 1313.290 1127.510 1314.470 ;
        RECT 1127.930 1313.290 1129.110 1314.470 ;
        RECT 1126.330 1311.690 1127.510 1312.870 ;
        RECT 1127.930 1311.690 1129.110 1312.870 ;
        RECT 1126.330 1133.290 1127.510 1134.470 ;
        RECT 1127.930 1133.290 1129.110 1134.470 ;
        RECT 1126.330 1131.690 1127.510 1132.870 ;
        RECT 1127.930 1131.690 1129.110 1132.870 ;
        RECT 46.330 953.290 47.510 954.470 ;
        RECT 47.930 953.290 49.110 954.470 ;
        RECT 46.330 951.690 47.510 952.870 ;
        RECT 47.930 951.690 49.110 952.870 ;
        RECT 46.330 773.290 47.510 774.470 ;
        RECT 47.930 773.290 49.110 774.470 ;
        RECT 46.330 771.690 47.510 772.870 ;
        RECT 47.930 771.690 49.110 772.870 ;
        RECT 46.330 593.290 47.510 594.470 ;
        RECT 47.930 593.290 49.110 594.470 ;
        RECT 46.330 591.690 47.510 592.870 ;
        RECT 47.930 591.690 49.110 592.870 ;
        RECT 46.330 413.290 47.510 414.470 ;
        RECT 47.930 413.290 49.110 414.470 ;
        RECT 46.330 411.690 47.510 412.870 ;
        RECT 47.930 411.690 49.110 412.870 ;
        RECT 1126.330 953.290 1127.510 954.470 ;
        RECT 1127.930 953.290 1129.110 954.470 ;
        RECT 1126.330 951.690 1127.510 952.870 ;
        RECT 1127.930 951.690 1129.110 952.870 ;
        RECT 1126.330 773.290 1127.510 774.470 ;
        RECT 1127.930 773.290 1129.110 774.470 ;
        RECT 1126.330 771.690 1127.510 772.870 ;
        RECT 1127.930 771.690 1129.110 772.870 ;
        RECT 1126.330 593.290 1127.510 594.470 ;
        RECT 1127.930 593.290 1129.110 594.470 ;
        RECT 1126.330 591.690 1127.510 592.870 ;
        RECT 1127.930 591.690 1129.110 592.870 ;
        RECT 1126.330 413.290 1127.510 414.470 ;
        RECT 1127.930 413.290 1129.110 414.470 ;
        RECT 1126.330 411.690 1127.510 412.870 ;
        RECT 1127.930 411.690 1129.110 412.870 ;
        RECT 46.330 233.290 47.510 234.470 ;
        RECT 47.930 233.290 49.110 234.470 ;
        RECT 46.330 231.690 47.510 232.870 ;
        RECT 47.930 231.690 49.110 232.870 ;
        RECT 46.330 53.290 47.510 54.470 ;
        RECT 47.930 53.290 49.110 54.470 ;
        RECT 46.330 51.690 47.510 52.870 ;
        RECT 47.930 51.690 49.110 52.870 ;
        RECT 46.330 -22.110 47.510 -20.930 ;
        RECT 47.930 -22.110 49.110 -20.930 ;
        RECT 46.330 -23.710 47.510 -22.530 ;
        RECT 47.930 -23.710 49.110 -22.530 ;
        RECT 226.330 233.290 227.510 234.470 ;
        RECT 227.930 233.290 229.110 234.470 ;
        RECT 226.330 231.690 227.510 232.870 ;
        RECT 227.930 231.690 229.110 232.870 ;
        RECT 226.330 53.290 227.510 54.470 ;
        RECT 227.930 53.290 229.110 54.470 ;
        RECT 226.330 51.690 227.510 52.870 ;
        RECT 227.930 51.690 229.110 52.870 ;
        RECT 226.330 -22.110 227.510 -20.930 ;
        RECT 227.930 -22.110 229.110 -20.930 ;
        RECT 226.330 -23.710 227.510 -22.530 ;
        RECT 227.930 -23.710 229.110 -22.530 ;
        RECT 406.330 233.290 407.510 234.470 ;
        RECT 407.930 233.290 409.110 234.470 ;
        RECT 406.330 231.690 407.510 232.870 ;
        RECT 407.930 231.690 409.110 232.870 ;
        RECT 406.330 53.290 407.510 54.470 ;
        RECT 407.930 53.290 409.110 54.470 ;
        RECT 406.330 51.690 407.510 52.870 ;
        RECT 407.930 51.690 409.110 52.870 ;
        RECT 406.330 -22.110 407.510 -20.930 ;
        RECT 407.930 -22.110 409.110 -20.930 ;
        RECT 406.330 -23.710 407.510 -22.530 ;
        RECT 407.930 -23.710 409.110 -22.530 ;
        RECT 586.330 233.290 587.510 234.470 ;
        RECT 587.930 233.290 589.110 234.470 ;
        RECT 586.330 231.690 587.510 232.870 ;
        RECT 587.930 231.690 589.110 232.870 ;
        RECT 586.330 53.290 587.510 54.470 ;
        RECT 587.930 53.290 589.110 54.470 ;
        RECT 586.330 51.690 587.510 52.870 ;
        RECT 587.930 51.690 589.110 52.870 ;
        RECT 586.330 -22.110 587.510 -20.930 ;
        RECT 587.930 -22.110 589.110 -20.930 ;
        RECT 586.330 -23.710 587.510 -22.530 ;
        RECT 587.930 -23.710 589.110 -22.530 ;
        RECT 766.330 233.290 767.510 234.470 ;
        RECT 767.930 233.290 769.110 234.470 ;
        RECT 766.330 231.690 767.510 232.870 ;
        RECT 767.930 231.690 769.110 232.870 ;
        RECT 766.330 53.290 767.510 54.470 ;
        RECT 767.930 53.290 769.110 54.470 ;
        RECT 766.330 51.690 767.510 52.870 ;
        RECT 767.930 51.690 769.110 52.870 ;
        RECT 766.330 -22.110 767.510 -20.930 ;
        RECT 767.930 -22.110 769.110 -20.930 ;
        RECT 766.330 -23.710 767.510 -22.530 ;
        RECT 767.930 -23.710 769.110 -22.530 ;
        RECT 946.330 233.290 947.510 234.470 ;
        RECT 947.930 233.290 949.110 234.470 ;
        RECT 946.330 231.690 947.510 232.870 ;
        RECT 947.930 231.690 949.110 232.870 ;
        RECT 946.330 53.290 947.510 54.470 ;
        RECT 947.930 53.290 949.110 54.470 ;
        RECT 946.330 51.690 947.510 52.870 ;
        RECT 947.930 51.690 949.110 52.870 ;
        RECT 946.330 -22.110 947.510 -20.930 ;
        RECT 947.930 -22.110 949.110 -20.930 ;
        RECT 946.330 -23.710 947.510 -22.530 ;
        RECT 947.930 -23.710 949.110 -22.530 ;
        RECT 1126.330 233.290 1127.510 234.470 ;
        RECT 1127.930 233.290 1129.110 234.470 ;
        RECT 1126.330 231.690 1127.510 232.870 ;
        RECT 1127.930 231.690 1129.110 232.870 ;
        RECT 1126.330 53.290 1127.510 54.470 ;
        RECT 1127.930 53.290 1129.110 54.470 ;
        RECT 1126.330 51.690 1127.510 52.870 ;
        RECT 1127.930 51.690 1129.110 52.870 ;
        RECT 1126.330 -22.110 1127.510 -20.930 ;
        RECT 1127.930 -22.110 1129.110 -20.930 ;
        RECT 1126.330 -23.710 1127.510 -22.530 ;
        RECT 1127.930 -23.710 1129.110 -22.530 ;
        RECT 1306.330 3542.210 1307.510 3543.390 ;
        RECT 1307.930 3542.210 1309.110 3543.390 ;
        RECT 1306.330 3540.610 1307.510 3541.790 ;
        RECT 1307.930 3540.610 1309.110 3541.790 ;
        RECT 1306.330 3473.290 1307.510 3474.470 ;
        RECT 1307.930 3473.290 1309.110 3474.470 ;
        RECT 1306.330 3471.690 1307.510 3472.870 ;
        RECT 1307.930 3471.690 1309.110 3472.870 ;
        RECT 1306.330 3293.290 1307.510 3294.470 ;
        RECT 1307.930 3293.290 1309.110 3294.470 ;
        RECT 1306.330 3291.690 1307.510 3292.870 ;
        RECT 1307.930 3291.690 1309.110 3292.870 ;
        RECT 1306.330 3113.290 1307.510 3114.470 ;
        RECT 1307.930 3113.290 1309.110 3114.470 ;
        RECT 1306.330 3111.690 1307.510 3112.870 ;
        RECT 1307.930 3111.690 1309.110 3112.870 ;
        RECT 1306.330 2933.290 1307.510 2934.470 ;
        RECT 1307.930 2933.290 1309.110 2934.470 ;
        RECT 1306.330 2931.690 1307.510 2932.870 ;
        RECT 1307.930 2931.690 1309.110 2932.870 ;
        RECT 1306.330 2753.290 1307.510 2754.470 ;
        RECT 1307.930 2753.290 1309.110 2754.470 ;
        RECT 1306.330 2751.690 1307.510 2752.870 ;
        RECT 1307.930 2751.690 1309.110 2752.870 ;
        RECT 1306.330 2573.290 1307.510 2574.470 ;
        RECT 1307.930 2573.290 1309.110 2574.470 ;
        RECT 1306.330 2571.690 1307.510 2572.870 ;
        RECT 1307.930 2571.690 1309.110 2572.870 ;
        RECT 1306.330 2393.290 1307.510 2394.470 ;
        RECT 1307.930 2393.290 1309.110 2394.470 ;
        RECT 1306.330 2391.690 1307.510 2392.870 ;
        RECT 1307.930 2391.690 1309.110 2392.870 ;
        RECT 1306.330 2213.290 1307.510 2214.470 ;
        RECT 1307.930 2213.290 1309.110 2214.470 ;
        RECT 1306.330 2211.690 1307.510 2212.870 ;
        RECT 1307.930 2211.690 1309.110 2212.870 ;
        RECT 1306.330 2033.290 1307.510 2034.470 ;
        RECT 1307.930 2033.290 1309.110 2034.470 ;
        RECT 1306.330 2031.690 1307.510 2032.870 ;
        RECT 1307.930 2031.690 1309.110 2032.870 ;
        RECT 1306.330 1853.290 1307.510 1854.470 ;
        RECT 1307.930 1853.290 1309.110 1854.470 ;
        RECT 1306.330 1851.690 1307.510 1852.870 ;
        RECT 1307.930 1851.690 1309.110 1852.870 ;
        RECT 1306.330 1673.290 1307.510 1674.470 ;
        RECT 1307.930 1673.290 1309.110 1674.470 ;
        RECT 1306.330 1671.690 1307.510 1672.870 ;
        RECT 1307.930 1671.690 1309.110 1672.870 ;
        RECT 1306.330 1493.290 1307.510 1494.470 ;
        RECT 1307.930 1493.290 1309.110 1494.470 ;
        RECT 1306.330 1491.690 1307.510 1492.870 ;
        RECT 1307.930 1491.690 1309.110 1492.870 ;
        RECT 1306.330 1313.290 1307.510 1314.470 ;
        RECT 1307.930 1313.290 1309.110 1314.470 ;
        RECT 1306.330 1311.690 1307.510 1312.870 ;
        RECT 1307.930 1311.690 1309.110 1312.870 ;
        RECT 1306.330 1133.290 1307.510 1134.470 ;
        RECT 1307.930 1133.290 1309.110 1134.470 ;
        RECT 1306.330 1131.690 1307.510 1132.870 ;
        RECT 1307.930 1131.690 1309.110 1132.870 ;
        RECT 1306.330 953.290 1307.510 954.470 ;
        RECT 1307.930 953.290 1309.110 954.470 ;
        RECT 1306.330 951.690 1307.510 952.870 ;
        RECT 1307.930 951.690 1309.110 952.870 ;
        RECT 1306.330 773.290 1307.510 774.470 ;
        RECT 1307.930 773.290 1309.110 774.470 ;
        RECT 1306.330 771.690 1307.510 772.870 ;
        RECT 1307.930 771.690 1309.110 772.870 ;
        RECT 1306.330 593.290 1307.510 594.470 ;
        RECT 1307.930 593.290 1309.110 594.470 ;
        RECT 1306.330 591.690 1307.510 592.870 ;
        RECT 1307.930 591.690 1309.110 592.870 ;
        RECT 1306.330 413.290 1307.510 414.470 ;
        RECT 1307.930 413.290 1309.110 414.470 ;
        RECT 1306.330 411.690 1307.510 412.870 ;
        RECT 1307.930 411.690 1309.110 412.870 ;
        RECT 1306.330 233.290 1307.510 234.470 ;
        RECT 1307.930 233.290 1309.110 234.470 ;
        RECT 1306.330 231.690 1307.510 232.870 ;
        RECT 1307.930 231.690 1309.110 232.870 ;
        RECT 1306.330 53.290 1307.510 54.470 ;
        RECT 1307.930 53.290 1309.110 54.470 ;
        RECT 1306.330 51.690 1307.510 52.870 ;
        RECT 1307.930 51.690 1309.110 52.870 ;
        RECT 1306.330 -22.110 1307.510 -20.930 ;
        RECT 1307.930 -22.110 1309.110 -20.930 ;
        RECT 1306.330 -23.710 1307.510 -22.530 ;
        RECT 1307.930 -23.710 1309.110 -22.530 ;
        RECT 1486.330 3542.210 1487.510 3543.390 ;
        RECT 1487.930 3542.210 1489.110 3543.390 ;
        RECT 1486.330 3540.610 1487.510 3541.790 ;
        RECT 1487.930 3540.610 1489.110 3541.790 ;
        RECT 1486.330 3473.290 1487.510 3474.470 ;
        RECT 1487.930 3473.290 1489.110 3474.470 ;
        RECT 1486.330 3471.690 1487.510 3472.870 ;
        RECT 1487.930 3471.690 1489.110 3472.870 ;
        RECT 1486.330 3293.290 1487.510 3294.470 ;
        RECT 1487.930 3293.290 1489.110 3294.470 ;
        RECT 1486.330 3291.690 1487.510 3292.870 ;
        RECT 1487.930 3291.690 1489.110 3292.870 ;
        RECT 1486.330 3113.290 1487.510 3114.470 ;
        RECT 1487.930 3113.290 1489.110 3114.470 ;
        RECT 1486.330 3111.690 1487.510 3112.870 ;
        RECT 1487.930 3111.690 1489.110 3112.870 ;
        RECT 1486.330 2933.290 1487.510 2934.470 ;
        RECT 1487.930 2933.290 1489.110 2934.470 ;
        RECT 1486.330 2931.690 1487.510 2932.870 ;
        RECT 1487.930 2931.690 1489.110 2932.870 ;
        RECT 1486.330 2753.290 1487.510 2754.470 ;
        RECT 1487.930 2753.290 1489.110 2754.470 ;
        RECT 1486.330 2751.690 1487.510 2752.870 ;
        RECT 1487.930 2751.690 1489.110 2752.870 ;
        RECT 1486.330 2573.290 1487.510 2574.470 ;
        RECT 1487.930 2573.290 1489.110 2574.470 ;
        RECT 1486.330 2571.690 1487.510 2572.870 ;
        RECT 1487.930 2571.690 1489.110 2572.870 ;
        RECT 1486.330 2393.290 1487.510 2394.470 ;
        RECT 1487.930 2393.290 1489.110 2394.470 ;
        RECT 1486.330 2391.690 1487.510 2392.870 ;
        RECT 1487.930 2391.690 1489.110 2392.870 ;
        RECT 1486.330 2213.290 1487.510 2214.470 ;
        RECT 1487.930 2213.290 1489.110 2214.470 ;
        RECT 1486.330 2211.690 1487.510 2212.870 ;
        RECT 1487.930 2211.690 1489.110 2212.870 ;
        RECT 1486.330 2033.290 1487.510 2034.470 ;
        RECT 1487.930 2033.290 1489.110 2034.470 ;
        RECT 1486.330 2031.690 1487.510 2032.870 ;
        RECT 1487.930 2031.690 1489.110 2032.870 ;
        RECT 1486.330 1853.290 1487.510 1854.470 ;
        RECT 1487.930 1853.290 1489.110 1854.470 ;
        RECT 1486.330 1851.690 1487.510 1852.870 ;
        RECT 1487.930 1851.690 1489.110 1852.870 ;
        RECT 1486.330 1673.290 1487.510 1674.470 ;
        RECT 1487.930 1673.290 1489.110 1674.470 ;
        RECT 1486.330 1671.690 1487.510 1672.870 ;
        RECT 1487.930 1671.690 1489.110 1672.870 ;
        RECT 1486.330 1493.290 1487.510 1494.470 ;
        RECT 1487.930 1493.290 1489.110 1494.470 ;
        RECT 1486.330 1491.690 1487.510 1492.870 ;
        RECT 1487.930 1491.690 1489.110 1492.870 ;
        RECT 1486.330 1313.290 1487.510 1314.470 ;
        RECT 1487.930 1313.290 1489.110 1314.470 ;
        RECT 1486.330 1311.690 1487.510 1312.870 ;
        RECT 1487.930 1311.690 1489.110 1312.870 ;
        RECT 1486.330 1133.290 1487.510 1134.470 ;
        RECT 1487.930 1133.290 1489.110 1134.470 ;
        RECT 1486.330 1131.690 1487.510 1132.870 ;
        RECT 1487.930 1131.690 1489.110 1132.870 ;
        RECT 1486.330 953.290 1487.510 954.470 ;
        RECT 1487.930 953.290 1489.110 954.470 ;
        RECT 1486.330 951.690 1487.510 952.870 ;
        RECT 1487.930 951.690 1489.110 952.870 ;
        RECT 1486.330 773.290 1487.510 774.470 ;
        RECT 1487.930 773.290 1489.110 774.470 ;
        RECT 1486.330 771.690 1487.510 772.870 ;
        RECT 1487.930 771.690 1489.110 772.870 ;
        RECT 1486.330 593.290 1487.510 594.470 ;
        RECT 1487.930 593.290 1489.110 594.470 ;
        RECT 1486.330 591.690 1487.510 592.870 ;
        RECT 1487.930 591.690 1489.110 592.870 ;
        RECT 1486.330 413.290 1487.510 414.470 ;
        RECT 1487.930 413.290 1489.110 414.470 ;
        RECT 1486.330 411.690 1487.510 412.870 ;
        RECT 1487.930 411.690 1489.110 412.870 ;
        RECT 1486.330 233.290 1487.510 234.470 ;
        RECT 1487.930 233.290 1489.110 234.470 ;
        RECT 1486.330 231.690 1487.510 232.870 ;
        RECT 1487.930 231.690 1489.110 232.870 ;
        RECT 1486.330 53.290 1487.510 54.470 ;
        RECT 1487.930 53.290 1489.110 54.470 ;
        RECT 1486.330 51.690 1487.510 52.870 ;
        RECT 1487.930 51.690 1489.110 52.870 ;
        RECT 1486.330 -22.110 1487.510 -20.930 ;
        RECT 1487.930 -22.110 1489.110 -20.930 ;
        RECT 1486.330 -23.710 1487.510 -22.530 ;
        RECT 1487.930 -23.710 1489.110 -22.530 ;
        RECT 1666.330 3542.210 1667.510 3543.390 ;
        RECT 1667.930 3542.210 1669.110 3543.390 ;
        RECT 1666.330 3540.610 1667.510 3541.790 ;
        RECT 1667.930 3540.610 1669.110 3541.790 ;
        RECT 1666.330 3473.290 1667.510 3474.470 ;
        RECT 1667.930 3473.290 1669.110 3474.470 ;
        RECT 1666.330 3471.690 1667.510 3472.870 ;
        RECT 1667.930 3471.690 1669.110 3472.870 ;
        RECT 1666.330 3293.290 1667.510 3294.470 ;
        RECT 1667.930 3293.290 1669.110 3294.470 ;
        RECT 1666.330 3291.690 1667.510 3292.870 ;
        RECT 1667.930 3291.690 1669.110 3292.870 ;
        RECT 1666.330 3113.290 1667.510 3114.470 ;
        RECT 1667.930 3113.290 1669.110 3114.470 ;
        RECT 1666.330 3111.690 1667.510 3112.870 ;
        RECT 1667.930 3111.690 1669.110 3112.870 ;
        RECT 1666.330 2933.290 1667.510 2934.470 ;
        RECT 1667.930 2933.290 1669.110 2934.470 ;
        RECT 1666.330 2931.690 1667.510 2932.870 ;
        RECT 1667.930 2931.690 1669.110 2932.870 ;
        RECT 1666.330 2753.290 1667.510 2754.470 ;
        RECT 1667.930 2753.290 1669.110 2754.470 ;
        RECT 1666.330 2751.690 1667.510 2752.870 ;
        RECT 1667.930 2751.690 1669.110 2752.870 ;
        RECT 1666.330 2573.290 1667.510 2574.470 ;
        RECT 1667.930 2573.290 1669.110 2574.470 ;
        RECT 1666.330 2571.690 1667.510 2572.870 ;
        RECT 1667.930 2571.690 1669.110 2572.870 ;
        RECT 1666.330 2393.290 1667.510 2394.470 ;
        RECT 1667.930 2393.290 1669.110 2394.470 ;
        RECT 1666.330 2391.690 1667.510 2392.870 ;
        RECT 1667.930 2391.690 1669.110 2392.870 ;
        RECT 1666.330 2213.290 1667.510 2214.470 ;
        RECT 1667.930 2213.290 1669.110 2214.470 ;
        RECT 1666.330 2211.690 1667.510 2212.870 ;
        RECT 1667.930 2211.690 1669.110 2212.870 ;
        RECT 1666.330 2033.290 1667.510 2034.470 ;
        RECT 1667.930 2033.290 1669.110 2034.470 ;
        RECT 1666.330 2031.690 1667.510 2032.870 ;
        RECT 1667.930 2031.690 1669.110 2032.870 ;
        RECT 1666.330 1853.290 1667.510 1854.470 ;
        RECT 1667.930 1853.290 1669.110 1854.470 ;
        RECT 1666.330 1851.690 1667.510 1852.870 ;
        RECT 1667.930 1851.690 1669.110 1852.870 ;
        RECT 1666.330 1673.290 1667.510 1674.470 ;
        RECT 1667.930 1673.290 1669.110 1674.470 ;
        RECT 1666.330 1671.690 1667.510 1672.870 ;
        RECT 1667.930 1671.690 1669.110 1672.870 ;
        RECT 1666.330 1493.290 1667.510 1494.470 ;
        RECT 1667.930 1493.290 1669.110 1494.470 ;
        RECT 1666.330 1491.690 1667.510 1492.870 ;
        RECT 1667.930 1491.690 1669.110 1492.870 ;
        RECT 1666.330 1313.290 1667.510 1314.470 ;
        RECT 1667.930 1313.290 1669.110 1314.470 ;
        RECT 1666.330 1311.690 1667.510 1312.870 ;
        RECT 1667.930 1311.690 1669.110 1312.870 ;
        RECT 1666.330 1133.290 1667.510 1134.470 ;
        RECT 1667.930 1133.290 1669.110 1134.470 ;
        RECT 1666.330 1131.690 1667.510 1132.870 ;
        RECT 1667.930 1131.690 1669.110 1132.870 ;
        RECT 1666.330 953.290 1667.510 954.470 ;
        RECT 1667.930 953.290 1669.110 954.470 ;
        RECT 1666.330 951.690 1667.510 952.870 ;
        RECT 1667.930 951.690 1669.110 952.870 ;
        RECT 1666.330 773.290 1667.510 774.470 ;
        RECT 1667.930 773.290 1669.110 774.470 ;
        RECT 1666.330 771.690 1667.510 772.870 ;
        RECT 1667.930 771.690 1669.110 772.870 ;
        RECT 1666.330 593.290 1667.510 594.470 ;
        RECT 1667.930 593.290 1669.110 594.470 ;
        RECT 1666.330 591.690 1667.510 592.870 ;
        RECT 1667.930 591.690 1669.110 592.870 ;
        RECT 1666.330 413.290 1667.510 414.470 ;
        RECT 1667.930 413.290 1669.110 414.470 ;
        RECT 1666.330 411.690 1667.510 412.870 ;
        RECT 1667.930 411.690 1669.110 412.870 ;
        RECT 1666.330 233.290 1667.510 234.470 ;
        RECT 1667.930 233.290 1669.110 234.470 ;
        RECT 1666.330 231.690 1667.510 232.870 ;
        RECT 1667.930 231.690 1669.110 232.870 ;
        RECT 1666.330 53.290 1667.510 54.470 ;
        RECT 1667.930 53.290 1669.110 54.470 ;
        RECT 1666.330 51.690 1667.510 52.870 ;
        RECT 1667.930 51.690 1669.110 52.870 ;
        RECT 1666.330 -22.110 1667.510 -20.930 ;
        RECT 1667.930 -22.110 1669.110 -20.930 ;
        RECT 1666.330 -23.710 1667.510 -22.530 ;
        RECT 1667.930 -23.710 1669.110 -22.530 ;
        RECT 1846.330 3542.210 1847.510 3543.390 ;
        RECT 1847.930 3542.210 1849.110 3543.390 ;
        RECT 1846.330 3540.610 1847.510 3541.790 ;
        RECT 1847.930 3540.610 1849.110 3541.790 ;
        RECT 1846.330 3473.290 1847.510 3474.470 ;
        RECT 1847.930 3473.290 1849.110 3474.470 ;
        RECT 1846.330 3471.690 1847.510 3472.870 ;
        RECT 1847.930 3471.690 1849.110 3472.870 ;
        RECT 1846.330 3293.290 1847.510 3294.470 ;
        RECT 1847.930 3293.290 1849.110 3294.470 ;
        RECT 1846.330 3291.690 1847.510 3292.870 ;
        RECT 1847.930 3291.690 1849.110 3292.870 ;
        RECT 1846.330 3113.290 1847.510 3114.470 ;
        RECT 1847.930 3113.290 1849.110 3114.470 ;
        RECT 1846.330 3111.690 1847.510 3112.870 ;
        RECT 1847.930 3111.690 1849.110 3112.870 ;
        RECT 1846.330 2933.290 1847.510 2934.470 ;
        RECT 1847.930 2933.290 1849.110 2934.470 ;
        RECT 1846.330 2931.690 1847.510 2932.870 ;
        RECT 1847.930 2931.690 1849.110 2932.870 ;
        RECT 1846.330 2753.290 1847.510 2754.470 ;
        RECT 1847.930 2753.290 1849.110 2754.470 ;
        RECT 1846.330 2751.690 1847.510 2752.870 ;
        RECT 1847.930 2751.690 1849.110 2752.870 ;
        RECT 1846.330 2573.290 1847.510 2574.470 ;
        RECT 1847.930 2573.290 1849.110 2574.470 ;
        RECT 1846.330 2571.690 1847.510 2572.870 ;
        RECT 1847.930 2571.690 1849.110 2572.870 ;
        RECT 1846.330 2393.290 1847.510 2394.470 ;
        RECT 1847.930 2393.290 1849.110 2394.470 ;
        RECT 1846.330 2391.690 1847.510 2392.870 ;
        RECT 1847.930 2391.690 1849.110 2392.870 ;
        RECT 1846.330 2213.290 1847.510 2214.470 ;
        RECT 1847.930 2213.290 1849.110 2214.470 ;
        RECT 1846.330 2211.690 1847.510 2212.870 ;
        RECT 1847.930 2211.690 1849.110 2212.870 ;
        RECT 1846.330 2033.290 1847.510 2034.470 ;
        RECT 1847.930 2033.290 1849.110 2034.470 ;
        RECT 1846.330 2031.690 1847.510 2032.870 ;
        RECT 1847.930 2031.690 1849.110 2032.870 ;
        RECT 1846.330 1853.290 1847.510 1854.470 ;
        RECT 1847.930 1853.290 1849.110 1854.470 ;
        RECT 1846.330 1851.690 1847.510 1852.870 ;
        RECT 1847.930 1851.690 1849.110 1852.870 ;
        RECT 1846.330 1673.290 1847.510 1674.470 ;
        RECT 1847.930 1673.290 1849.110 1674.470 ;
        RECT 1846.330 1671.690 1847.510 1672.870 ;
        RECT 1847.930 1671.690 1849.110 1672.870 ;
        RECT 1846.330 1493.290 1847.510 1494.470 ;
        RECT 1847.930 1493.290 1849.110 1494.470 ;
        RECT 1846.330 1491.690 1847.510 1492.870 ;
        RECT 1847.930 1491.690 1849.110 1492.870 ;
        RECT 1846.330 1313.290 1847.510 1314.470 ;
        RECT 1847.930 1313.290 1849.110 1314.470 ;
        RECT 1846.330 1311.690 1847.510 1312.870 ;
        RECT 1847.930 1311.690 1849.110 1312.870 ;
        RECT 1846.330 1133.290 1847.510 1134.470 ;
        RECT 1847.930 1133.290 1849.110 1134.470 ;
        RECT 1846.330 1131.690 1847.510 1132.870 ;
        RECT 1847.930 1131.690 1849.110 1132.870 ;
        RECT 1846.330 953.290 1847.510 954.470 ;
        RECT 1847.930 953.290 1849.110 954.470 ;
        RECT 1846.330 951.690 1847.510 952.870 ;
        RECT 1847.930 951.690 1849.110 952.870 ;
        RECT 1846.330 773.290 1847.510 774.470 ;
        RECT 1847.930 773.290 1849.110 774.470 ;
        RECT 1846.330 771.690 1847.510 772.870 ;
        RECT 1847.930 771.690 1849.110 772.870 ;
        RECT 1846.330 593.290 1847.510 594.470 ;
        RECT 1847.930 593.290 1849.110 594.470 ;
        RECT 1846.330 591.690 1847.510 592.870 ;
        RECT 1847.930 591.690 1849.110 592.870 ;
        RECT 1846.330 413.290 1847.510 414.470 ;
        RECT 1847.930 413.290 1849.110 414.470 ;
        RECT 1846.330 411.690 1847.510 412.870 ;
        RECT 1847.930 411.690 1849.110 412.870 ;
        RECT 1846.330 233.290 1847.510 234.470 ;
        RECT 1847.930 233.290 1849.110 234.470 ;
        RECT 1846.330 231.690 1847.510 232.870 ;
        RECT 1847.930 231.690 1849.110 232.870 ;
        RECT 1846.330 53.290 1847.510 54.470 ;
        RECT 1847.930 53.290 1849.110 54.470 ;
        RECT 1846.330 51.690 1847.510 52.870 ;
        RECT 1847.930 51.690 1849.110 52.870 ;
        RECT 1846.330 -22.110 1847.510 -20.930 ;
        RECT 1847.930 -22.110 1849.110 -20.930 ;
        RECT 1846.330 -23.710 1847.510 -22.530 ;
        RECT 1847.930 -23.710 1849.110 -22.530 ;
        RECT 2026.330 3542.210 2027.510 3543.390 ;
        RECT 2027.930 3542.210 2029.110 3543.390 ;
        RECT 2026.330 3540.610 2027.510 3541.790 ;
        RECT 2027.930 3540.610 2029.110 3541.790 ;
        RECT 2026.330 3473.290 2027.510 3474.470 ;
        RECT 2027.930 3473.290 2029.110 3474.470 ;
        RECT 2026.330 3471.690 2027.510 3472.870 ;
        RECT 2027.930 3471.690 2029.110 3472.870 ;
        RECT 2026.330 3293.290 2027.510 3294.470 ;
        RECT 2027.930 3293.290 2029.110 3294.470 ;
        RECT 2026.330 3291.690 2027.510 3292.870 ;
        RECT 2027.930 3291.690 2029.110 3292.870 ;
        RECT 2026.330 3113.290 2027.510 3114.470 ;
        RECT 2027.930 3113.290 2029.110 3114.470 ;
        RECT 2026.330 3111.690 2027.510 3112.870 ;
        RECT 2027.930 3111.690 2029.110 3112.870 ;
        RECT 2026.330 2933.290 2027.510 2934.470 ;
        RECT 2027.930 2933.290 2029.110 2934.470 ;
        RECT 2026.330 2931.690 2027.510 2932.870 ;
        RECT 2027.930 2931.690 2029.110 2932.870 ;
        RECT 2026.330 2753.290 2027.510 2754.470 ;
        RECT 2027.930 2753.290 2029.110 2754.470 ;
        RECT 2026.330 2751.690 2027.510 2752.870 ;
        RECT 2027.930 2751.690 2029.110 2752.870 ;
        RECT 2026.330 2573.290 2027.510 2574.470 ;
        RECT 2027.930 2573.290 2029.110 2574.470 ;
        RECT 2026.330 2571.690 2027.510 2572.870 ;
        RECT 2027.930 2571.690 2029.110 2572.870 ;
        RECT 2026.330 2393.290 2027.510 2394.470 ;
        RECT 2027.930 2393.290 2029.110 2394.470 ;
        RECT 2026.330 2391.690 2027.510 2392.870 ;
        RECT 2027.930 2391.690 2029.110 2392.870 ;
        RECT 2026.330 2213.290 2027.510 2214.470 ;
        RECT 2027.930 2213.290 2029.110 2214.470 ;
        RECT 2026.330 2211.690 2027.510 2212.870 ;
        RECT 2027.930 2211.690 2029.110 2212.870 ;
        RECT 2026.330 2033.290 2027.510 2034.470 ;
        RECT 2027.930 2033.290 2029.110 2034.470 ;
        RECT 2026.330 2031.690 2027.510 2032.870 ;
        RECT 2027.930 2031.690 2029.110 2032.870 ;
        RECT 2026.330 1853.290 2027.510 1854.470 ;
        RECT 2027.930 1853.290 2029.110 1854.470 ;
        RECT 2026.330 1851.690 2027.510 1852.870 ;
        RECT 2027.930 1851.690 2029.110 1852.870 ;
        RECT 2026.330 1673.290 2027.510 1674.470 ;
        RECT 2027.930 1673.290 2029.110 1674.470 ;
        RECT 2026.330 1671.690 2027.510 1672.870 ;
        RECT 2027.930 1671.690 2029.110 1672.870 ;
        RECT 2026.330 1493.290 2027.510 1494.470 ;
        RECT 2027.930 1493.290 2029.110 1494.470 ;
        RECT 2026.330 1491.690 2027.510 1492.870 ;
        RECT 2027.930 1491.690 2029.110 1492.870 ;
        RECT 2026.330 1313.290 2027.510 1314.470 ;
        RECT 2027.930 1313.290 2029.110 1314.470 ;
        RECT 2026.330 1311.690 2027.510 1312.870 ;
        RECT 2027.930 1311.690 2029.110 1312.870 ;
        RECT 2026.330 1133.290 2027.510 1134.470 ;
        RECT 2027.930 1133.290 2029.110 1134.470 ;
        RECT 2026.330 1131.690 2027.510 1132.870 ;
        RECT 2027.930 1131.690 2029.110 1132.870 ;
        RECT 2026.330 953.290 2027.510 954.470 ;
        RECT 2027.930 953.290 2029.110 954.470 ;
        RECT 2026.330 951.690 2027.510 952.870 ;
        RECT 2027.930 951.690 2029.110 952.870 ;
        RECT 2026.330 773.290 2027.510 774.470 ;
        RECT 2027.930 773.290 2029.110 774.470 ;
        RECT 2026.330 771.690 2027.510 772.870 ;
        RECT 2027.930 771.690 2029.110 772.870 ;
        RECT 2026.330 593.290 2027.510 594.470 ;
        RECT 2027.930 593.290 2029.110 594.470 ;
        RECT 2026.330 591.690 2027.510 592.870 ;
        RECT 2027.930 591.690 2029.110 592.870 ;
        RECT 2026.330 413.290 2027.510 414.470 ;
        RECT 2027.930 413.290 2029.110 414.470 ;
        RECT 2026.330 411.690 2027.510 412.870 ;
        RECT 2027.930 411.690 2029.110 412.870 ;
        RECT 2026.330 233.290 2027.510 234.470 ;
        RECT 2027.930 233.290 2029.110 234.470 ;
        RECT 2026.330 231.690 2027.510 232.870 ;
        RECT 2027.930 231.690 2029.110 232.870 ;
        RECT 2026.330 53.290 2027.510 54.470 ;
        RECT 2027.930 53.290 2029.110 54.470 ;
        RECT 2026.330 51.690 2027.510 52.870 ;
        RECT 2027.930 51.690 2029.110 52.870 ;
        RECT 2026.330 -22.110 2027.510 -20.930 ;
        RECT 2027.930 -22.110 2029.110 -20.930 ;
        RECT 2026.330 -23.710 2027.510 -22.530 ;
        RECT 2027.930 -23.710 2029.110 -22.530 ;
        RECT 2206.330 3542.210 2207.510 3543.390 ;
        RECT 2207.930 3542.210 2209.110 3543.390 ;
        RECT 2206.330 3540.610 2207.510 3541.790 ;
        RECT 2207.930 3540.610 2209.110 3541.790 ;
        RECT 2206.330 3473.290 2207.510 3474.470 ;
        RECT 2207.930 3473.290 2209.110 3474.470 ;
        RECT 2206.330 3471.690 2207.510 3472.870 ;
        RECT 2207.930 3471.690 2209.110 3472.870 ;
        RECT 2206.330 3293.290 2207.510 3294.470 ;
        RECT 2207.930 3293.290 2209.110 3294.470 ;
        RECT 2206.330 3291.690 2207.510 3292.870 ;
        RECT 2207.930 3291.690 2209.110 3292.870 ;
        RECT 2206.330 3113.290 2207.510 3114.470 ;
        RECT 2207.930 3113.290 2209.110 3114.470 ;
        RECT 2206.330 3111.690 2207.510 3112.870 ;
        RECT 2207.930 3111.690 2209.110 3112.870 ;
        RECT 2206.330 2933.290 2207.510 2934.470 ;
        RECT 2207.930 2933.290 2209.110 2934.470 ;
        RECT 2206.330 2931.690 2207.510 2932.870 ;
        RECT 2207.930 2931.690 2209.110 2932.870 ;
        RECT 2206.330 2753.290 2207.510 2754.470 ;
        RECT 2207.930 2753.290 2209.110 2754.470 ;
        RECT 2206.330 2751.690 2207.510 2752.870 ;
        RECT 2207.930 2751.690 2209.110 2752.870 ;
        RECT 2206.330 2573.290 2207.510 2574.470 ;
        RECT 2207.930 2573.290 2209.110 2574.470 ;
        RECT 2206.330 2571.690 2207.510 2572.870 ;
        RECT 2207.930 2571.690 2209.110 2572.870 ;
        RECT 2206.330 2393.290 2207.510 2394.470 ;
        RECT 2207.930 2393.290 2209.110 2394.470 ;
        RECT 2206.330 2391.690 2207.510 2392.870 ;
        RECT 2207.930 2391.690 2209.110 2392.870 ;
        RECT 2206.330 2213.290 2207.510 2214.470 ;
        RECT 2207.930 2213.290 2209.110 2214.470 ;
        RECT 2206.330 2211.690 2207.510 2212.870 ;
        RECT 2207.930 2211.690 2209.110 2212.870 ;
        RECT 2206.330 2033.290 2207.510 2034.470 ;
        RECT 2207.930 2033.290 2209.110 2034.470 ;
        RECT 2206.330 2031.690 2207.510 2032.870 ;
        RECT 2207.930 2031.690 2209.110 2032.870 ;
        RECT 2206.330 1853.290 2207.510 1854.470 ;
        RECT 2207.930 1853.290 2209.110 1854.470 ;
        RECT 2206.330 1851.690 2207.510 1852.870 ;
        RECT 2207.930 1851.690 2209.110 1852.870 ;
        RECT 2206.330 1673.290 2207.510 1674.470 ;
        RECT 2207.930 1673.290 2209.110 1674.470 ;
        RECT 2206.330 1671.690 2207.510 1672.870 ;
        RECT 2207.930 1671.690 2209.110 1672.870 ;
        RECT 2206.330 1493.290 2207.510 1494.470 ;
        RECT 2207.930 1493.290 2209.110 1494.470 ;
        RECT 2206.330 1491.690 2207.510 1492.870 ;
        RECT 2207.930 1491.690 2209.110 1492.870 ;
        RECT 2206.330 1313.290 2207.510 1314.470 ;
        RECT 2207.930 1313.290 2209.110 1314.470 ;
        RECT 2206.330 1311.690 2207.510 1312.870 ;
        RECT 2207.930 1311.690 2209.110 1312.870 ;
        RECT 2206.330 1133.290 2207.510 1134.470 ;
        RECT 2207.930 1133.290 2209.110 1134.470 ;
        RECT 2206.330 1131.690 2207.510 1132.870 ;
        RECT 2207.930 1131.690 2209.110 1132.870 ;
        RECT 2206.330 953.290 2207.510 954.470 ;
        RECT 2207.930 953.290 2209.110 954.470 ;
        RECT 2206.330 951.690 2207.510 952.870 ;
        RECT 2207.930 951.690 2209.110 952.870 ;
        RECT 2206.330 773.290 2207.510 774.470 ;
        RECT 2207.930 773.290 2209.110 774.470 ;
        RECT 2206.330 771.690 2207.510 772.870 ;
        RECT 2207.930 771.690 2209.110 772.870 ;
        RECT 2206.330 593.290 2207.510 594.470 ;
        RECT 2207.930 593.290 2209.110 594.470 ;
        RECT 2206.330 591.690 2207.510 592.870 ;
        RECT 2207.930 591.690 2209.110 592.870 ;
        RECT 2206.330 413.290 2207.510 414.470 ;
        RECT 2207.930 413.290 2209.110 414.470 ;
        RECT 2206.330 411.690 2207.510 412.870 ;
        RECT 2207.930 411.690 2209.110 412.870 ;
        RECT 2206.330 233.290 2207.510 234.470 ;
        RECT 2207.930 233.290 2209.110 234.470 ;
        RECT 2206.330 231.690 2207.510 232.870 ;
        RECT 2207.930 231.690 2209.110 232.870 ;
        RECT 2206.330 53.290 2207.510 54.470 ;
        RECT 2207.930 53.290 2209.110 54.470 ;
        RECT 2206.330 51.690 2207.510 52.870 ;
        RECT 2207.930 51.690 2209.110 52.870 ;
        RECT 2206.330 -22.110 2207.510 -20.930 ;
        RECT 2207.930 -22.110 2209.110 -20.930 ;
        RECT 2206.330 -23.710 2207.510 -22.530 ;
        RECT 2207.930 -23.710 2209.110 -22.530 ;
        RECT 2386.330 3542.210 2387.510 3543.390 ;
        RECT 2387.930 3542.210 2389.110 3543.390 ;
        RECT 2386.330 3540.610 2387.510 3541.790 ;
        RECT 2387.930 3540.610 2389.110 3541.790 ;
        RECT 2386.330 3473.290 2387.510 3474.470 ;
        RECT 2387.930 3473.290 2389.110 3474.470 ;
        RECT 2386.330 3471.690 2387.510 3472.870 ;
        RECT 2387.930 3471.690 2389.110 3472.870 ;
        RECT 2386.330 3293.290 2387.510 3294.470 ;
        RECT 2387.930 3293.290 2389.110 3294.470 ;
        RECT 2386.330 3291.690 2387.510 3292.870 ;
        RECT 2387.930 3291.690 2389.110 3292.870 ;
        RECT 2386.330 3113.290 2387.510 3114.470 ;
        RECT 2387.930 3113.290 2389.110 3114.470 ;
        RECT 2386.330 3111.690 2387.510 3112.870 ;
        RECT 2387.930 3111.690 2389.110 3112.870 ;
        RECT 2386.330 2933.290 2387.510 2934.470 ;
        RECT 2387.930 2933.290 2389.110 2934.470 ;
        RECT 2386.330 2931.690 2387.510 2932.870 ;
        RECT 2387.930 2931.690 2389.110 2932.870 ;
        RECT 2386.330 2753.290 2387.510 2754.470 ;
        RECT 2387.930 2753.290 2389.110 2754.470 ;
        RECT 2386.330 2751.690 2387.510 2752.870 ;
        RECT 2387.930 2751.690 2389.110 2752.870 ;
        RECT 2386.330 2573.290 2387.510 2574.470 ;
        RECT 2387.930 2573.290 2389.110 2574.470 ;
        RECT 2386.330 2571.690 2387.510 2572.870 ;
        RECT 2387.930 2571.690 2389.110 2572.870 ;
        RECT 2386.330 2393.290 2387.510 2394.470 ;
        RECT 2387.930 2393.290 2389.110 2394.470 ;
        RECT 2386.330 2391.690 2387.510 2392.870 ;
        RECT 2387.930 2391.690 2389.110 2392.870 ;
        RECT 2386.330 2213.290 2387.510 2214.470 ;
        RECT 2387.930 2213.290 2389.110 2214.470 ;
        RECT 2386.330 2211.690 2387.510 2212.870 ;
        RECT 2387.930 2211.690 2389.110 2212.870 ;
        RECT 2386.330 2033.290 2387.510 2034.470 ;
        RECT 2387.930 2033.290 2389.110 2034.470 ;
        RECT 2386.330 2031.690 2387.510 2032.870 ;
        RECT 2387.930 2031.690 2389.110 2032.870 ;
        RECT 2386.330 1853.290 2387.510 1854.470 ;
        RECT 2387.930 1853.290 2389.110 1854.470 ;
        RECT 2386.330 1851.690 2387.510 1852.870 ;
        RECT 2387.930 1851.690 2389.110 1852.870 ;
        RECT 2386.330 1673.290 2387.510 1674.470 ;
        RECT 2387.930 1673.290 2389.110 1674.470 ;
        RECT 2386.330 1671.690 2387.510 1672.870 ;
        RECT 2387.930 1671.690 2389.110 1672.870 ;
        RECT 2386.330 1493.290 2387.510 1494.470 ;
        RECT 2387.930 1493.290 2389.110 1494.470 ;
        RECT 2386.330 1491.690 2387.510 1492.870 ;
        RECT 2387.930 1491.690 2389.110 1492.870 ;
        RECT 2386.330 1313.290 2387.510 1314.470 ;
        RECT 2387.930 1313.290 2389.110 1314.470 ;
        RECT 2386.330 1311.690 2387.510 1312.870 ;
        RECT 2387.930 1311.690 2389.110 1312.870 ;
        RECT 2386.330 1133.290 2387.510 1134.470 ;
        RECT 2387.930 1133.290 2389.110 1134.470 ;
        RECT 2386.330 1131.690 2387.510 1132.870 ;
        RECT 2387.930 1131.690 2389.110 1132.870 ;
        RECT 2386.330 953.290 2387.510 954.470 ;
        RECT 2387.930 953.290 2389.110 954.470 ;
        RECT 2386.330 951.690 2387.510 952.870 ;
        RECT 2387.930 951.690 2389.110 952.870 ;
        RECT 2386.330 773.290 2387.510 774.470 ;
        RECT 2387.930 773.290 2389.110 774.470 ;
        RECT 2386.330 771.690 2387.510 772.870 ;
        RECT 2387.930 771.690 2389.110 772.870 ;
        RECT 2386.330 593.290 2387.510 594.470 ;
        RECT 2387.930 593.290 2389.110 594.470 ;
        RECT 2386.330 591.690 2387.510 592.870 ;
        RECT 2387.930 591.690 2389.110 592.870 ;
        RECT 2386.330 413.290 2387.510 414.470 ;
        RECT 2387.930 413.290 2389.110 414.470 ;
        RECT 2386.330 411.690 2387.510 412.870 ;
        RECT 2387.930 411.690 2389.110 412.870 ;
        RECT 2386.330 233.290 2387.510 234.470 ;
        RECT 2387.930 233.290 2389.110 234.470 ;
        RECT 2386.330 231.690 2387.510 232.870 ;
        RECT 2387.930 231.690 2389.110 232.870 ;
        RECT 2386.330 53.290 2387.510 54.470 ;
        RECT 2387.930 53.290 2389.110 54.470 ;
        RECT 2386.330 51.690 2387.510 52.870 ;
        RECT 2387.930 51.690 2389.110 52.870 ;
        RECT 2386.330 -22.110 2387.510 -20.930 ;
        RECT 2387.930 -22.110 2389.110 -20.930 ;
        RECT 2386.330 -23.710 2387.510 -22.530 ;
        RECT 2387.930 -23.710 2389.110 -22.530 ;
        RECT 2566.330 3542.210 2567.510 3543.390 ;
        RECT 2567.930 3542.210 2569.110 3543.390 ;
        RECT 2566.330 3540.610 2567.510 3541.790 ;
        RECT 2567.930 3540.610 2569.110 3541.790 ;
        RECT 2566.330 3473.290 2567.510 3474.470 ;
        RECT 2567.930 3473.290 2569.110 3474.470 ;
        RECT 2566.330 3471.690 2567.510 3472.870 ;
        RECT 2567.930 3471.690 2569.110 3472.870 ;
        RECT 2566.330 3293.290 2567.510 3294.470 ;
        RECT 2567.930 3293.290 2569.110 3294.470 ;
        RECT 2566.330 3291.690 2567.510 3292.870 ;
        RECT 2567.930 3291.690 2569.110 3292.870 ;
        RECT 2566.330 3113.290 2567.510 3114.470 ;
        RECT 2567.930 3113.290 2569.110 3114.470 ;
        RECT 2566.330 3111.690 2567.510 3112.870 ;
        RECT 2567.930 3111.690 2569.110 3112.870 ;
        RECT 2566.330 2933.290 2567.510 2934.470 ;
        RECT 2567.930 2933.290 2569.110 2934.470 ;
        RECT 2566.330 2931.690 2567.510 2932.870 ;
        RECT 2567.930 2931.690 2569.110 2932.870 ;
        RECT 2566.330 2753.290 2567.510 2754.470 ;
        RECT 2567.930 2753.290 2569.110 2754.470 ;
        RECT 2566.330 2751.690 2567.510 2752.870 ;
        RECT 2567.930 2751.690 2569.110 2752.870 ;
        RECT 2566.330 2573.290 2567.510 2574.470 ;
        RECT 2567.930 2573.290 2569.110 2574.470 ;
        RECT 2566.330 2571.690 2567.510 2572.870 ;
        RECT 2567.930 2571.690 2569.110 2572.870 ;
        RECT 2566.330 2393.290 2567.510 2394.470 ;
        RECT 2567.930 2393.290 2569.110 2394.470 ;
        RECT 2566.330 2391.690 2567.510 2392.870 ;
        RECT 2567.930 2391.690 2569.110 2392.870 ;
        RECT 2566.330 2213.290 2567.510 2214.470 ;
        RECT 2567.930 2213.290 2569.110 2214.470 ;
        RECT 2566.330 2211.690 2567.510 2212.870 ;
        RECT 2567.930 2211.690 2569.110 2212.870 ;
        RECT 2566.330 2033.290 2567.510 2034.470 ;
        RECT 2567.930 2033.290 2569.110 2034.470 ;
        RECT 2566.330 2031.690 2567.510 2032.870 ;
        RECT 2567.930 2031.690 2569.110 2032.870 ;
        RECT 2566.330 1853.290 2567.510 1854.470 ;
        RECT 2567.930 1853.290 2569.110 1854.470 ;
        RECT 2566.330 1851.690 2567.510 1852.870 ;
        RECT 2567.930 1851.690 2569.110 1852.870 ;
        RECT 2566.330 1673.290 2567.510 1674.470 ;
        RECT 2567.930 1673.290 2569.110 1674.470 ;
        RECT 2566.330 1671.690 2567.510 1672.870 ;
        RECT 2567.930 1671.690 2569.110 1672.870 ;
        RECT 2566.330 1493.290 2567.510 1494.470 ;
        RECT 2567.930 1493.290 2569.110 1494.470 ;
        RECT 2566.330 1491.690 2567.510 1492.870 ;
        RECT 2567.930 1491.690 2569.110 1492.870 ;
        RECT 2566.330 1313.290 2567.510 1314.470 ;
        RECT 2567.930 1313.290 2569.110 1314.470 ;
        RECT 2566.330 1311.690 2567.510 1312.870 ;
        RECT 2567.930 1311.690 2569.110 1312.870 ;
        RECT 2566.330 1133.290 2567.510 1134.470 ;
        RECT 2567.930 1133.290 2569.110 1134.470 ;
        RECT 2566.330 1131.690 2567.510 1132.870 ;
        RECT 2567.930 1131.690 2569.110 1132.870 ;
        RECT 2566.330 953.290 2567.510 954.470 ;
        RECT 2567.930 953.290 2569.110 954.470 ;
        RECT 2566.330 951.690 2567.510 952.870 ;
        RECT 2567.930 951.690 2569.110 952.870 ;
        RECT 2566.330 773.290 2567.510 774.470 ;
        RECT 2567.930 773.290 2569.110 774.470 ;
        RECT 2566.330 771.690 2567.510 772.870 ;
        RECT 2567.930 771.690 2569.110 772.870 ;
        RECT 2566.330 593.290 2567.510 594.470 ;
        RECT 2567.930 593.290 2569.110 594.470 ;
        RECT 2566.330 591.690 2567.510 592.870 ;
        RECT 2567.930 591.690 2569.110 592.870 ;
        RECT 2566.330 413.290 2567.510 414.470 ;
        RECT 2567.930 413.290 2569.110 414.470 ;
        RECT 2566.330 411.690 2567.510 412.870 ;
        RECT 2567.930 411.690 2569.110 412.870 ;
        RECT 2566.330 233.290 2567.510 234.470 ;
        RECT 2567.930 233.290 2569.110 234.470 ;
        RECT 2566.330 231.690 2567.510 232.870 ;
        RECT 2567.930 231.690 2569.110 232.870 ;
        RECT 2566.330 53.290 2567.510 54.470 ;
        RECT 2567.930 53.290 2569.110 54.470 ;
        RECT 2566.330 51.690 2567.510 52.870 ;
        RECT 2567.930 51.690 2569.110 52.870 ;
        RECT 2566.330 -22.110 2567.510 -20.930 ;
        RECT 2567.930 -22.110 2569.110 -20.930 ;
        RECT 2566.330 -23.710 2567.510 -22.530 ;
        RECT 2567.930 -23.710 2569.110 -22.530 ;
        RECT 2746.330 3542.210 2747.510 3543.390 ;
        RECT 2747.930 3542.210 2749.110 3543.390 ;
        RECT 2746.330 3540.610 2747.510 3541.790 ;
        RECT 2747.930 3540.610 2749.110 3541.790 ;
        RECT 2746.330 3473.290 2747.510 3474.470 ;
        RECT 2747.930 3473.290 2749.110 3474.470 ;
        RECT 2746.330 3471.690 2747.510 3472.870 ;
        RECT 2747.930 3471.690 2749.110 3472.870 ;
        RECT 2746.330 3293.290 2747.510 3294.470 ;
        RECT 2747.930 3293.290 2749.110 3294.470 ;
        RECT 2746.330 3291.690 2747.510 3292.870 ;
        RECT 2747.930 3291.690 2749.110 3292.870 ;
        RECT 2746.330 3113.290 2747.510 3114.470 ;
        RECT 2747.930 3113.290 2749.110 3114.470 ;
        RECT 2746.330 3111.690 2747.510 3112.870 ;
        RECT 2747.930 3111.690 2749.110 3112.870 ;
        RECT 2746.330 2933.290 2747.510 2934.470 ;
        RECT 2747.930 2933.290 2749.110 2934.470 ;
        RECT 2746.330 2931.690 2747.510 2932.870 ;
        RECT 2747.930 2931.690 2749.110 2932.870 ;
        RECT 2746.330 2753.290 2747.510 2754.470 ;
        RECT 2747.930 2753.290 2749.110 2754.470 ;
        RECT 2746.330 2751.690 2747.510 2752.870 ;
        RECT 2747.930 2751.690 2749.110 2752.870 ;
        RECT 2746.330 2573.290 2747.510 2574.470 ;
        RECT 2747.930 2573.290 2749.110 2574.470 ;
        RECT 2746.330 2571.690 2747.510 2572.870 ;
        RECT 2747.930 2571.690 2749.110 2572.870 ;
        RECT 2746.330 2393.290 2747.510 2394.470 ;
        RECT 2747.930 2393.290 2749.110 2394.470 ;
        RECT 2746.330 2391.690 2747.510 2392.870 ;
        RECT 2747.930 2391.690 2749.110 2392.870 ;
        RECT 2746.330 2213.290 2747.510 2214.470 ;
        RECT 2747.930 2213.290 2749.110 2214.470 ;
        RECT 2746.330 2211.690 2747.510 2212.870 ;
        RECT 2747.930 2211.690 2749.110 2212.870 ;
        RECT 2746.330 2033.290 2747.510 2034.470 ;
        RECT 2747.930 2033.290 2749.110 2034.470 ;
        RECT 2746.330 2031.690 2747.510 2032.870 ;
        RECT 2747.930 2031.690 2749.110 2032.870 ;
        RECT 2746.330 1853.290 2747.510 1854.470 ;
        RECT 2747.930 1853.290 2749.110 1854.470 ;
        RECT 2746.330 1851.690 2747.510 1852.870 ;
        RECT 2747.930 1851.690 2749.110 1852.870 ;
        RECT 2746.330 1673.290 2747.510 1674.470 ;
        RECT 2747.930 1673.290 2749.110 1674.470 ;
        RECT 2746.330 1671.690 2747.510 1672.870 ;
        RECT 2747.930 1671.690 2749.110 1672.870 ;
        RECT 2746.330 1493.290 2747.510 1494.470 ;
        RECT 2747.930 1493.290 2749.110 1494.470 ;
        RECT 2746.330 1491.690 2747.510 1492.870 ;
        RECT 2747.930 1491.690 2749.110 1492.870 ;
        RECT 2746.330 1313.290 2747.510 1314.470 ;
        RECT 2747.930 1313.290 2749.110 1314.470 ;
        RECT 2746.330 1311.690 2747.510 1312.870 ;
        RECT 2747.930 1311.690 2749.110 1312.870 ;
        RECT 2746.330 1133.290 2747.510 1134.470 ;
        RECT 2747.930 1133.290 2749.110 1134.470 ;
        RECT 2746.330 1131.690 2747.510 1132.870 ;
        RECT 2747.930 1131.690 2749.110 1132.870 ;
        RECT 2746.330 953.290 2747.510 954.470 ;
        RECT 2747.930 953.290 2749.110 954.470 ;
        RECT 2746.330 951.690 2747.510 952.870 ;
        RECT 2747.930 951.690 2749.110 952.870 ;
        RECT 2746.330 773.290 2747.510 774.470 ;
        RECT 2747.930 773.290 2749.110 774.470 ;
        RECT 2746.330 771.690 2747.510 772.870 ;
        RECT 2747.930 771.690 2749.110 772.870 ;
        RECT 2746.330 593.290 2747.510 594.470 ;
        RECT 2747.930 593.290 2749.110 594.470 ;
        RECT 2746.330 591.690 2747.510 592.870 ;
        RECT 2747.930 591.690 2749.110 592.870 ;
        RECT 2746.330 413.290 2747.510 414.470 ;
        RECT 2747.930 413.290 2749.110 414.470 ;
        RECT 2746.330 411.690 2747.510 412.870 ;
        RECT 2747.930 411.690 2749.110 412.870 ;
        RECT 2746.330 233.290 2747.510 234.470 ;
        RECT 2747.930 233.290 2749.110 234.470 ;
        RECT 2746.330 231.690 2747.510 232.870 ;
        RECT 2747.930 231.690 2749.110 232.870 ;
        RECT 2746.330 53.290 2747.510 54.470 ;
        RECT 2747.930 53.290 2749.110 54.470 ;
        RECT 2746.330 51.690 2747.510 52.870 ;
        RECT 2747.930 51.690 2749.110 52.870 ;
        RECT 2746.330 -22.110 2747.510 -20.930 ;
        RECT 2747.930 -22.110 2749.110 -20.930 ;
        RECT 2746.330 -23.710 2747.510 -22.530 ;
        RECT 2747.930 -23.710 2749.110 -22.530 ;
        RECT 2945.910 3542.210 2947.090 3543.390 ;
        RECT 2947.510 3542.210 2948.690 3543.390 ;
        RECT 2945.910 3540.610 2947.090 3541.790 ;
        RECT 2947.510 3540.610 2948.690 3541.790 ;
        RECT 2945.910 3473.290 2947.090 3474.470 ;
        RECT 2947.510 3473.290 2948.690 3474.470 ;
        RECT 2945.910 3471.690 2947.090 3472.870 ;
        RECT 2947.510 3471.690 2948.690 3472.870 ;
        RECT 2945.910 3293.290 2947.090 3294.470 ;
        RECT 2947.510 3293.290 2948.690 3294.470 ;
        RECT 2945.910 3291.690 2947.090 3292.870 ;
        RECT 2947.510 3291.690 2948.690 3292.870 ;
        RECT 2945.910 3113.290 2947.090 3114.470 ;
        RECT 2947.510 3113.290 2948.690 3114.470 ;
        RECT 2945.910 3111.690 2947.090 3112.870 ;
        RECT 2947.510 3111.690 2948.690 3112.870 ;
        RECT 2945.910 2933.290 2947.090 2934.470 ;
        RECT 2947.510 2933.290 2948.690 2934.470 ;
        RECT 2945.910 2931.690 2947.090 2932.870 ;
        RECT 2947.510 2931.690 2948.690 2932.870 ;
        RECT 2945.910 2753.290 2947.090 2754.470 ;
        RECT 2947.510 2753.290 2948.690 2754.470 ;
        RECT 2945.910 2751.690 2947.090 2752.870 ;
        RECT 2947.510 2751.690 2948.690 2752.870 ;
        RECT 2945.910 2573.290 2947.090 2574.470 ;
        RECT 2947.510 2573.290 2948.690 2574.470 ;
        RECT 2945.910 2571.690 2947.090 2572.870 ;
        RECT 2947.510 2571.690 2948.690 2572.870 ;
        RECT 2945.910 2393.290 2947.090 2394.470 ;
        RECT 2947.510 2393.290 2948.690 2394.470 ;
        RECT 2945.910 2391.690 2947.090 2392.870 ;
        RECT 2947.510 2391.690 2948.690 2392.870 ;
        RECT 2945.910 2213.290 2947.090 2214.470 ;
        RECT 2947.510 2213.290 2948.690 2214.470 ;
        RECT 2945.910 2211.690 2947.090 2212.870 ;
        RECT 2947.510 2211.690 2948.690 2212.870 ;
        RECT 2945.910 2033.290 2947.090 2034.470 ;
        RECT 2947.510 2033.290 2948.690 2034.470 ;
        RECT 2945.910 2031.690 2947.090 2032.870 ;
        RECT 2947.510 2031.690 2948.690 2032.870 ;
        RECT 2945.910 1853.290 2947.090 1854.470 ;
        RECT 2947.510 1853.290 2948.690 1854.470 ;
        RECT 2945.910 1851.690 2947.090 1852.870 ;
        RECT 2947.510 1851.690 2948.690 1852.870 ;
        RECT 2945.910 1673.290 2947.090 1674.470 ;
        RECT 2947.510 1673.290 2948.690 1674.470 ;
        RECT 2945.910 1671.690 2947.090 1672.870 ;
        RECT 2947.510 1671.690 2948.690 1672.870 ;
        RECT 2945.910 1493.290 2947.090 1494.470 ;
        RECT 2947.510 1493.290 2948.690 1494.470 ;
        RECT 2945.910 1491.690 2947.090 1492.870 ;
        RECT 2947.510 1491.690 2948.690 1492.870 ;
        RECT 2945.910 1313.290 2947.090 1314.470 ;
        RECT 2947.510 1313.290 2948.690 1314.470 ;
        RECT 2945.910 1311.690 2947.090 1312.870 ;
        RECT 2947.510 1311.690 2948.690 1312.870 ;
        RECT 2945.910 1133.290 2947.090 1134.470 ;
        RECT 2947.510 1133.290 2948.690 1134.470 ;
        RECT 2945.910 1131.690 2947.090 1132.870 ;
        RECT 2947.510 1131.690 2948.690 1132.870 ;
        RECT 2945.910 953.290 2947.090 954.470 ;
        RECT 2947.510 953.290 2948.690 954.470 ;
        RECT 2945.910 951.690 2947.090 952.870 ;
        RECT 2947.510 951.690 2948.690 952.870 ;
        RECT 2945.910 773.290 2947.090 774.470 ;
        RECT 2947.510 773.290 2948.690 774.470 ;
        RECT 2945.910 771.690 2947.090 772.870 ;
        RECT 2947.510 771.690 2948.690 772.870 ;
        RECT 2945.910 593.290 2947.090 594.470 ;
        RECT 2947.510 593.290 2948.690 594.470 ;
        RECT 2945.910 591.690 2947.090 592.870 ;
        RECT 2947.510 591.690 2948.690 592.870 ;
        RECT 2945.910 413.290 2947.090 414.470 ;
        RECT 2947.510 413.290 2948.690 414.470 ;
        RECT 2945.910 411.690 2947.090 412.870 ;
        RECT 2947.510 411.690 2948.690 412.870 ;
        RECT 2945.910 233.290 2947.090 234.470 ;
        RECT 2947.510 233.290 2948.690 234.470 ;
        RECT 2945.910 231.690 2947.090 232.870 ;
        RECT 2947.510 231.690 2948.690 232.870 ;
        RECT 2945.910 53.290 2947.090 54.470 ;
        RECT 2947.510 53.290 2948.690 54.470 ;
        RECT 2945.910 51.690 2947.090 52.870 ;
        RECT 2947.510 51.690 2948.690 52.870 ;
        RECT 2945.910 -22.110 2947.090 -20.930 ;
        RECT 2947.510 -22.110 2948.690 -20.930 ;
        RECT 2945.910 -23.710 2947.090 -22.530 ;
        RECT 2947.510 -23.710 2948.690 -22.530 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
        RECT -34.030 951.530 2953.650 954.630 ;
        RECT -34.030 771.530 2953.650 774.630 ;
        RECT -34.030 591.530 2953.650 594.630 ;
        RECT -34.030 411.530 2953.650 414.630 ;
        RECT -34.030 231.530 2953.650 234.630 ;
        RECT -34.030 51.530 2953.650 54.630 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
        RECT 244.770 1010.000 247.870 3557.950 ;
        RECT 424.770 1010.000 427.870 3557.950 ;
        RECT 604.770 1010.000 607.870 3557.950 ;
        RECT 784.770 1010.000 787.870 3557.950 ;
        RECT 964.770 1010.000 967.870 3557.950 ;
        RECT 244.770 -38.270 247.870 390.000 ;
        RECT 424.770 -38.270 427.870 390.000 ;
        RECT 604.770 -38.270 607.870 390.000 ;
        RECT 784.770 -38.270 787.870 390.000 ;
        RECT 964.770 -38.270 967.870 390.000 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER via4 ;
        RECT -38.670 3551.810 -37.490 3552.990 ;
        RECT -37.070 3551.810 -35.890 3552.990 ;
        RECT -38.670 3550.210 -37.490 3551.390 ;
        RECT -37.070 3550.210 -35.890 3551.390 ;
        RECT -38.670 3491.890 -37.490 3493.070 ;
        RECT -37.070 3491.890 -35.890 3493.070 ;
        RECT -38.670 3490.290 -37.490 3491.470 ;
        RECT -37.070 3490.290 -35.890 3491.470 ;
        RECT -38.670 3311.890 -37.490 3313.070 ;
        RECT -37.070 3311.890 -35.890 3313.070 ;
        RECT -38.670 3310.290 -37.490 3311.470 ;
        RECT -37.070 3310.290 -35.890 3311.470 ;
        RECT -38.670 3131.890 -37.490 3133.070 ;
        RECT -37.070 3131.890 -35.890 3133.070 ;
        RECT -38.670 3130.290 -37.490 3131.470 ;
        RECT -37.070 3130.290 -35.890 3131.470 ;
        RECT -38.670 2951.890 -37.490 2953.070 ;
        RECT -37.070 2951.890 -35.890 2953.070 ;
        RECT -38.670 2950.290 -37.490 2951.470 ;
        RECT -37.070 2950.290 -35.890 2951.470 ;
        RECT -38.670 2771.890 -37.490 2773.070 ;
        RECT -37.070 2771.890 -35.890 2773.070 ;
        RECT -38.670 2770.290 -37.490 2771.470 ;
        RECT -37.070 2770.290 -35.890 2771.470 ;
        RECT -38.670 2591.890 -37.490 2593.070 ;
        RECT -37.070 2591.890 -35.890 2593.070 ;
        RECT -38.670 2590.290 -37.490 2591.470 ;
        RECT -37.070 2590.290 -35.890 2591.470 ;
        RECT -38.670 2411.890 -37.490 2413.070 ;
        RECT -37.070 2411.890 -35.890 2413.070 ;
        RECT -38.670 2410.290 -37.490 2411.470 ;
        RECT -37.070 2410.290 -35.890 2411.470 ;
        RECT -38.670 2231.890 -37.490 2233.070 ;
        RECT -37.070 2231.890 -35.890 2233.070 ;
        RECT -38.670 2230.290 -37.490 2231.470 ;
        RECT -37.070 2230.290 -35.890 2231.470 ;
        RECT -38.670 2051.890 -37.490 2053.070 ;
        RECT -37.070 2051.890 -35.890 2053.070 ;
        RECT -38.670 2050.290 -37.490 2051.470 ;
        RECT -37.070 2050.290 -35.890 2051.470 ;
        RECT -38.670 1871.890 -37.490 1873.070 ;
        RECT -37.070 1871.890 -35.890 1873.070 ;
        RECT -38.670 1870.290 -37.490 1871.470 ;
        RECT -37.070 1870.290 -35.890 1871.470 ;
        RECT -38.670 1691.890 -37.490 1693.070 ;
        RECT -37.070 1691.890 -35.890 1693.070 ;
        RECT -38.670 1690.290 -37.490 1691.470 ;
        RECT -37.070 1690.290 -35.890 1691.470 ;
        RECT -38.670 1511.890 -37.490 1513.070 ;
        RECT -37.070 1511.890 -35.890 1513.070 ;
        RECT -38.670 1510.290 -37.490 1511.470 ;
        RECT -37.070 1510.290 -35.890 1511.470 ;
        RECT -38.670 1331.890 -37.490 1333.070 ;
        RECT -37.070 1331.890 -35.890 1333.070 ;
        RECT -38.670 1330.290 -37.490 1331.470 ;
        RECT -37.070 1330.290 -35.890 1331.470 ;
        RECT -38.670 1151.890 -37.490 1153.070 ;
        RECT -37.070 1151.890 -35.890 1153.070 ;
        RECT -38.670 1150.290 -37.490 1151.470 ;
        RECT -37.070 1150.290 -35.890 1151.470 ;
        RECT -38.670 971.890 -37.490 973.070 ;
        RECT -37.070 971.890 -35.890 973.070 ;
        RECT -38.670 970.290 -37.490 971.470 ;
        RECT -37.070 970.290 -35.890 971.470 ;
        RECT -38.670 791.890 -37.490 793.070 ;
        RECT -37.070 791.890 -35.890 793.070 ;
        RECT -38.670 790.290 -37.490 791.470 ;
        RECT -37.070 790.290 -35.890 791.470 ;
        RECT -38.670 611.890 -37.490 613.070 ;
        RECT -37.070 611.890 -35.890 613.070 ;
        RECT -38.670 610.290 -37.490 611.470 ;
        RECT -37.070 610.290 -35.890 611.470 ;
        RECT -38.670 431.890 -37.490 433.070 ;
        RECT -37.070 431.890 -35.890 433.070 ;
        RECT -38.670 430.290 -37.490 431.470 ;
        RECT -37.070 430.290 -35.890 431.470 ;
        RECT -38.670 251.890 -37.490 253.070 ;
        RECT -37.070 251.890 -35.890 253.070 ;
        RECT -38.670 250.290 -37.490 251.470 ;
        RECT -37.070 250.290 -35.890 251.470 ;
        RECT -38.670 71.890 -37.490 73.070 ;
        RECT -37.070 71.890 -35.890 73.070 ;
        RECT -38.670 70.290 -37.490 71.470 ;
        RECT -37.070 70.290 -35.890 71.470 ;
        RECT -38.670 -31.710 -37.490 -30.530 ;
        RECT -37.070 -31.710 -35.890 -30.530 ;
        RECT -38.670 -33.310 -37.490 -32.130 ;
        RECT -37.070 -33.310 -35.890 -32.130 ;
        RECT 64.930 3551.810 66.110 3552.990 ;
        RECT 66.530 3551.810 67.710 3552.990 ;
        RECT 64.930 3550.210 66.110 3551.390 ;
        RECT 66.530 3550.210 67.710 3551.390 ;
        RECT 64.930 3491.890 66.110 3493.070 ;
        RECT 66.530 3491.890 67.710 3493.070 ;
        RECT 64.930 3490.290 66.110 3491.470 ;
        RECT 66.530 3490.290 67.710 3491.470 ;
        RECT 64.930 3311.890 66.110 3313.070 ;
        RECT 66.530 3311.890 67.710 3313.070 ;
        RECT 64.930 3310.290 66.110 3311.470 ;
        RECT 66.530 3310.290 67.710 3311.470 ;
        RECT 64.930 3131.890 66.110 3133.070 ;
        RECT 66.530 3131.890 67.710 3133.070 ;
        RECT 64.930 3130.290 66.110 3131.470 ;
        RECT 66.530 3130.290 67.710 3131.470 ;
        RECT 64.930 2951.890 66.110 2953.070 ;
        RECT 66.530 2951.890 67.710 2953.070 ;
        RECT 64.930 2950.290 66.110 2951.470 ;
        RECT 66.530 2950.290 67.710 2951.470 ;
        RECT 64.930 2771.890 66.110 2773.070 ;
        RECT 66.530 2771.890 67.710 2773.070 ;
        RECT 64.930 2770.290 66.110 2771.470 ;
        RECT 66.530 2770.290 67.710 2771.470 ;
        RECT 64.930 2591.890 66.110 2593.070 ;
        RECT 66.530 2591.890 67.710 2593.070 ;
        RECT 64.930 2590.290 66.110 2591.470 ;
        RECT 66.530 2590.290 67.710 2591.470 ;
        RECT 64.930 2411.890 66.110 2413.070 ;
        RECT 66.530 2411.890 67.710 2413.070 ;
        RECT 64.930 2410.290 66.110 2411.470 ;
        RECT 66.530 2410.290 67.710 2411.470 ;
        RECT 64.930 2231.890 66.110 2233.070 ;
        RECT 66.530 2231.890 67.710 2233.070 ;
        RECT 64.930 2230.290 66.110 2231.470 ;
        RECT 66.530 2230.290 67.710 2231.470 ;
        RECT 64.930 2051.890 66.110 2053.070 ;
        RECT 66.530 2051.890 67.710 2053.070 ;
        RECT 64.930 2050.290 66.110 2051.470 ;
        RECT 66.530 2050.290 67.710 2051.470 ;
        RECT 64.930 1871.890 66.110 1873.070 ;
        RECT 66.530 1871.890 67.710 1873.070 ;
        RECT 64.930 1870.290 66.110 1871.470 ;
        RECT 66.530 1870.290 67.710 1871.470 ;
        RECT 64.930 1691.890 66.110 1693.070 ;
        RECT 66.530 1691.890 67.710 1693.070 ;
        RECT 64.930 1690.290 66.110 1691.470 ;
        RECT 66.530 1690.290 67.710 1691.470 ;
        RECT 64.930 1511.890 66.110 1513.070 ;
        RECT 66.530 1511.890 67.710 1513.070 ;
        RECT 64.930 1510.290 66.110 1511.470 ;
        RECT 66.530 1510.290 67.710 1511.470 ;
        RECT 64.930 1331.890 66.110 1333.070 ;
        RECT 66.530 1331.890 67.710 1333.070 ;
        RECT 64.930 1330.290 66.110 1331.470 ;
        RECT 66.530 1330.290 67.710 1331.470 ;
        RECT 64.930 1151.890 66.110 1153.070 ;
        RECT 66.530 1151.890 67.710 1153.070 ;
        RECT 64.930 1150.290 66.110 1151.470 ;
        RECT 66.530 1150.290 67.710 1151.470 ;
        RECT 244.930 3551.810 246.110 3552.990 ;
        RECT 246.530 3551.810 247.710 3552.990 ;
        RECT 244.930 3550.210 246.110 3551.390 ;
        RECT 246.530 3550.210 247.710 3551.390 ;
        RECT 244.930 3491.890 246.110 3493.070 ;
        RECT 246.530 3491.890 247.710 3493.070 ;
        RECT 244.930 3490.290 246.110 3491.470 ;
        RECT 246.530 3490.290 247.710 3491.470 ;
        RECT 244.930 3311.890 246.110 3313.070 ;
        RECT 246.530 3311.890 247.710 3313.070 ;
        RECT 244.930 3310.290 246.110 3311.470 ;
        RECT 246.530 3310.290 247.710 3311.470 ;
        RECT 244.930 3131.890 246.110 3133.070 ;
        RECT 246.530 3131.890 247.710 3133.070 ;
        RECT 244.930 3130.290 246.110 3131.470 ;
        RECT 246.530 3130.290 247.710 3131.470 ;
        RECT 244.930 2951.890 246.110 2953.070 ;
        RECT 246.530 2951.890 247.710 2953.070 ;
        RECT 244.930 2950.290 246.110 2951.470 ;
        RECT 246.530 2950.290 247.710 2951.470 ;
        RECT 244.930 2771.890 246.110 2773.070 ;
        RECT 246.530 2771.890 247.710 2773.070 ;
        RECT 244.930 2770.290 246.110 2771.470 ;
        RECT 246.530 2770.290 247.710 2771.470 ;
        RECT 244.930 2591.890 246.110 2593.070 ;
        RECT 246.530 2591.890 247.710 2593.070 ;
        RECT 244.930 2590.290 246.110 2591.470 ;
        RECT 246.530 2590.290 247.710 2591.470 ;
        RECT 244.930 2411.890 246.110 2413.070 ;
        RECT 246.530 2411.890 247.710 2413.070 ;
        RECT 244.930 2410.290 246.110 2411.470 ;
        RECT 246.530 2410.290 247.710 2411.470 ;
        RECT 244.930 2231.890 246.110 2233.070 ;
        RECT 246.530 2231.890 247.710 2233.070 ;
        RECT 244.930 2230.290 246.110 2231.470 ;
        RECT 246.530 2230.290 247.710 2231.470 ;
        RECT 244.930 2051.890 246.110 2053.070 ;
        RECT 246.530 2051.890 247.710 2053.070 ;
        RECT 244.930 2050.290 246.110 2051.470 ;
        RECT 246.530 2050.290 247.710 2051.470 ;
        RECT 244.930 1871.890 246.110 1873.070 ;
        RECT 246.530 1871.890 247.710 1873.070 ;
        RECT 244.930 1870.290 246.110 1871.470 ;
        RECT 246.530 1870.290 247.710 1871.470 ;
        RECT 244.930 1691.890 246.110 1693.070 ;
        RECT 246.530 1691.890 247.710 1693.070 ;
        RECT 244.930 1690.290 246.110 1691.470 ;
        RECT 246.530 1690.290 247.710 1691.470 ;
        RECT 244.930 1511.890 246.110 1513.070 ;
        RECT 246.530 1511.890 247.710 1513.070 ;
        RECT 244.930 1510.290 246.110 1511.470 ;
        RECT 246.530 1510.290 247.710 1511.470 ;
        RECT 244.930 1331.890 246.110 1333.070 ;
        RECT 246.530 1331.890 247.710 1333.070 ;
        RECT 244.930 1330.290 246.110 1331.470 ;
        RECT 246.530 1330.290 247.710 1331.470 ;
        RECT 244.930 1151.890 246.110 1153.070 ;
        RECT 246.530 1151.890 247.710 1153.070 ;
        RECT 244.930 1150.290 246.110 1151.470 ;
        RECT 246.530 1150.290 247.710 1151.470 ;
        RECT 424.930 3551.810 426.110 3552.990 ;
        RECT 426.530 3551.810 427.710 3552.990 ;
        RECT 424.930 3550.210 426.110 3551.390 ;
        RECT 426.530 3550.210 427.710 3551.390 ;
        RECT 424.930 3491.890 426.110 3493.070 ;
        RECT 426.530 3491.890 427.710 3493.070 ;
        RECT 424.930 3490.290 426.110 3491.470 ;
        RECT 426.530 3490.290 427.710 3491.470 ;
        RECT 424.930 3311.890 426.110 3313.070 ;
        RECT 426.530 3311.890 427.710 3313.070 ;
        RECT 424.930 3310.290 426.110 3311.470 ;
        RECT 426.530 3310.290 427.710 3311.470 ;
        RECT 424.930 3131.890 426.110 3133.070 ;
        RECT 426.530 3131.890 427.710 3133.070 ;
        RECT 424.930 3130.290 426.110 3131.470 ;
        RECT 426.530 3130.290 427.710 3131.470 ;
        RECT 424.930 2951.890 426.110 2953.070 ;
        RECT 426.530 2951.890 427.710 2953.070 ;
        RECT 424.930 2950.290 426.110 2951.470 ;
        RECT 426.530 2950.290 427.710 2951.470 ;
        RECT 424.930 2771.890 426.110 2773.070 ;
        RECT 426.530 2771.890 427.710 2773.070 ;
        RECT 424.930 2770.290 426.110 2771.470 ;
        RECT 426.530 2770.290 427.710 2771.470 ;
        RECT 424.930 2591.890 426.110 2593.070 ;
        RECT 426.530 2591.890 427.710 2593.070 ;
        RECT 424.930 2590.290 426.110 2591.470 ;
        RECT 426.530 2590.290 427.710 2591.470 ;
        RECT 424.930 2411.890 426.110 2413.070 ;
        RECT 426.530 2411.890 427.710 2413.070 ;
        RECT 424.930 2410.290 426.110 2411.470 ;
        RECT 426.530 2410.290 427.710 2411.470 ;
        RECT 424.930 2231.890 426.110 2233.070 ;
        RECT 426.530 2231.890 427.710 2233.070 ;
        RECT 424.930 2230.290 426.110 2231.470 ;
        RECT 426.530 2230.290 427.710 2231.470 ;
        RECT 424.930 2051.890 426.110 2053.070 ;
        RECT 426.530 2051.890 427.710 2053.070 ;
        RECT 424.930 2050.290 426.110 2051.470 ;
        RECT 426.530 2050.290 427.710 2051.470 ;
        RECT 424.930 1871.890 426.110 1873.070 ;
        RECT 426.530 1871.890 427.710 1873.070 ;
        RECT 424.930 1870.290 426.110 1871.470 ;
        RECT 426.530 1870.290 427.710 1871.470 ;
        RECT 424.930 1691.890 426.110 1693.070 ;
        RECT 426.530 1691.890 427.710 1693.070 ;
        RECT 424.930 1690.290 426.110 1691.470 ;
        RECT 426.530 1690.290 427.710 1691.470 ;
        RECT 424.930 1511.890 426.110 1513.070 ;
        RECT 426.530 1511.890 427.710 1513.070 ;
        RECT 424.930 1510.290 426.110 1511.470 ;
        RECT 426.530 1510.290 427.710 1511.470 ;
        RECT 424.930 1331.890 426.110 1333.070 ;
        RECT 426.530 1331.890 427.710 1333.070 ;
        RECT 424.930 1330.290 426.110 1331.470 ;
        RECT 426.530 1330.290 427.710 1331.470 ;
        RECT 424.930 1151.890 426.110 1153.070 ;
        RECT 426.530 1151.890 427.710 1153.070 ;
        RECT 424.930 1150.290 426.110 1151.470 ;
        RECT 426.530 1150.290 427.710 1151.470 ;
        RECT 604.930 3551.810 606.110 3552.990 ;
        RECT 606.530 3551.810 607.710 3552.990 ;
        RECT 604.930 3550.210 606.110 3551.390 ;
        RECT 606.530 3550.210 607.710 3551.390 ;
        RECT 604.930 3491.890 606.110 3493.070 ;
        RECT 606.530 3491.890 607.710 3493.070 ;
        RECT 604.930 3490.290 606.110 3491.470 ;
        RECT 606.530 3490.290 607.710 3491.470 ;
        RECT 604.930 3311.890 606.110 3313.070 ;
        RECT 606.530 3311.890 607.710 3313.070 ;
        RECT 604.930 3310.290 606.110 3311.470 ;
        RECT 606.530 3310.290 607.710 3311.470 ;
        RECT 604.930 3131.890 606.110 3133.070 ;
        RECT 606.530 3131.890 607.710 3133.070 ;
        RECT 604.930 3130.290 606.110 3131.470 ;
        RECT 606.530 3130.290 607.710 3131.470 ;
        RECT 604.930 2951.890 606.110 2953.070 ;
        RECT 606.530 2951.890 607.710 2953.070 ;
        RECT 604.930 2950.290 606.110 2951.470 ;
        RECT 606.530 2950.290 607.710 2951.470 ;
        RECT 604.930 2771.890 606.110 2773.070 ;
        RECT 606.530 2771.890 607.710 2773.070 ;
        RECT 604.930 2770.290 606.110 2771.470 ;
        RECT 606.530 2770.290 607.710 2771.470 ;
        RECT 604.930 2591.890 606.110 2593.070 ;
        RECT 606.530 2591.890 607.710 2593.070 ;
        RECT 604.930 2590.290 606.110 2591.470 ;
        RECT 606.530 2590.290 607.710 2591.470 ;
        RECT 604.930 2411.890 606.110 2413.070 ;
        RECT 606.530 2411.890 607.710 2413.070 ;
        RECT 604.930 2410.290 606.110 2411.470 ;
        RECT 606.530 2410.290 607.710 2411.470 ;
        RECT 604.930 2231.890 606.110 2233.070 ;
        RECT 606.530 2231.890 607.710 2233.070 ;
        RECT 604.930 2230.290 606.110 2231.470 ;
        RECT 606.530 2230.290 607.710 2231.470 ;
        RECT 604.930 2051.890 606.110 2053.070 ;
        RECT 606.530 2051.890 607.710 2053.070 ;
        RECT 604.930 2050.290 606.110 2051.470 ;
        RECT 606.530 2050.290 607.710 2051.470 ;
        RECT 604.930 1871.890 606.110 1873.070 ;
        RECT 606.530 1871.890 607.710 1873.070 ;
        RECT 604.930 1870.290 606.110 1871.470 ;
        RECT 606.530 1870.290 607.710 1871.470 ;
        RECT 604.930 1691.890 606.110 1693.070 ;
        RECT 606.530 1691.890 607.710 1693.070 ;
        RECT 604.930 1690.290 606.110 1691.470 ;
        RECT 606.530 1690.290 607.710 1691.470 ;
        RECT 604.930 1511.890 606.110 1513.070 ;
        RECT 606.530 1511.890 607.710 1513.070 ;
        RECT 604.930 1510.290 606.110 1511.470 ;
        RECT 606.530 1510.290 607.710 1511.470 ;
        RECT 604.930 1331.890 606.110 1333.070 ;
        RECT 606.530 1331.890 607.710 1333.070 ;
        RECT 604.930 1330.290 606.110 1331.470 ;
        RECT 606.530 1330.290 607.710 1331.470 ;
        RECT 604.930 1151.890 606.110 1153.070 ;
        RECT 606.530 1151.890 607.710 1153.070 ;
        RECT 604.930 1150.290 606.110 1151.470 ;
        RECT 606.530 1150.290 607.710 1151.470 ;
        RECT 784.930 3551.810 786.110 3552.990 ;
        RECT 786.530 3551.810 787.710 3552.990 ;
        RECT 784.930 3550.210 786.110 3551.390 ;
        RECT 786.530 3550.210 787.710 3551.390 ;
        RECT 784.930 3491.890 786.110 3493.070 ;
        RECT 786.530 3491.890 787.710 3493.070 ;
        RECT 784.930 3490.290 786.110 3491.470 ;
        RECT 786.530 3490.290 787.710 3491.470 ;
        RECT 784.930 3311.890 786.110 3313.070 ;
        RECT 786.530 3311.890 787.710 3313.070 ;
        RECT 784.930 3310.290 786.110 3311.470 ;
        RECT 786.530 3310.290 787.710 3311.470 ;
        RECT 784.930 3131.890 786.110 3133.070 ;
        RECT 786.530 3131.890 787.710 3133.070 ;
        RECT 784.930 3130.290 786.110 3131.470 ;
        RECT 786.530 3130.290 787.710 3131.470 ;
        RECT 784.930 2951.890 786.110 2953.070 ;
        RECT 786.530 2951.890 787.710 2953.070 ;
        RECT 784.930 2950.290 786.110 2951.470 ;
        RECT 786.530 2950.290 787.710 2951.470 ;
        RECT 784.930 2771.890 786.110 2773.070 ;
        RECT 786.530 2771.890 787.710 2773.070 ;
        RECT 784.930 2770.290 786.110 2771.470 ;
        RECT 786.530 2770.290 787.710 2771.470 ;
        RECT 784.930 2591.890 786.110 2593.070 ;
        RECT 786.530 2591.890 787.710 2593.070 ;
        RECT 784.930 2590.290 786.110 2591.470 ;
        RECT 786.530 2590.290 787.710 2591.470 ;
        RECT 784.930 2411.890 786.110 2413.070 ;
        RECT 786.530 2411.890 787.710 2413.070 ;
        RECT 784.930 2410.290 786.110 2411.470 ;
        RECT 786.530 2410.290 787.710 2411.470 ;
        RECT 784.930 2231.890 786.110 2233.070 ;
        RECT 786.530 2231.890 787.710 2233.070 ;
        RECT 784.930 2230.290 786.110 2231.470 ;
        RECT 786.530 2230.290 787.710 2231.470 ;
        RECT 784.930 2051.890 786.110 2053.070 ;
        RECT 786.530 2051.890 787.710 2053.070 ;
        RECT 784.930 2050.290 786.110 2051.470 ;
        RECT 786.530 2050.290 787.710 2051.470 ;
        RECT 784.930 1871.890 786.110 1873.070 ;
        RECT 786.530 1871.890 787.710 1873.070 ;
        RECT 784.930 1870.290 786.110 1871.470 ;
        RECT 786.530 1870.290 787.710 1871.470 ;
        RECT 784.930 1691.890 786.110 1693.070 ;
        RECT 786.530 1691.890 787.710 1693.070 ;
        RECT 784.930 1690.290 786.110 1691.470 ;
        RECT 786.530 1690.290 787.710 1691.470 ;
        RECT 784.930 1511.890 786.110 1513.070 ;
        RECT 786.530 1511.890 787.710 1513.070 ;
        RECT 784.930 1510.290 786.110 1511.470 ;
        RECT 786.530 1510.290 787.710 1511.470 ;
        RECT 784.930 1331.890 786.110 1333.070 ;
        RECT 786.530 1331.890 787.710 1333.070 ;
        RECT 784.930 1330.290 786.110 1331.470 ;
        RECT 786.530 1330.290 787.710 1331.470 ;
        RECT 784.930 1151.890 786.110 1153.070 ;
        RECT 786.530 1151.890 787.710 1153.070 ;
        RECT 784.930 1150.290 786.110 1151.470 ;
        RECT 786.530 1150.290 787.710 1151.470 ;
        RECT 964.930 3551.810 966.110 3552.990 ;
        RECT 966.530 3551.810 967.710 3552.990 ;
        RECT 964.930 3550.210 966.110 3551.390 ;
        RECT 966.530 3550.210 967.710 3551.390 ;
        RECT 964.930 3491.890 966.110 3493.070 ;
        RECT 966.530 3491.890 967.710 3493.070 ;
        RECT 964.930 3490.290 966.110 3491.470 ;
        RECT 966.530 3490.290 967.710 3491.470 ;
        RECT 964.930 3311.890 966.110 3313.070 ;
        RECT 966.530 3311.890 967.710 3313.070 ;
        RECT 964.930 3310.290 966.110 3311.470 ;
        RECT 966.530 3310.290 967.710 3311.470 ;
        RECT 964.930 3131.890 966.110 3133.070 ;
        RECT 966.530 3131.890 967.710 3133.070 ;
        RECT 964.930 3130.290 966.110 3131.470 ;
        RECT 966.530 3130.290 967.710 3131.470 ;
        RECT 964.930 2951.890 966.110 2953.070 ;
        RECT 966.530 2951.890 967.710 2953.070 ;
        RECT 964.930 2950.290 966.110 2951.470 ;
        RECT 966.530 2950.290 967.710 2951.470 ;
        RECT 964.930 2771.890 966.110 2773.070 ;
        RECT 966.530 2771.890 967.710 2773.070 ;
        RECT 964.930 2770.290 966.110 2771.470 ;
        RECT 966.530 2770.290 967.710 2771.470 ;
        RECT 964.930 2591.890 966.110 2593.070 ;
        RECT 966.530 2591.890 967.710 2593.070 ;
        RECT 964.930 2590.290 966.110 2591.470 ;
        RECT 966.530 2590.290 967.710 2591.470 ;
        RECT 964.930 2411.890 966.110 2413.070 ;
        RECT 966.530 2411.890 967.710 2413.070 ;
        RECT 964.930 2410.290 966.110 2411.470 ;
        RECT 966.530 2410.290 967.710 2411.470 ;
        RECT 964.930 2231.890 966.110 2233.070 ;
        RECT 966.530 2231.890 967.710 2233.070 ;
        RECT 964.930 2230.290 966.110 2231.470 ;
        RECT 966.530 2230.290 967.710 2231.470 ;
        RECT 964.930 2051.890 966.110 2053.070 ;
        RECT 966.530 2051.890 967.710 2053.070 ;
        RECT 964.930 2050.290 966.110 2051.470 ;
        RECT 966.530 2050.290 967.710 2051.470 ;
        RECT 964.930 1871.890 966.110 1873.070 ;
        RECT 966.530 1871.890 967.710 1873.070 ;
        RECT 964.930 1870.290 966.110 1871.470 ;
        RECT 966.530 1870.290 967.710 1871.470 ;
        RECT 964.930 1691.890 966.110 1693.070 ;
        RECT 966.530 1691.890 967.710 1693.070 ;
        RECT 964.930 1690.290 966.110 1691.470 ;
        RECT 966.530 1690.290 967.710 1691.470 ;
        RECT 964.930 1511.890 966.110 1513.070 ;
        RECT 966.530 1511.890 967.710 1513.070 ;
        RECT 964.930 1510.290 966.110 1511.470 ;
        RECT 966.530 1510.290 967.710 1511.470 ;
        RECT 964.930 1331.890 966.110 1333.070 ;
        RECT 966.530 1331.890 967.710 1333.070 ;
        RECT 964.930 1330.290 966.110 1331.470 ;
        RECT 966.530 1330.290 967.710 1331.470 ;
        RECT 964.930 1151.890 966.110 1153.070 ;
        RECT 966.530 1151.890 967.710 1153.070 ;
        RECT 964.930 1150.290 966.110 1151.470 ;
        RECT 966.530 1150.290 967.710 1151.470 ;
        RECT 1144.930 3551.810 1146.110 3552.990 ;
        RECT 1146.530 3551.810 1147.710 3552.990 ;
        RECT 1144.930 3550.210 1146.110 3551.390 ;
        RECT 1146.530 3550.210 1147.710 3551.390 ;
        RECT 1144.930 3491.890 1146.110 3493.070 ;
        RECT 1146.530 3491.890 1147.710 3493.070 ;
        RECT 1144.930 3490.290 1146.110 3491.470 ;
        RECT 1146.530 3490.290 1147.710 3491.470 ;
        RECT 1144.930 3311.890 1146.110 3313.070 ;
        RECT 1146.530 3311.890 1147.710 3313.070 ;
        RECT 1144.930 3310.290 1146.110 3311.470 ;
        RECT 1146.530 3310.290 1147.710 3311.470 ;
        RECT 1144.930 3131.890 1146.110 3133.070 ;
        RECT 1146.530 3131.890 1147.710 3133.070 ;
        RECT 1144.930 3130.290 1146.110 3131.470 ;
        RECT 1146.530 3130.290 1147.710 3131.470 ;
        RECT 1144.930 2951.890 1146.110 2953.070 ;
        RECT 1146.530 2951.890 1147.710 2953.070 ;
        RECT 1144.930 2950.290 1146.110 2951.470 ;
        RECT 1146.530 2950.290 1147.710 2951.470 ;
        RECT 1144.930 2771.890 1146.110 2773.070 ;
        RECT 1146.530 2771.890 1147.710 2773.070 ;
        RECT 1144.930 2770.290 1146.110 2771.470 ;
        RECT 1146.530 2770.290 1147.710 2771.470 ;
        RECT 1144.930 2591.890 1146.110 2593.070 ;
        RECT 1146.530 2591.890 1147.710 2593.070 ;
        RECT 1144.930 2590.290 1146.110 2591.470 ;
        RECT 1146.530 2590.290 1147.710 2591.470 ;
        RECT 1144.930 2411.890 1146.110 2413.070 ;
        RECT 1146.530 2411.890 1147.710 2413.070 ;
        RECT 1144.930 2410.290 1146.110 2411.470 ;
        RECT 1146.530 2410.290 1147.710 2411.470 ;
        RECT 1144.930 2231.890 1146.110 2233.070 ;
        RECT 1146.530 2231.890 1147.710 2233.070 ;
        RECT 1144.930 2230.290 1146.110 2231.470 ;
        RECT 1146.530 2230.290 1147.710 2231.470 ;
        RECT 1144.930 2051.890 1146.110 2053.070 ;
        RECT 1146.530 2051.890 1147.710 2053.070 ;
        RECT 1144.930 2050.290 1146.110 2051.470 ;
        RECT 1146.530 2050.290 1147.710 2051.470 ;
        RECT 1144.930 1871.890 1146.110 1873.070 ;
        RECT 1146.530 1871.890 1147.710 1873.070 ;
        RECT 1144.930 1870.290 1146.110 1871.470 ;
        RECT 1146.530 1870.290 1147.710 1871.470 ;
        RECT 1144.930 1691.890 1146.110 1693.070 ;
        RECT 1146.530 1691.890 1147.710 1693.070 ;
        RECT 1144.930 1690.290 1146.110 1691.470 ;
        RECT 1146.530 1690.290 1147.710 1691.470 ;
        RECT 1144.930 1511.890 1146.110 1513.070 ;
        RECT 1146.530 1511.890 1147.710 1513.070 ;
        RECT 1144.930 1510.290 1146.110 1511.470 ;
        RECT 1146.530 1510.290 1147.710 1511.470 ;
        RECT 1144.930 1331.890 1146.110 1333.070 ;
        RECT 1146.530 1331.890 1147.710 1333.070 ;
        RECT 1144.930 1330.290 1146.110 1331.470 ;
        RECT 1146.530 1330.290 1147.710 1331.470 ;
        RECT 1144.930 1151.890 1146.110 1153.070 ;
        RECT 1146.530 1151.890 1147.710 1153.070 ;
        RECT 1144.930 1150.290 1146.110 1151.470 ;
        RECT 1146.530 1150.290 1147.710 1151.470 ;
        RECT 64.930 971.890 66.110 973.070 ;
        RECT 66.530 971.890 67.710 973.070 ;
        RECT 64.930 970.290 66.110 971.470 ;
        RECT 66.530 970.290 67.710 971.470 ;
        RECT 64.930 791.890 66.110 793.070 ;
        RECT 66.530 791.890 67.710 793.070 ;
        RECT 64.930 790.290 66.110 791.470 ;
        RECT 66.530 790.290 67.710 791.470 ;
        RECT 64.930 611.890 66.110 613.070 ;
        RECT 66.530 611.890 67.710 613.070 ;
        RECT 64.930 610.290 66.110 611.470 ;
        RECT 66.530 610.290 67.710 611.470 ;
        RECT 64.930 431.890 66.110 433.070 ;
        RECT 66.530 431.890 67.710 433.070 ;
        RECT 64.930 430.290 66.110 431.470 ;
        RECT 66.530 430.290 67.710 431.470 ;
        RECT 1144.930 971.890 1146.110 973.070 ;
        RECT 1146.530 971.890 1147.710 973.070 ;
        RECT 1144.930 970.290 1146.110 971.470 ;
        RECT 1146.530 970.290 1147.710 971.470 ;
        RECT 1144.930 791.890 1146.110 793.070 ;
        RECT 1146.530 791.890 1147.710 793.070 ;
        RECT 1144.930 790.290 1146.110 791.470 ;
        RECT 1146.530 790.290 1147.710 791.470 ;
        RECT 1144.930 611.890 1146.110 613.070 ;
        RECT 1146.530 611.890 1147.710 613.070 ;
        RECT 1144.930 610.290 1146.110 611.470 ;
        RECT 1146.530 610.290 1147.710 611.470 ;
        RECT 1144.930 431.890 1146.110 433.070 ;
        RECT 1146.530 431.890 1147.710 433.070 ;
        RECT 1144.930 430.290 1146.110 431.470 ;
        RECT 1146.530 430.290 1147.710 431.470 ;
        RECT 64.930 251.890 66.110 253.070 ;
        RECT 66.530 251.890 67.710 253.070 ;
        RECT 64.930 250.290 66.110 251.470 ;
        RECT 66.530 250.290 67.710 251.470 ;
        RECT 64.930 71.890 66.110 73.070 ;
        RECT 66.530 71.890 67.710 73.070 ;
        RECT 64.930 70.290 66.110 71.470 ;
        RECT 66.530 70.290 67.710 71.470 ;
        RECT 64.930 -31.710 66.110 -30.530 ;
        RECT 66.530 -31.710 67.710 -30.530 ;
        RECT 64.930 -33.310 66.110 -32.130 ;
        RECT 66.530 -33.310 67.710 -32.130 ;
        RECT 244.930 251.890 246.110 253.070 ;
        RECT 246.530 251.890 247.710 253.070 ;
        RECT 244.930 250.290 246.110 251.470 ;
        RECT 246.530 250.290 247.710 251.470 ;
        RECT 244.930 71.890 246.110 73.070 ;
        RECT 246.530 71.890 247.710 73.070 ;
        RECT 244.930 70.290 246.110 71.470 ;
        RECT 246.530 70.290 247.710 71.470 ;
        RECT 244.930 -31.710 246.110 -30.530 ;
        RECT 246.530 -31.710 247.710 -30.530 ;
        RECT 244.930 -33.310 246.110 -32.130 ;
        RECT 246.530 -33.310 247.710 -32.130 ;
        RECT 424.930 251.890 426.110 253.070 ;
        RECT 426.530 251.890 427.710 253.070 ;
        RECT 424.930 250.290 426.110 251.470 ;
        RECT 426.530 250.290 427.710 251.470 ;
        RECT 424.930 71.890 426.110 73.070 ;
        RECT 426.530 71.890 427.710 73.070 ;
        RECT 424.930 70.290 426.110 71.470 ;
        RECT 426.530 70.290 427.710 71.470 ;
        RECT 424.930 -31.710 426.110 -30.530 ;
        RECT 426.530 -31.710 427.710 -30.530 ;
        RECT 424.930 -33.310 426.110 -32.130 ;
        RECT 426.530 -33.310 427.710 -32.130 ;
        RECT 604.930 251.890 606.110 253.070 ;
        RECT 606.530 251.890 607.710 253.070 ;
        RECT 604.930 250.290 606.110 251.470 ;
        RECT 606.530 250.290 607.710 251.470 ;
        RECT 604.930 71.890 606.110 73.070 ;
        RECT 606.530 71.890 607.710 73.070 ;
        RECT 604.930 70.290 606.110 71.470 ;
        RECT 606.530 70.290 607.710 71.470 ;
        RECT 604.930 -31.710 606.110 -30.530 ;
        RECT 606.530 -31.710 607.710 -30.530 ;
        RECT 604.930 -33.310 606.110 -32.130 ;
        RECT 606.530 -33.310 607.710 -32.130 ;
        RECT 784.930 251.890 786.110 253.070 ;
        RECT 786.530 251.890 787.710 253.070 ;
        RECT 784.930 250.290 786.110 251.470 ;
        RECT 786.530 250.290 787.710 251.470 ;
        RECT 784.930 71.890 786.110 73.070 ;
        RECT 786.530 71.890 787.710 73.070 ;
        RECT 784.930 70.290 786.110 71.470 ;
        RECT 786.530 70.290 787.710 71.470 ;
        RECT 784.930 -31.710 786.110 -30.530 ;
        RECT 786.530 -31.710 787.710 -30.530 ;
        RECT 784.930 -33.310 786.110 -32.130 ;
        RECT 786.530 -33.310 787.710 -32.130 ;
        RECT 964.930 251.890 966.110 253.070 ;
        RECT 966.530 251.890 967.710 253.070 ;
        RECT 964.930 250.290 966.110 251.470 ;
        RECT 966.530 250.290 967.710 251.470 ;
        RECT 964.930 71.890 966.110 73.070 ;
        RECT 966.530 71.890 967.710 73.070 ;
        RECT 964.930 70.290 966.110 71.470 ;
        RECT 966.530 70.290 967.710 71.470 ;
        RECT 964.930 -31.710 966.110 -30.530 ;
        RECT 966.530 -31.710 967.710 -30.530 ;
        RECT 964.930 -33.310 966.110 -32.130 ;
        RECT 966.530 -33.310 967.710 -32.130 ;
        RECT 1144.930 251.890 1146.110 253.070 ;
        RECT 1146.530 251.890 1147.710 253.070 ;
        RECT 1144.930 250.290 1146.110 251.470 ;
        RECT 1146.530 250.290 1147.710 251.470 ;
        RECT 1144.930 71.890 1146.110 73.070 ;
        RECT 1146.530 71.890 1147.710 73.070 ;
        RECT 1144.930 70.290 1146.110 71.470 ;
        RECT 1146.530 70.290 1147.710 71.470 ;
        RECT 1144.930 -31.710 1146.110 -30.530 ;
        RECT 1146.530 -31.710 1147.710 -30.530 ;
        RECT 1144.930 -33.310 1146.110 -32.130 ;
        RECT 1146.530 -33.310 1147.710 -32.130 ;
        RECT 1324.930 3551.810 1326.110 3552.990 ;
        RECT 1326.530 3551.810 1327.710 3552.990 ;
        RECT 1324.930 3550.210 1326.110 3551.390 ;
        RECT 1326.530 3550.210 1327.710 3551.390 ;
        RECT 1324.930 3491.890 1326.110 3493.070 ;
        RECT 1326.530 3491.890 1327.710 3493.070 ;
        RECT 1324.930 3490.290 1326.110 3491.470 ;
        RECT 1326.530 3490.290 1327.710 3491.470 ;
        RECT 1324.930 3311.890 1326.110 3313.070 ;
        RECT 1326.530 3311.890 1327.710 3313.070 ;
        RECT 1324.930 3310.290 1326.110 3311.470 ;
        RECT 1326.530 3310.290 1327.710 3311.470 ;
        RECT 1324.930 3131.890 1326.110 3133.070 ;
        RECT 1326.530 3131.890 1327.710 3133.070 ;
        RECT 1324.930 3130.290 1326.110 3131.470 ;
        RECT 1326.530 3130.290 1327.710 3131.470 ;
        RECT 1324.930 2951.890 1326.110 2953.070 ;
        RECT 1326.530 2951.890 1327.710 2953.070 ;
        RECT 1324.930 2950.290 1326.110 2951.470 ;
        RECT 1326.530 2950.290 1327.710 2951.470 ;
        RECT 1324.930 2771.890 1326.110 2773.070 ;
        RECT 1326.530 2771.890 1327.710 2773.070 ;
        RECT 1324.930 2770.290 1326.110 2771.470 ;
        RECT 1326.530 2770.290 1327.710 2771.470 ;
        RECT 1324.930 2591.890 1326.110 2593.070 ;
        RECT 1326.530 2591.890 1327.710 2593.070 ;
        RECT 1324.930 2590.290 1326.110 2591.470 ;
        RECT 1326.530 2590.290 1327.710 2591.470 ;
        RECT 1324.930 2411.890 1326.110 2413.070 ;
        RECT 1326.530 2411.890 1327.710 2413.070 ;
        RECT 1324.930 2410.290 1326.110 2411.470 ;
        RECT 1326.530 2410.290 1327.710 2411.470 ;
        RECT 1324.930 2231.890 1326.110 2233.070 ;
        RECT 1326.530 2231.890 1327.710 2233.070 ;
        RECT 1324.930 2230.290 1326.110 2231.470 ;
        RECT 1326.530 2230.290 1327.710 2231.470 ;
        RECT 1324.930 2051.890 1326.110 2053.070 ;
        RECT 1326.530 2051.890 1327.710 2053.070 ;
        RECT 1324.930 2050.290 1326.110 2051.470 ;
        RECT 1326.530 2050.290 1327.710 2051.470 ;
        RECT 1324.930 1871.890 1326.110 1873.070 ;
        RECT 1326.530 1871.890 1327.710 1873.070 ;
        RECT 1324.930 1870.290 1326.110 1871.470 ;
        RECT 1326.530 1870.290 1327.710 1871.470 ;
        RECT 1324.930 1691.890 1326.110 1693.070 ;
        RECT 1326.530 1691.890 1327.710 1693.070 ;
        RECT 1324.930 1690.290 1326.110 1691.470 ;
        RECT 1326.530 1690.290 1327.710 1691.470 ;
        RECT 1324.930 1511.890 1326.110 1513.070 ;
        RECT 1326.530 1511.890 1327.710 1513.070 ;
        RECT 1324.930 1510.290 1326.110 1511.470 ;
        RECT 1326.530 1510.290 1327.710 1511.470 ;
        RECT 1324.930 1331.890 1326.110 1333.070 ;
        RECT 1326.530 1331.890 1327.710 1333.070 ;
        RECT 1324.930 1330.290 1326.110 1331.470 ;
        RECT 1326.530 1330.290 1327.710 1331.470 ;
        RECT 1324.930 1151.890 1326.110 1153.070 ;
        RECT 1326.530 1151.890 1327.710 1153.070 ;
        RECT 1324.930 1150.290 1326.110 1151.470 ;
        RECT 1326.530 1150.290 1327.710 1151.470 ;
        RECT 1324.930 971.890 1326.110 973.070 ;
        RECT 1326.530 971.890 1327.710 973.070 ;
        RECT 1324.930 970.290 1326.110 971.470 ;
        RECT 1326.530 970.290 1327.710 971.470 ;
        RECT 1324.930 791.890 1326.110 793.070 ;
        RECT 1326.530 791.890 1327.710 793.070 ;
        RECT 1324.930 790.290 1326.110 791.470 ;
        RECT 1326.530 790.290 1327.710 791.470 ;
        RECT 1324.930 611.890 1326.110 613.070 ;
        RECT 1326.530 611.890 1327.710 613.070 ;
        RECT 1324.930 610.290 1326.110 611.470 ;
        RECT 1326.530 610.290 1327.710 611.470 ;
        RECT 1324.930 431.890 1326.110 433.070 ;
        RECT 1326.530 431.890 1327.710 433.070 ;
        RECT 1324.930 430.290 1326.110 431.470 ;
        RECT 1326.530 430.290 1327.710 431.470 ;
        RECT 1324.930 251.890 1326.110 253.070 ;
        RECT 1326.530 251.890 1327.710 253.070 ;
        RECT 1324.930 250.290 1326.110 251.470 ;
        RECT 1326.530 250.290 1327.710 251.470 ;
        RECT 1324.930 71.890 1326.110 73.070 ;
        RECT 1326.530 71.890 1327.710 73.070 ;
        RECT 1324.930 70.290 1326.110 71.470 ;
        RECT 1326.530 70.290 1327.710 71.470 ;
        RECT 1324.930 -31.710 1326.110 -30.530 ;
        RECT 1326.530 -31.710 1327.710 -30.530 ;
        RECT 1324.930 -33.310 1326.110 -32.130 ;
        RECT 1326.530 -33.310 1327.710 -32.130 ;
        RECT 1504.930 3551.810 1506.110 3552.990 ;
        RECT 1506.530 3551.810 1507.710 3552.990 ;
        RECT 1504.930 3550.210 1506.110 3551.390 ;
        RECT 1506.530 3550.210 1507.710 3551.390 ;
        RECT 1504.930 3491.890 1506.110 3493.070 ;
        RECT 1506.530 3491.890 1507.710 3493.070 ;
        RECT 1504.930 3490.290 1506.110 3491.470 ;
        RECT 1506.530 3490.290 1507.710 3491.470 ;
        RECT 1504.930 3311.890 1506.110 3313.070 ;
        RECT 1506.530 3311.890 1507.710 3313.070 ;
        RECT 1504.930 3310.290 1506.110 3311.470 ;
        RECT 1506.530 3310.290 1507.710 3311.470 ;
        RECT 1504.930 3131.890 1506.110 3133.070 ;
        RECT 1506.530 3131.890 1507.710 3133.070 ;
        RECT 1504.930 3130.290 1506.110 3131.470 ;
        RECT 1506.530 3130.290 1507.710 3131.470 ;
        RECT 1504.930 2951.890 1506.110 2953.070 ;
        RECT 1506.530 2951.890 1507.710 2953.070 ;
        RECT 1504.930 2950.290 1506.110 2951.470 ;
        RECT 1506.530 2950.290 1507.710 2951.470 ;
        RECT 1504.930 2771.890 1506.110 2773.070 ;
        RECT 1506.530 2771.890 1507.710 2773.070 ;
        RECT 1504.930 2770.290 1506.110 2771.470 ;
        RECT 1506.530 2770.290 1507.710 2771.470 ;
        RECT 1504.930 2591.890 1506.110 2593.070 ;
        RECT 1506.530 2591.890 1507.710 2593.070 ;
        RECT 1504.930 2590.290 1506.110 2591.470 ;
        RECT 1506.530 2590.290 1507.710 2591.470 ;
        RECT 1504.930 2411.890 1506.110 2413.070 ;
        RECT 1506.530 2411.890 1507.710 2413.070 ;
        RECT 1504.930 2410.290 1506.110 2411.470 ;
        RECT 1506.530 2410.290 1507.710 2411.470 ;
        RECT 1504.930 2231.890 1506.110 2233.070 ;
        RECT 1506.530 2231.890 1507.710 2233.070 ;
        RECT 1504.930 2230.290 1506.110 2231.470 ;
        RECT 1506.530 2230.290 1507.710 2231.470 ;
        RECT 1504.930 2051.890 1506.110 2053.070 ;
        RECT 1506.530 2051.890 1507.710 2053.070 ;
        RECT 1504.930 2050.290 1506.110 2051.470 ;
        RECT 1506.530 2050.290 1507.710 2051.470 ;
        RECT 1504.930 1871.890 1506.110 1873.070 ;
        RECT 1506.530 1871.890 1507.710 1873.070 ;
        RECT 1504.930 1870.290 1506.110 1871.470 ;
        RECT 1506.530 1870.290 1507.710 1871.470 ;
        RECT 1504.930 1691.890 1506.110 1693.070 ;
        RECT 1506.530 1691.890 1507.710 1693.070 ;
        RECT 1504.930 1690.290 1506.110 1691.470 ;
        RECT 1506.530 1690.290 1507.710 1691.470 ;
        RECT 1504.930 1511.890 1506.110 1513.070 ;
        RECT 1506.530 1511.890 1507.710 1513.070 ;
        RECT 1504.930 1510.290 1506.110 1511.470 ;
        RECT 1506.530 1510.290 1507.710 1511.470 ;
        RECT 1504.930 1331.890 1506.110 1333.070 ;
        RECT 1506.530 1331.890 1507.710 1333.070 ;
        RECT 1504.930 1330.290 1506.110 1331.470 ;
        RECT 1506.530 1330.290 1507.710 1331.470 ;
        RECT 1504.930 1151.890 1506.110 1153.070 ;
        RECT 1506.530 1151.890 1507.710 1153.070 ;
        RECT 1504.930 1150.290 1506.110 1151.470 ;
        RECT 1506.530 1150.290 1507.710 1151.470 ;
        RECT 1504.930 971.890 1506.110 973.070 ;
        RECT 1506.530 971.890 1507.710 973.070 ;
        RECT 1504.930 970.290 1506.110 971.470 ;
        RECT 1506.530 970.290 1507.710 971.470 ;
        RECT 1504.930 791.890 1506.110 793.070 ;
        RECT 1506.530 791.890 1507.710 793.070 ;
        RECT 1504.930 790.290 1506.110 791.470 ;
        RECT 1506.530 790.290 1507.710 791.470 ;
        RECT 1504.930 611.890 1506.110 613.070 ;
        RECT 1506.530 611.890 1507.710 613.070 ;
        RECT 1504.930 610.290 1506.110 611.470 ;
        RECT 1506.530 610.290 1507.710 611.470 ;
        RECT 1504.930 431.890 1506.110 433.070 ;
        RECT 1506.530 431.890 1507.710 433.070 ;
        RECT 1504.930 430.290 1506.110 431.470 ;
        RECT 1506.530 430.290 1507.710 431.470 ;
        RECT 1504.930 251.890 1506.110 253.070 ;
        RECT 1506.530 251.890 1507.710 253.070 ;
        RECT 1504.930 250.290 1506.110 251.470 ;
        RECT 1506.530 250.290 1507.710 251.470 ;
        RECT 1504.930 71.890 1506.110 73.070 ;
        RECT 1506.530 71.890 1507.710 73.070 ;
        RECT 1504.930 70.290 1506.110 71.470 ;
        RECT 1506.530 70.290 1507.710 71.470 ;
        RECT 1504.930 -31.710 1506.110 -30.530 ;
        RECT 1506.530 -31.710 1507.710 -30.530 ;
        RECT 1504.930 -33.310 1506.110 -32.130 ;
        RECT 1506.530 -33.310 1507.710 -32.130 ;
        RECT 1684.930 3551.810 1686.110 3552.990 ;
        RECT 1686.530 3551.810 1687.710 3552.990 ;
        RECT 1684.930 3550.210 1686.110 3551.390 ;
        RECT 1686.530 3550.210 1687.710 3551.390 ;
        RECT 1684.930 3491.890 1686.110 3493.070 ;
        RECT 1686.530 3491.890 1687.710 3493.070 ;
        RECT 1684.930 3490.290 1686.110 3491.470 ;
        RECT 1686.530 3490.290 1687.710 3491.470 ;
        RECT 1684.930 3311.890 1686.110 3313.070 ;
        RECT 1686.530 3311.890 1687.710 3313.070 ;
        RECT 1684.930 3310.290 1686.110 3311.470 ;
        RECT 1686.530 3310.290 1687.710 3311.470 ;
        RECT 1684.930 3131.890 1686.110 3133.070 ;
        RECT 1686.530 3131.890 1687.710 3133.070 ;
        RECT 1684.930 3130.290 1686.110 3131.470 ;
        RECT 1686.530 3130.290 1687.710 3131.470 ;
        RECT 1684.930 2951.890 1686.110 2953.070 ;
        RECT 1686.530 2951.890 1687.710 2953.070 ;
        RECT 1684.930 2950.290 1686.110 2951.470 ;
        RECT 1686.530 2950.290 1687.710 2951.470 ;
        RECT 1684.930 2771.890 1686.110 2773.070 ;
        RECT 1686.530 2771.890 1687.710 2773.070 ;
        RECT 1684.930 2770.290 1686.110 2771.470 ;
        RECT 1686.530 2770.290 1687.710 2771.470 ;
        RECT 1684.930 2591.890 1686.110 2593.070 ;
        RECT 1686.530 2591.890 1687.710 2593.070 ;
        RECT 1684.930 2590.290 1686.110 2591.470 ;
        RECT 1686.530 2590.290 1687.710 2591.470 ;
        RECT 1684.930 2411.890 1686.110 2413.070 ;
        RECT 1686.530 2411.890 1687.710 2413.070 ;
        RECT 1684.930 2410.290 1686.110 2411.470 ;
        RECT 1686.530 2410.290 1687.710 2411.470 ;
        RECT 1684.930 2231.890 1686.110 2233.070 ;
        RECT 1686.530 2231.890 1687.710 2233.070 ;
        RECT 1684.930 2230.290 1686.110 2231.470 ;
        RECT 1686.530 2230.290 1687.710 2231.470 ;
        RECT 1684.930 2051.890 1686.110 2053.070 ;
        RECT 1686.530 2051.890 1687.710 2053.070 ;
        RECT 1684.930 2050.290 1686.110 2051.470 ;
        RECT 1686.530 2050.290 1687.710 2051.470 ;
        RECT 1684.930 1871.890 1686.110 1873.070 ;
        RECT 1686.530 1871.890 1687.710 1873.070 ;
        RECT 1684.930 1870.290 1686.110 1871.470 ;
        RECT 1686.530 1870.290 1687.710 1871.470 ;
        RECT 1684.930 1691.890 1686.110 1693.070 ;
        RECT 1686.530 1691.890 1687.710 1693.070 ;
        RECT 1684.930 1690.290 1686.110 1691.470 ;
        RECT 1686.530 1690.290 1687.710 1691.470 ;
        RECT 1684.930 1511.890 1686.110 1513.070 ;
        RECT 1686.530 1511.890 1687.710 1513.070 ;
        RECT 1684.930 1510.290 1686.110 1511.470 ;
        RECT 1686.530 1510.290 1687.710 1511.470 ;
        RECT 1684.930 1331.890 1686.110 1333.070 ;
        RECT 1686.530 1331.890 1687.710 1333.070 ;
        RECT 1684.930 1330.290 1686.110 1331.470 ;
        RECT 1686.530 1330.290 1687.710 1331.470 ;
        RECT 1684.930 1151.890 1686.110 1153.070 ;
        RECT 1686.530 1151.890 1687.710 1153.070 ;
        RECT 1684.930 1150.290 1686.110 1151.470 ;
        RECT 1686.530 1150.290 1687.710 1151.470 ;
        RECT 1684.930 971.890 1686.110 973.070 ;
        RECT 1686.530 971.890 1687.710 973.070 ;
        RECT 1684.930 970.290 1686.110 971.470 ;
        RECT 1686.530 970.290 1687.710 971.470 ;
        RECT 1684.930 791.890 1686.110 793.070 ;
        RECT 1686.530 791.890 1687.710 793.070 ;
        RECT 1684.930 790.290 1686.110 791.470 ;
        RECT 1686.530 790.290 1687.710 791.470 ;
        RECT 1684.930 611.890 1686.110 613.070 ;
        RECT 1686.530 611.890 1687.710 613.070 ;
        RECT 1684.930 610.290 1686.110 611.470 ;
        RECT 1686.530 610.290 1687.710 611.470 ;
        RECT 1684.930 431.890 1686.110 433.070 ;
        RECT 1686.530 431.890 1687.710 433.070 ;
        RECT 1684.930 430.290 1686.110 431.470 ;
        RECT 1686.530 430.290 1687.710 431.470 ;
        RECT 1684.930 251.890 1686.110 253.070 ;
        RECT 1686.530 251.890 1687.710 253.070 ;
        RECT 1684.930 250.290 1686.110 251.470 ;
        RECT 1686.530 250.290 1687.710 251.470 ;
        RECT 1684.930 71.890 1686.110 73.070 ;
        RECT 1686.530 71.890 1687.710 73.070 ;
        RECT 1684.930 70.290 1686.110 71.470 ;
        RECT 1686.530 70.290 1687.710 71.470 ;
        RECT 1684.930 -31.710 1686.110 -30.530 ;
        RECT 1686.530 -31.710 1687.710 -30.530 ;
        RECT 1684.930 -33.310 1686.110 -32.130 ;
        RECT 1686.530 -33.310 1687.710 -32.130 ;
        RECT 1864.930 3551.810 1866.110 3552.990 ;
        RECT 1866.530 3551.810 1867.710 3552.990 ;
        RECT 1864.930 3550.210 1866.110 3551.390 ;
        RECT 1866.530 3550.210 1867.710 3551.390 ;
        RECT 1864.930 3491.890 1866.110 3493.070 ;
        RECT 1866.530 3491.890 1867.710 3493.070 ;
        RECT 1864.930 3490.290 1866.110 3491.470 ;
        RECT 1866.530 3490.290 1867.710 3491.470 ;
        RECT 1864.930 3311.890 1866.110 3313.070 ;
        RECT 1866.530 3311.890 1867.710 3313.070 ;
        RECT 1864.930 3310.290 1866.110 3311.470 ;
        RECT 1866.530 3310.290 1867.710 3311.470 ;
        RECT 1864.930 3131.890 1866.110 3133.070 ;
        RECT 1866.530 3131.890 1867.710 3133.070 ;
        RECT 1864.930 3130.290 1866.110 3131.470 ;
        RECT 1866.530 3130.290 1867.710 3131.470 ;
        RECT 1864.930 2951.890 1866.110 2953.070 ;
        RECT 1866.530 2951.890 1867.710 2953.070 ;
        RECT 1864.930 2950.290 1866.110 2951.470 ;
        RECT 1866.530 2950.290 1867.710 2951.470 ;
        RECT 1864.930 2771.890 1866.110 2773.070 ;
        RECT 1866.530 2771.890 1867.710 2773.070 ;
        RECT 1864.930 2770.290 1866.110 2771.470 ;
        RECT 1866.530 2770.290 1867.710 2771.470 ;
        RECT 1864.930 2591.890 1866.110 2593.070 ;
        RECT 1866.530 2591.890 1867.710 2593.070 ;
        RECT 1864.930 2590.290 1866.110 2591.470 ;
        RECT 1866.530 2590.290 1867.710 2591.470 ;
        RECT 1864.930 2411.890 1866.110 2413.070 ;
        RECT 1866.530 2411.890 1867.710 2413.070 ;
        RECT 1864.930 2410.290 1866.110 2411.470 ;
        RECT 1866.530 2410.290 1867.710 2411.470 ;
        RECT 1864.930 2231.890 1866.110 2233.070 ;
        RECT 1866.530 2231.890 1867.710 2233.070 ;
        RECT 1864.930 2230.290 1866.110 2231.470 ;
        RECT 1866.530 2230.290 1867.710 2231.470 ;
        RECT 1864.930 2051.890 1866.110 2053.070 ;
        RECT 1866.530 2051.890 1867.710 2053.070 ;
        RECT 1864.930 2050.290 1866.110 2051.470 ;
        RECT 1866.530 2050.290 1867.710 2051.470 ;
        RECT 1864.930 1871.890 1866.110 1873.070 ;
        RECT 1866.530 1871.890 1867.710 1873.070 ;
        RECT 1864.930 1870.290 1866.110 1871.470 ;
        RECT 1866.530 1870.290 1867.710 1871.470 ;
        RECT 1864.930 1691.890 1866.110 1693.070 ;
        RECT 1866.530 1691.890 1867.710 1693.070 ;
        RECT 1864.930 1690.290 1866.110 1691.470 ;
        RECT 1866.530 1690.290 1867.710 1691.470 ;
        RECT 1864.930 1511.890 1866.110 1513.070 ;
        RECT 1866.530 1511.890 1867.710 1513.070 ;
        RECT 1864.930 1510.290 1866.110 1511.470 ;
        RECT 1866.530 1510.290 1867.710 1511.470 ;
        RECT 1864.930 1331.890 1866.110 1333.070 ;
        RECT 1866.530 1331.890 1867.710 1333.070 ;
        RECT 1864.930 1330.290 1866.110 1331.470 ;
        RECT 1866.530 1330.290 1867.710 1331.470 ;
        RECT 1864.930 1151.890 1866.110 1153.070 ;
        RECT 1866.530 1151.890 1867.710 1153.070 ;
        RECT 1864.930 1150.290 1866.110 1151.470 ;
        RECT 1866.530 1150.290 1867.710 1151.470 ;
        RECT 1864.930 971.890 1866.110 973.070 ;
        RECT 1866.530 971.890 1867.710 973.070 ;
        RECT 1864.930 970.290 1866.110 971.470 ;
        RECT 1866.530 970.290 1867.710 971.470 ;
        RECT 1864.930 791.890 1866.110 793.070 ;
        RECT 1866.530 791.890 1867.710 793.070 ;
        RECT 1864.930 790.290 1866.110 791.470 ;
        RECT 1866.530 790.290 1867.710 791.470 ;
        RECT 1864.930 611.890 1866.110 613.070 ;
        RECT 1866.530 611.890 1867.710 613.070 ;
        RECT 1864.930 610.290 1866.110 611.470 ;
        RECT 1866.530 610.290 1867.710 611.470 ;
        RECT 1864.930 431.890 1866.110 433.070 ;
        RECT 1866.530 431.890 1867.710 433.070 ;
        RECT 1864.930 430.290 1866.110 431.470 ;
        RECT 1866.530 430.290 1867.710 431.470 ;
        RECT 1864.930 251.890 1866.110 253.070 ;
        RECT 1866.530 251.890 1867.710 253.070 ;
        RECT 1864.930 250.290 1866.110 251.470 ;
        RECT 1866.530 250.290 1867.710 251.470 ;
        RECT 1864.930 71.890 1866.110 73.070 ;
        RECT 1866.530 71.890 1867.710 73.070 ;
        RECT 1864.930 70.290 1866.110 71.470 ;
        RECT 1866.530 70.290 1867.710 71.470 ;
        RECT 1864.930 -31.710 1866.110 -30.530 ;
        RECT 1866.530 -31.710 1867.710 -30.530 ;
        RECT 1864.930 -33.310 1866.110 -32.130 ;
        RECT 1866.530 -33.310 1867.710 -32.130 ;
        RECT 2044.930 3551.810 2046.110 3552.990 ;
        RECT 2046.530 3551.810 2047.710 3552.990 ;
        RECT 2044.930 3550.210 2046.110 3551.390 ;
        RECT 2046.530 3550.210 2047.710 3551.390 ;
        RECT 2044.930 3491.890 2046.110 3493.070 ;
        RECT 2046.530 3491.890 2047.710 3493.070 ;
        RECT 2044.930 3490.290 2046.110 3491.470 ;
        RECT 2046.530 3490.290 2047.710 3491.470 ;
        RECT 2044.930 3311.890 2046.110 3313.070 ;
        RECT 2046.530 3311.890 2047.710 3313.070 ;
        RECT 2044.930 3310.290 2046.110 3311.470 ;
        RECT 2046.530 3310.290 2047.710 3311.470 ;
        RECT 2044.930 3131.890 2046.110 3133.070 ;
        RECT 2046.530 3131.890 2047.710 3133.070 ;
        RECT 2044.930 3130.290 2046.110 3131.470 ;
        RECT 2046.530 3130.290 2047.710 3131.470 ;
        RECT 2044.930 2951.890 2046.110 2953.070 ;
        RECT 2046.530 2951.890 2047.710 2953.070 ;
        RECT 2044.930 2950.290 2046.110 2951.470 ;
        RECT 2046.530 2950.290 2047.710 2951.470 ;
        RECT 2044.930 2771.890 2046.110 2773.070 ;
        RECT 2046.530 2771.890 2047.710 2773.070 ;
        RECT 2044.930 2770.290 2046.110 2771.470 ;
        RECT 2046.530 2770.290 2047.710 2771.470 ;
        RECT 2044.930 2591.890 2046.110 2593.070 ;
        RECT 2046.530 2591.890 2047.710 2593.070 ;
        RECT 2044.930 2590.290 2046.110 2591.470 ;
        RECT 2046.530 2590.290 2047.710 2591.470 ;
        RECT 2044.930 2411.890 2046.110 2413.070 ;
        RECT 2046.530 2411.890 2047.710 2413.070 ;
        RECT 2044.930 2410.290 2046.110 2411.470 ;
        RECT 2046.530 2410.290 2047.710 2411.470 ;
        RECT 2044.930 2231.890 2046.110 2233.070 ;
        RECT 2046.530 2231.890 2047.710 2233.070 ;
        RECT 2044.930 2230.290 2046.110 2231.470 ;
        RECT 2046.530 2230.290 2047.710 2231.470 ;
        RECT 2044.930 2051.890 2046.110 2053.070 ;
        RECT 2046.530 2051.890 2047.710 2053.070 ;
        RECT 2044.930 2050.290 2046.110 2051.470 ;
        RECT 2046.530 2050.290 2047.710 2051.470 ;
        RECT 2044.930 1871.890 2046.110 1873.070 ;
        RECT 2046.530 1871.890 2047.710 1873.070 ;
        RECT 2044.930 1870.290 2046.110 1871.470 ;
        RECT 2046.530 1870.290 2047.710 1871.470 ;
        RECT 2044.930 1691.890 2046.110 1693.070 ;
        RECT 2046.530 1691.890 2047.710 1693.070 ;
        RECT 2044.930 1690.290 2046.110 1691.470 ;
        RECT 2046.530 1690.290 2047.710 1691.470 ;
        RECT 2044.930 1511.890 2046.110 1513.070 ;
        RECT 2046.530 1511.890 2047.710 1513.070 ;
        RECT 2044.930 1510.290 2046.110 1511.470 ;
        RECT 2046.530 1510.290 2047.710 1511.470 ;
        RECT 2044.930 1331.890 2046.110 1333.070 ;
        RECT 2046.530 1331.890 2047.710 1333.070 ;
        RECT 2044.930 1330.290 2046.110 1331.470 ;
        RECT 2046.530 1330.290 2047.710 1331.470 ;
        RECT 2044.930 1151.890 2046.110 1153.070 ;
        RECT 2046.530 1151.890 2047.710 1153.070 ;
        RECT 2044.930 1150.290 2046.110 1151.470 ;
        RECT 2046.530 1150.290 2047.710 1151.470 ;
        RECT 2044.930 971.890 2046.110 973.070 ;
        RECT 2046.530 971.890 2047.710 973.070 ;
        RECT 2044.930 970.290 2046.110 971.470 ;
        RECT 2046.530 970.290 2047.710 971.470 ;
        RECT 2044.930 791.890 2046.110 793.070 ;
        RECT 2046.530 791.890 2047.710 793.070 ;
        RECT 2044.930 790.290 2046.110 791.470 ;
        RECT 2046.530 790.290 2047.710 791.470 ;
        RECT 2044.930 611.890 2046.110 613.070 ;
        RECT 2046.530 611.890 2047.710 613.070 ;
        RECT 2044.930 610.290 2046.110 611.470 ;
        RECT 2046.530 610.290 2047.710 611.470 ;
        RECT 2044.930 431.890 2046.110 433.070 ;
        RECT 2046.530 431.890 2047.710 433.070 ;
        RECT 2044.930 430.290 2046.110 431.470 ;
        RECT 2046.530 430.290 2047.710 431.470 ;
        RECT 2044.930 251.890 2046.110 253.070 ;
        RECT 2046.530 251.890 2047.710 253.070 ;
        RECT 2044.930 250.290 2046.110 251.470 ;
        RECT 2046.530 250.290 2047.710 251.470 ;
        RECT 2044.930 71.890 2046.110 73.070 ;
        RECT 2046.530 71.890 2047.710 73.070 ;
        RECT 2044.930 70.290 2046.110 71.470 ;
        RECT 2046.530 70.290 2047.710 71.470 ;
        RECT 2044.930 -31.710 2046.110 -30.530 ;
        RECT 2046.530 -31.710 2047.710 -30.530 ;
        RECT 2044.930 -33.310 2046.110 -32.130 ;
        RECT 2046.530 -33.310 2047.710 -32.130 ;
        RECT 2224.930 3551.810 2226.110 3552.990 ;
        RECT 2226.530 3551.810 2227.710 3552.990 ;
        RECT 2224.930 3550.210 2226.110 3551.390 ;
        RECT 2226.530 3550.210 2227.710 3551.390 ;
        RECT 2224.930 3491.890 2226.110 3493.070 ;
        RECT 2226.530 3491.890 2227.710 3493.070 ;
        RECT 2224.930 3490.290 2226.110 3491.470 ;
        RECT 2226.530 3490.290 2227.710 3491.470 ;
        RECT 2224.930 3311.890 2226.110 3313.070 ;
        RECT 2226.530 3311.890 2227.710 3313.070 ;
        RECT 2224.930 3310.290 2226.110 3311.470 ;
        RECT 2226.530 3310.290 2227.710 3311.470 ;
        RECT 2224.930 3131.890 2226.110 3133.070 ;
        RECT 2226.530 3131.890 2227.710 3133.070 ;
        RECT 2224.930 3130.290 2226.110 3131.470 ;
        RECT 2226.530 3130.290 2227.710 3131.470 ;
        RECT 2224.930 2951.890 2226.110 2953.070 ;
        RECT 2226.530 2951.890 2227.710 2953.070 ;
        RECT 2224.930 2950.290 2226.110 2951.470 ;
        RECT 2226.530 2950.290 2227.710 2951.470 ;
        RECT 2224.930 2771.890 2226.110 2773.070 ;
        RECT 2226.530 2771.890 2227.710 2773.070 ;
        RECT 2224.930 2770.290 2226.110 2771.470 ;
        RECT 2226.530 2770.290 2227.710 2771.470 ;
        RECT 2224.930 2591.890 2226.110 2593.070 ;
        RECT 2226.530 2591.890 2227.710 2593.070 ;
        RECT 2224.930 2590.290 2226.110 2591.470 ;
        RECT 2226.530 2590.290 2227.710 2591.470 ;
        RECT 2224.930 2411.890 2226.110 2413.070 ;
        RECT 2226.530 2411.890 2227.710 2413.070 ;
        RECT 2224.930 2410.290 2226.110 2411.470 ;
        RECT 2226.530 2410.290 2227.710 2411.470 ;
        RECT 2224.930 2231.890 2226.110 2233.070 ;
        RECT 2226.530 2231.890 2227.710 2233.070 ;
        RECT 2224.930 2230.290 2226.110 2231.470 ;
        RECT 2226.530 2230.290 2227.710 2231.470 ;
        RECT 2224.930 2051.890 2226.110 2053.070 ;
        RECT 2226.530 2051.890 2227.710 2053.070 ;
        RECT 2224.930 2050.290 2226.110 2051.470 ;
        RECT 2226.530 2050.290 2227.710 2051.470 ;
        RECT 2224.930 1871.890 2226.110 1873.070 ;
        RECT 2226.530 1871.890 2227.710 1873.070 ;
        RECT 2224.930 1870.290 2226.110 1871.470 ;
        RECT 2226.530 1870.290 2227.710 1871.470 ;
        RECT 2224.930 1691.890 2226.110 1693.070 ;
        RECT 2226.530 1691.890 2227.710 1693.070 ;
        RECT 2224.930 1690.290 2226.110 1691.470 ;
        RECT 2226.530 1690.290 2227.710 1691.470 ;
        RECT 2224.930 1511.890 2226.110 1513.070 ;
        RECT 2226.530 1511.890 2227.710 1513.070 ;
        RECT 2224.930 1510.290 2226.110 1511.470 ;
        RECT 2226.530 1510.290 2227.710 1511.470 ;
        RECT 2224.930 1331.890 2226.110 1333.070 ;
        RECT 2226.530 1331.890 2227.710 1333.070 ;
        RECT 2224.930 1330.290 2226.110 1331.470 ;
        RECT 2226.530 1330.290 2227.710 1331.470 ;
        RECT 2224.930 1151.890 2226.110 1153.070 ;
        RECT 2226.530 1151.890 2227.710 1153.070 ;
        RECT 2224.930 1150.290 2226.110 1151.470 ;
        RECT 2226.530 1150.290 2227.710 1151.470 ;
        RECT 2224.930 971.890 2226.110 973.070 ;
        RECT 2226.530 971.890 2227.710 973.070 ;
        RECT 2224.930 970.290 2226.110 971.470 ;
        RECT 2226.530 970.290 2227.710 971.470 ;
        RECT 2224.930 791.890 2226.110 793.070 ;
        RECT 2226.530 791.890 2227.710 793.070 ;
        RECT 2224.930 790.290 2226.110 791.470 ;
        RECT 2226.530 790.290 2227.710 791.470 ;
        RECT 2224.930 611.890 2226.110 613.070 ;
        RECT 2226.530 611.890 2227.710 613.070 ;
        RECT 2224.930 610.290 2226.110 611.470 ;
        RECT 2226.530 610.290 2227.710 611.470 ;
        RECT 2224.930 431.890 2226.110 433.070 ;
        RECT 2226.530 431.890 2227.710 433.070 ;
        RECT 2224.930 430.290 2226.110 431.470 ;
        RECT 2226.530 430.290 2227.710 431.470 ;
        RECT 2224.930 251.890 2226.110 253.070 ;
        RECT 2226.530 251.890 2227.710 253.070 ;
        RECT 2224.930 250.290 2226.110 251.470 ;
        RECT 2226.530 250.290 2227.710 251.470 ;
        RECT 2224.930 71.890 2226.110 73.070 ;
        RECT 2226.530 71.890 2227.710 73.070 ;
        RECT 2224.930 70.290 2226.110 71.470 ;
        RECT 2226.530 70.290 2227.710 71.470 ;
        RECT 2224.930 -31.710 2226.110 -30.530 ;
        RECT 2226.530 -31.710 2227.710 -30.530 ;
        RECT 2224.930 -33.310 2226.110 -32.130 ;
        RECT 2226.530 -33.310 2227.710 -32.130 ;
        RECT 2404.930 3551.810 2406.110 3552.990 ;
        RECT 2406.530 3551.810 2407.710 3552.990 ;
        RECT 2404.930 3550.210 2406.110 3551.390 ;
        RECT 2406.530 3550.210 2407.710 3551.390 ;
        RECT 2404.930 3491.890 2406.110 3493.070 ;
        RECT 2406.530 3491.890 2407.710 3493.070 ;
        RECT 2404.930 3490.290 2406.110 3491.470 ;
        RECT 2406.530 3490.290 2407.710 3491.470 ;
        RECT 2404.930 3311.890 2406.110 3313.070 ;
        RECT 2406.530 3311.890 2407.710 3313.070 ;
        RECT 2404.930 3310.290 2406.110 3311.470 ;
        RECT 2406.530 3310.290 2407.710 3311.470 ;
        RECT 2404.930 3131.890 2406.110 3133.070 ;
        RECT 2406.530 3131.890 2407.710 3133.070 ;
        RECT 2404.930 3130.290 2406.110 3131.470 ;
        RECT 2406.530 3130.290 2407.710 3131.470 ;
        RECT 2404.930 2951.890 2406.110 2953.070 ;
        RECT 2406.530 2951.890 2407.710 2953.070 ;
        RECT 2404.930 2950.290 2406.110 2951.470 ;
        RECT 2406.530 2950.290 2407.710 2951.470 ;
        RECT 2404.930 2771.890 2406.110 2773.070 ;
        RECT 2406.530 2771.890 2407.710 2773.070 ;
        RECT 2404.930 2770.290 2406.110 2771.470 ;
        RECT 2406.530 2770.290 2407.710 2771.470 ;
        RECT 2404.930 2591.890 2406.110 2593.070 ;
        RECT 2406.530 2591.890 2407.710 2593.070 ;
        RECT 2404.930 2590.290 2406.110 2591.470 ;
        RECT 2406.530 2590.290 2407.710 2591.470 ;
        RECT 2404.930 2411.890 2406.110 2413.070 ;
        RECT 2406.530 2411.890 2407.710 2413.070 ;
        RECT 2404.930 2410.290 2406.110 2411.470 ;
        RECT 2406.530 2410.290 2407.710 2411.470 ;
        RECT 2404.930 2231.890 2406.110 2233.070 ;
        RECT 2406.530 2231.890 2407.710 2233.070 ;
        RECT 2404.930 2230.290 2406.110 2231.470 ;
        RECT 2406.530 2230.290 2407.710 2231.470 ;
        RECT 2404.930 2051.890 2406.110 2053.070 ;
        RECT 2406.530 2051.890 2407.710 2053.070 ;
        RECT 2404.930 2050.290 2406.110 2051.470 ;
        RECT 2406.530 2050.290 2407.710 2051.470 ;
        RECT 2404.930 1871.890 2406.110 1873.070 ;
        RECT 2406.530 1871.890 2407.710 1873.070 ;
        RECT 2404.930 1870.290 2406.110 1871.470 ;
        RECT 2406.530 1870.290 2407.710 1871.470 ;
        RECT 2404.930 1691.890 2406.110 1693.070 ;
        RECT 2406.530 1691.890 2407.710 1693.070 ;
        RECT 2404.930 1690.290 2406.110 1691.470 ;
        RECT 2406.530 1690.290 2407.710 1691.470 ;
        RECT 2404.930 1511.890 2406.110 1513.070 ;
        RECT 2406.530 1511.890 2407.710 1513.070 ;
        RECT 2404.930 1510.290 2406.110 1511.470 ;
        RECT 2406.530 1510.290 2407.710 1511.470 ;
        RECT 2404.930 1331.890 2406.110 1333.070 ;
        RECT 2406.530 1331.890 2407.710 1333.070 ;
        RECT 2404.930 1330.290 2406.110 1331.470 ;
        RECT 2406.530 1330.290 2407.710 1331.470 ;
        RECT 2404.930 1151.890 2406.110 1153.070 ;
        RECT 2406.530 1151.890 2407.710 1153.070 ;
        RECT 2404.930 1150.290 2406.110 1151.470 ;
        RECT 2406.530 1150.290 2407.710 1151.470 ;
        RECT 2404.930 971.890 2406.110 973.070 ;
        RECT 2406.530 971.890 2407.710 973.070 ;
        RECT 2404.930 970.290 2406.110 971.470 ;
        RECT 2406.530 970.290 2407.710 971.470 ;
        RECT 2404.930 791.890 2406.110 793.070 ;
        RECT 2406.530 791.890 2407.710 793.070 ;
        RECT 2404.930 790.290 2406.110 791.470 ;
        RECT 2406.530 790.290 2407.710 791.470 ;
        RECT 2404.930 611.890 2406.110 613.070 ;
        RECT 2406.530 611.890 2407.710 613.070 ;
        RECT 2404.930 610.290 2406.110 611.470 ;
        RECT 2406.530 610.290 2407.710 611.470 ;
        RECT 2404.930 431.890 2406.110 433.070 ;
        RECT 2406.530 431.890 2407.710 433.070 ;
        RECT 2404.930 430.290 2406.110 431.470 ;
        RECT 2406.530 430.290 2407.710 431.470 ;
        RECT 2404.930 251.890 2406.110 253.070 ;
        RECT 2406.530 251.890 2407.710 253.070 ;
        RECT 2404.930 250.290 2406.110 251.470 ;
        RECT 2406.530 250.290 2407.710 251.470 ;
        RECT 2404.930 71.890 2406.110 73.070 ;
        RECT 2406.530 71.890 2407.710 73.070 ;
        RECT 2404.930 70.290 2406.110 71.470 ;
        RECT 2406.530 70.290 2407.710 71.470 ;
        RECT 2404.930 -31.710 2406.110 -30.530 ;
        RECT 2406.530 -31.710 2407.710 -30.530 ;
        RECT 2404.930 -33.310 2406.110 -32.130 ;
        RECT 2406.530 -33.310 2407.710 -32.130 ;
        RECT 2584.930 3551.810 2586.110 3552.990 ;
        RECT 2586.530 3551.810 2587.710 3552.990 ;
        RECT 2584.930 3550.210 2586.110 3551.390 ;
        RECT 2586.530 3550.210 2587.710 3551.390 ;
        RECT 2584.930 3491.890 2586.110 3493.070 ;
        RECT 2586.530 3491.890 2587.710 3493.070 ;
        RECT 2584.930 3490.290 2586.110 3491.470 ;
        RECT 2586.530 3490.290 2587.710 3491.470 ;
        RECT 2584.930 3311.890 2586.110 3313.070 ;
        RECT 2586.530 3311.890 2587.710 3313.070 ;
        RECT 2584.930 3310.290 2586.110 3311.470 ;
        RECT 2586.530 3310.290 2587.710 3311.470 ;
        RECT 2584.930 3131.890 2586.110 3133.070 ;
        RECT 2586.530 3131.890 2587.710 3133.070 ;
        RECT 2584.930 3130.290 2586.110 3131.470 ;
        RECT 2586.530 3130.290 2587.710 3131.470 ;
        RECT 2584.930 2951.890 2586.110 2953.070 ;
        RECT 2586.530 2951.890 2587.710 2953.070 ;
        RECT 2584.930 2950.290 2586.110 2951.470 ;
        RECT 2586.530 2950.290 2587.710 2951.470 ;
        RECT 2584.930 2771.890 2586.110 2773.070 ;
        RECT 2586.530 2771.890 2587.710 2773.070 ;
        RECT 2584.930 2770.290 2586.110 2771.470 ;
        RECT 2586.530 2770.290 2587.710 2771.470 ;
        RECT 2584.930 2591.890 2586.110 2593.070 ;
        RECT 2586.530 2591.890 2587.710 2593.070 ;
        RECT 2584.930 2590.290 2586.110 2591.470 ;
        RECT 2586.530 2590.290 2587.710 2591.470 ;
        RECT 2584.930 2411.890 2586.110 2413.070 ;
        RECT 2586.530 2411.890 2587.710 2413.070 ;
        RECT 2584.930 2410.290 2586.110 2411.470 ;
        RECT 2586.530 2410.290 2587.710 2411.470 ;
        RECT 2584.930 2231.890 2586.110 2233.070 ;
        RECT 2586.530 2231.890 2587.710 2233.070 ;
        RECT 2584.930 2230.290 2586.110 2231.470 ;
        RECT 2586.530 2230.290 2587.710 2231.470 ;
        RECT 2584.930 2051.890 2586.110 2053.070 ;
        RECT 2586.530 2051.890 2587.710 2053.070 ;
        RECT 2584.930 2050.290 2586.110 2051.470 ;
        RECT 2586.530 2050.290 2587.710 2051.470 ;
        RECT 2584.930 1871.890 2586.110 1873.070 ;
        RECT 2586.530 1871.890 2587.710 1873.070 ;
        RECT 2584.930 1870.290 2586.110 1871.470 ;
        RECT 2586.530 1870.290 2587.710 1871.470 ;
        RECT 2584.930 1691.890 2586.110 1693.070 ;
        RECT 2586.530 1691.890 2587.710 1693.070 ;
        RECT 2584.930 1690.290 2586.110 1691.470 ;
        RECT 2586.530 1690.290 2587.710 1691.470 ;
        RECT 2584.930 1511.890 2586.110 1513.070 ;
        RECT 2586.530 1511.890 2587.710 1513.070 ;
        RECT 2584.930 1510.290 2586.110 1511.470 ;
        RECT 2586.530 1510.290 2587.710 1511.470 ;
        RECT 2584.930 1331.890 2586.110 1333.070 ;
        RECT 2586.530 1331.890 2587.710 1333.070 ;
        RECT 2584.930 1330.290 2586.110 1331.470 ;
        RECT 2586.530 1330.290 2587.710 1331.470 ;
        RECT 2584.930 1151.890 2586.110 1153.070 ;
        RECT 2586.530 1151.890 2587.710 1153.070 ;
        RECT 2584.930 1150.290 2586.110 1151.470 ;
        RECT 2586.530 1150.290 2587.710 1151.470 ;
        RECT 2584.930 971.890 2586.110 973.070 ;
        RECT 2586.530 971.890 2587.710 973.070 ;
        RECT 2584.930 970.290 2586.110 971.470 ;
        RECT 2586.530 970.290 2587.710 971.470 ;
        RECT 2584.930 791.890 2586.110 793.070 ;
        RECT 2586.530 791.890 2587.710 793.070 ;
        RECT 2584.930 790.290 2586.110 791.470 ;
        RECT 2586.530 790.290 2587.710 791.470 ;
        RECT 2584.930 611.890 2586.110 613.070 ;
        RECT 2586.530 611.890 2587.710 613.070 ;
        RECT 2584.930 610.290 2586.110 611.470 ;
        RECT 2586.530 610.290 2587.710 611.470 ;
        RECT 2584.930 431.890 2586.110 433.070 ;
        RECT 2586.530 431.890 2587.710 433.070 ;
        RECT 2584.930 430.290 2586.110 431.470 ;
        RECT 2586.530 430.290 2587.710 431.470 ;
        RECT 2584.930 251.890 2586.110 253.070 ;
        RECT 2586.530 251.890 2587.710 253.070 ;
        RECT 2584.930 250.290 2586.110 251.470 ;
        RECT 2586.530 250.290 2587.710 251.470 ;
        RECT 2584.930 71.890 2586.110 73.070 ;
        RECT 2586.530 71.890 2587.710 73.070 ;
        RECT 2584.930 70.290 2586.110 71.470 ;
        RECT 2586.530 70.290 2587.710 71.470 ;
        RECT 2584.930 -31.710 2586.110 -30.530 ;
        RECT 2586.530 -31.710 2587.710 -30.530 ;
        RECT 2584.930 -33.310 2586.110 -32.130 ;
        RECT 2586.530 -33.310 2587.710 -32.130 ;
        RECT 2764.930 3551.810 2766.110 3552.990 ;
        RECT 2766.530 3551.810 2767.710 3552.990 ;
        RECT 2764.930 3550.210 2766.110 3551.390 ;
        RECT 2766.530 3550.210 2767.710 3551.390 ;
        RECT 2764.930 3491.890 2766.110 3493.070 ;
        RECT 2766.530 3491.890 2767.710 3493.070 ;
        RECT 2764.930 3490.290 2766.110 3491.470 ;
        RECT 2766.530 3490.290 2767.710 3491.470 ;
        RECT 2764.930 3311.890 2766.110 3313.070 ;
        RECT 2766.530 3311.890 2767.710 3313.070 ;
        RECT 2764.930 3310.290 2766.110 3311.470 ;
        RECT 2766.530 3310.290 2767.710 3311.470 ;
        RECT 2764.930 3131.890 2766.110 3133.070 ;
        RECT 2766.530 3131.890 2767.710 3133.070 ;
        RECT 2764.930 3130.290 2766.110 3131.470 ;
        RECT 2766.530 3130.290 2767.710 3131.470 ;
        RECT 2764.930 2951.890 2766.110 2953.070 ;
        RECT 2766.530 2951.890 2767.710 2953.070 ;
        RECT 2764.930 2950.290 2766.110 2951.470 ;
        RECT 2766.530 2950.290 2767.710 2951.470 ;
        RECT 2764.930 2771.890 2766.110 2773.070 ;
        RECT 2766.530 2771.890 2767.710 2773.070 ;
        RECT 2764.930 2770.290 2766.110 2771.470 ;
        RECT 2766.530 2770.290 2767.710 2771.470 ;
        RECT 2764.930 2591.890 2766.110 2593.070 ;
        RECT 2766.530 2591.890 2767.710 2593.070 ;
        RECT 2764.930 2590.290 2766.110 2591.470 ;
        RECT 2766.530 2590.290 2767.710 2591.470 ;
        RECT 2764.930 2411.890 2766.110 2413.070 ;
        RECT 2766.530 2411.890 2767.710 2413.070 ;
        RECT 2764.930 2410.290 2766.110 2411.470 ;
        RECT 2766.530 2410.290 2767.710 2411.470 ;
        RECT 2764.930 2231.890 2766.110 2233.070 ;
        RECT 2766.530 2231.890 2767.710 2233.070 ;
        RECT 2764.930 2230.290 2766.110 2231.470 ;
        RECT 2766.530 2230.290 2767.710 2231.470 ;
        RECT 2764.930 2051.890 2766.110 2053.070 ;
        RECT 2766.530 2051.890 2767.710 2053.070 ;
        RECT 2764.930 2050.290 2766.110 2051.470 ;
        RECT 2766.530 2050.290 2767.710 2051.470 ;
        RECT 2764.930 1871.890 2766.110 1873.070 ;
        RECT 2766.530 1871.890 2767.710 1873.070 ;
        RECT 2764.930 1870.290 2766.110 1871.470 ;
        RECT 2766.530 1870.290 2767.710 1871.470 ;
        RECT 2764.930 1691.890 2766.110 1693.070 ;
        RECT 2766.530 1691.890 2767.710 1693.070 ;
        RECT 2764.930 1690.290 2766.110 1691.470 ;
        RECT 2766.530 1690.290 2767.710 1691.470 ;
        RECT 2764.930 1511.890 2766.110 1513.070 ;
        RECT 2766.530 1511.890 2767.710 1513.070 ;
        RECT 2764.930 1510.290 2766.110 1511.470 ;
        RECT 2766.530 1510.290 2767.710 1511.470 ;
        RECT 2764.930 1331.890 2766.110 1333.070 ;
        RECT 2766.530 1331.890 2767.710 1333.070 ;
        RECT 2764.930 1330.290 2766.110 1331.470 ;
        RECT 2766.530 1330.290 2767.710 1331.470 ;
        RECT 2764.930 1151.890 2766.110 1153.070 ;
        RECT 2766.530 1151.890 2767.710 1153.070 ;
        RECT 2764.930 1150.290 2766.110 1151.470 ;
        RECT 2766.530 1150.290 2767.710 1151.470 ;
        RECT 2764.930 971.890 2766.110 973.070 ;
        RECT 2766.530 971.890 2767.710 973.070 ;
        RECT 2764.930 970.290 2766.110 971.470 ;
        RECT 2766.530 970.290 2767.710 971.470 ;
        RECT 2764.930 791.890 2766.110 793.070 ;
        RECT 2766.530 791.890 2767.710 793.070 ;
        RECT 2764.930 790.290 2766.110 791.470 ;
        RECT 2766.530 790.290 2767.710 791.470 ;
        RECT 2764.930 611.890 2766.110 613.070 ;
        RECT 2766.530 611.890 2767.710 613.070 ;
        RECT 2764.930 610.290 2766.110 611.470 ;
        RECT 2766.530 610.290 2767.710 611.470 ;
        RECT 2764.930 431.890 2766.110 433.070 ;
        RECT 2766.530 431.890 2767.710 433.070 ;
        RECT 2764.930 430.290 2766.110 431.470 ;
        RECT 2766.530 430.290 2767.710 431.470 ;
        RECT 2764.930 251.890 2766.110 253.070 ;
        RECT 2766.530 251.890 2767.710 253.070 ;
        RECT 2764.930 250.290 2766.110 251.470 ;
        RECT 2766.530 250.290 2767.710 251.470 ;
        RECT 2764.930 71.890 2766.110 73.070 ;
        RECT 2766.530 71.890 2767.710 73.070 ;
        RECT 2764.930 70.290 2766.110 71.470 ;
        RECT 2766.530 70.290 2767.710 71.470 ;
        RECT 2764.930 -31.710 2766.110 -30.530 ;
        RECT 2766.530 -31.710 2767.710 -30.530 ;
        RECT 2764.930 -33.310 2766.110 -32.130 ;
        RECT 2766.530 -33.310 2767.710 -32.130 ;
        RECT 2955.510 3551.810 2956.690 3552.990 ;
        RECT 2957.110 3551.810 2958.290 3552.990 ;
        RECT 2955.510 3550.210 2956.690 3551.390 ;
        RECT 2957.110 3550.210 2958.290 3551.390 ;
        RECT 2955.510 3491.890 2956.690 3493.070 ;
        RECT 2957.110 3491.890 2958.290 3493.070 ;
        RECT 2955.510 3490.290 2956.690 3491.470 ;
        RECT 2957.110 3490.290 2958.290 3491.470 ;
        RECT 2955.510 3311.890 2956.690 3313.070 ;
        RECT 2957.110 3311.890 2958.290 3313.070 ;
        RECT 2955.510 3310.290 2956.690 3311.470 ;
        RECT 2957.110 3310.290 2958.290 3311.470 ;
        RECT 2955.510 3131.890 2956.690 3133.070 ;
        RECT 2957.110 3131.890 2958.290 3133.070 ;
        RECT 2955.510 3130.290 2956.690 3131.470 ;
        RECT 2957.110 3130.290 2958.290 3131.470 ;
        RECT 2955.510 2951.890 2956.690 2953.070 ;
        RECT 2957.110 2951.890 2958.290 2953.070 ;
        RECT 2955.510 2950.290 2956.690 2951.470 ;
        RECT 2957.110 2950.290 2958.290 2951.470 ;
        RECT 2955.510 2771.890 2956.690 2773.070 ;
        RECT 2957.110 2771.890 2958.290 2773.070 ;
        RECT 2955.510 2770.290 2956.690 2771.470 ;
        RECT 2957.110 2770.290 2958.290 2771.470 ;
        RECT 2955.510 2591.890 2956.690 2593.070 ;
        RECT 2957.110 2591.890 2958.290 2593.070 ;
        RECT 2955.510 2590.290 2956.690 2591.470 ;
        RECT 2957.110 2590.290 2958.290 2591.470 ;
        RECT 2955.510 2411.890 2956.690 2413.070 ;
        RECT 2957.110 2411.890 2958.290 2413.070 ;
        RECT 2955.510 2410.290 2956.690 2411.470 ;
        RECT 2957.110 2410.290 2958.290 2411.470 ;
        RECT 2955.510 2231.890 2956.690 2233.070 ;
        RECT 2957.110 2231.890 2958.290 2233.070 ;
        RECT 2955.510 2230.290 2956.690 2231.470 ;
        RECT 2957.110 2230.290 2958.290 2231.470 ;
        RECT 2955.510 2051.890 2956.690 2053.070 ;
        RECT 2957.110 2051.890 2958.290 2053.070 ;
        RECT 2955.510 2050.290 2956.690 2051.470 ;
        RECT 2957.110 2050.290 2958.290 2051.470 ;
        RECT 2955.510 1871.890 2956.690 1873.070 ;
        RECT 2957.110 1871.890 2958.290 1873.070 ;
        RECT 2955.510 1870.290 2956.690 1871.470 ;
        RECT 2957.110 1870.290 2958.290 1871.470 ;
        RECT 2955.510 1691.890 2956.690 1693.070 ;
        RECT 2957.110 1691.890 2958.290 1693.070 ;
        RECT 2955.510 1690.290 2956.690 1691.470 ;
        RECT 2957.110 1690.290 2958.290 1691.470 ;
        RECT 2955.510 1511.890 2956.690 1513.070 ;
        RECT 2957.110 1511.890 2958.290 1513.070 ;
        RECT 2955.510 1510.290 2956.690 1511.470 ;
        RECT 2957.110 1510.290 2958.290 1511.470 ;
        RECT 2955.510 1331.890 2956.690 1333.070 ;
        RECT 2957.110 1331.890 2958.290 1333.070 ;
        RECT 2955.510 1330.290 2956.690 1331.470 ;
        RECT 2957.110 1330.290 2958.290 1331.470 ;
        RECT 2955.510 1151.890 2956.690 1153.070 ;
        RECT 2957.110 1151.890 2958.290 1153.070 ;
        RECT 2955.510 1150.290 2956.690 1151.470 ;
        RECT 2957.110 1150.290 2958.290 1151.470 ;
        RECT 2955.510 971.890 2956.690 973.070 ;
        RECT 2957.110 971.890 2958.290 973.070 ;
        RECT 2955.510 970.290 2956.690 971.470 ;
        RECT 2957.110 970.290 2958.290 971.470 ;
        RECT 2955.510 791.890 2956.690 793.070 ;
        RECT 2957.110 791.890 2958.290 793.070 ;
        RECT 2955.510 790.290 2956.690 791.470 ;
        RECT 2957.110 790.290 2958.290 791.470 ;
        RECT 2955.510 611.890 2956.690 613.070 ;
        RECT 2957.110 611.890 2958.290 613.070 ;
        RECT 2955.510 610.290 2956.690 611.470 ;
        RECT 2957.110 610.290 2958.290 611.470 ;
        RECT 2955.510 431.890 2956.690 433.070 ;
        RECT 2957.110 431.890 2958.290 433.070 ;
        RECT 2955.510 430.290 2956.690 431.470 ;
        RECT 2957.110 430.290 2958.290 431.470 ;
        RECT 2955.510 251.890 2956.690 253.070 ;
        RECT 2957.110 251.890 2958.290 253.070 ;
        RECT 2955.510 250.290 2956.690 251.470 ;
        RECT 2957.110 250.290 2958.290 251.470 ;
        RECT 2955.510 71.890 2956.690 73.070 ;
        RECT 2957.110 71.890 2958.290 73.070 ;
        RECT 2955.510 70.290 2956.690 71.470 ;
        RECT 2957.110 70.290 2958.290 71.470 ;
        RECT 2955.510 -31.710 2956.690 -30.530 ;
        RECT 2957.110 -31.710 2958.290 -30.530 ;
        RECT 2955.510 -33.310 2956.690 -32.130 ;
        RECT 2957.110 -33.310 2958.290 -32.130 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
        RECT -43.630 970.130 2963.250 973.230 ;
        RECT -43.630 790.130 2963.250 793.230 ;
        RECT -43.630 610.130 2963.250 613.230 ;
        RECT -43.630 430.130 2963.250 433.230 ;
        RECT -43.630 250.130 2963.250 253.230 ;
        RECT -43.630 70.130 2963.250 73.230 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
        RECT 316.170 1010.000 319.270 3548.350 ;
        RECT 496.170 1010.000 499.270 3548.350 ;
        RECT 676.170 1010.000 679.270 3548.350 ;
        RECT 856.170 1010.000 859.270 3548.350 ;
        RECT 1036.170 1010.000 1039.270 3548.350 ;
        RECT 316.170 -28.670 319.270 390.000 ;
        RECT 496.170 -28.670 499.270 390.000 ;
        RECT 676.170 -28.670 679.270 390.000 ;
        RECT 856.170 -28.670 859.270 390.000 ;
        RECT 1036.170 -28.670 1039.270 390.000 ;
        RECT 1216.170 -28.670 1219.270 3548.350 ;
        RECT 1396.170 -28.670 1399.270 3548.350 ;
        RECT 1576.170 -28.670 1579.270 3548.350 ;
        RECT 1756.170 -28.670 1759.270 3548.350 ;
        RECT 1936.170 -28.670 1939.270 3548.350 ;
        RECT 2116.170 -28.670 2119.270 3548.350 ;
        RECT 2296.170 -28.670 2299.270 3548.350 ;
        RECT 2476.170 -28.670 2479.270 3548.350 ;
        RECT 2656.170 -28.670 2659.270 3548.350 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER via4 ;
        RECT -33.870 3547.010 -32.690 3548.190 ;
        RECT -32.270 3547.010 -31.090 3548.190 ;
        RECT -33.870 3545.410 -32.690 3546.590 ;
        RECT -32.270 3545.410 -31.090 3546.590 ;
        RECT -33.870 3383.290 -32.690 3384.470 ;
        RECT -32.270 3383.290 -31.090 3384.470 ;
        RECT -33.870 3381.690 -32.690 3382.870 ;
        RECT -32.270 3381.690 -31.090 3382.870 ;
        RECT -33.870 3203.290 -32.690 3204.470 ;
        RECT -32.270 3203.290 -31.090 3204.470 ;
        RECT -33.870 3201.690 -32.690 3202.870 ;
        RECT -32.270 3201.690 -31.090 3202.870 ;
        RECT -33.870 3023.290 -32.690 3024.470 ;
        RECT -32.270 3023.290 -31.090 3024.470 ;
        RECT -33.870 3021.690 -32.690 3022.870 ;
        RECT -32.270 3021.690 -31.090 3022.870 ;
        RECT -33.870 2843.290 -32.690 2844.470 ;
        RECT -32.270 2843.290 -31.090 2844.470 ;
        RECT -33.870 2841.690 -32.690 2842.870 ;
        RECT -32.270 2841.690 -31.090 2842.870 ;
        RECT -33.870 2663.290 -32.690 2664.470 ;
        RECT -32.270 2663.290 -31.090 2664.470 ;
        RECT -33.870 2661.690 -32.690 2662.870 ;
        RECT -32.270 2661.690 -31.090 2662.870 ;
        RECT -33.870 2483.290 -32.690 2484.470 ;
        RECT -32.270 2483.290 -31.090 2484.470 ;
        RECT -33.870 2481.690 -32.690 2482.870 ;
        RECT -32.270 2481.690 -31.090 2482.870 ;
        RECT -33.870 2303.290 -32.690 2304.470 ;
        RECT -32.270 2303.290 -31.090 2304.470 ;
        RECT -33.870 2301.690 -32.690 2302.870 ;
        RECT -32.270 2301.690 -31.090 2302.870 ;
        RECT -33.870 2123.290 -32.690 2124.470 ;
        RECT -32.270 2123.290 -31.090 2124.470 ;
        RECT -33.870 2121.690 -32.690 2122.870 ;
        RECT -32.270 2121.690 -31.090 2122.870 ;
        RECT -33.870 1943.290 -32.690 1944.470 ;
        RECT -32.270 1943.290 -31.090 1944.470 ;
        RECT -33.870 1941.690 -32.690 1942.870 ;
        RECT -32.270 1941.690 -31.090 1942.870 ;
        RECT -33.870 1763.290 -32.690 1764.470 ;
        RECT -32.270 1763.290 -31.090 1764.470 ;
        RECT -33.870 1761.690 -32.690 1762.870 ;
        RECT -32.270 1761.690 -31.090 1762.870 ;
        RECT -33.870 1583.290 -32.690 1584.470 ;
        RECT -32.270 1583.290 -31.090 1584.470 ;
        RECT -33.870 1581.690 -32.690 1582.870 ;
        RECT -32.270 1581.690 -31.090 1582.870 ;
        RECT -33.870 1403.290 -32.690 1404.470 ;
        RECT -32.270 1403.290 -31.090 1404.470 ;
        RECT -33.870 1401.690 -32.690 1402.870 ;
        RECT -32.270 1401.690 -31.090 1402.870 ;
        RECT -33.870 1223.290 -32.690 1224.470 ;
        RECT -32.270 1223.290 -31.090 1224.470 ;
        RECT -33.870 1221.690 -32.690 1222.870 ;
        RECT -32.270 1221.690 -31.090 1222.870 ;
        RECT -33.870 1043.290 -32.690 1044.470 ;
        RECT -32.270 1043.290 -31.090 1044.470 ;
        RECT -33.870 1041.690 -32.690 1042.870 ;
        RECT -32.270 1041.690 -31.090 1042.870 ;
        RECT -33.870 863.290 -32.690 864.470 ;
        RECT -32.270 863.290 -31.090 864.470 ;
        RECT -33.870 861.690 -32.690 862.870 ;
        RECT -32.270 861.690 -31.090 862.870 ;
        RECT -33.870 683.290 -32.690 684.470 ;
        RECT -32.270 683.290 -31.090 684.470 ;
        RECT -33.870 681.690 -32.690 682.870 ;
        RECT -32.270 681.690 -31.090 682.870 ;
        RECT -33.870 503.290 -32.690 504.470 ;
        RECT -32.270 503.290 -31.090 504.470 ;
        RECT -33.870 501.690 -32.690 502.870 ;
        RECT -32.270 501.690 -31.090 502.870 ;
        RECT -33.870 323.290 -32.690 324.470 ;
        RECT -32.270 323.290 -31.090 324.470 ;
        RECT -33.870 321.690 -32.690 322.870 ;
        RECT -32.270 321.690 -31.090 322.870 ;
        RECT -33.870 143.290 -32.690 144.470 ;
        RECT -32.270 143.290 -31.090 144.470 ;
        RECT -33.870 141.690 -32.690 142.870 ;
        RECT -32.270 141.690 -31.090 142.870 ;
        RECT -33.870 -26.910 -32.690 -25.730 ;
        RECT -32.270 -26.910 -31.090 -25.730 ;
        RECT -33.870 -28.510 -32.690 -27.330 ;
        RECT -32.270 -28.510 -31.090 -27.330 ;
        RECT 136.330 3547.010 137.510 3548.190 ;
        RECT 137.930 3547.010 139.110 3548.190 ;
        RECT 136.330 3545.410 137.510 3546.590 ;
        RECT 137.930 3545.410 139.110 3546.590 ;
        RECT 136.330 3383.290 137.510 3384.470 ;
        RECT 137.930 3383.290 139.110 3384.470 ;
        RECT 136.330 3381.690 137.510 3382.870 ;
        RECT 137.930 3381.690 139.110 3382.870 ;
        RECT 136.330 3203.290 137.510 3204.470 ;
        RECT 137.930 3203.290 139.110 3204.470 ;
        RECT 136.330 3201.690 137.510 3202.870 ;
        RECT 137.930 3201.690 139.110 3202.870 ;
        RECT 136.330 3023.290 137.510 3024.470 ;
        RECT 137.930 3023.290 139.110 3024.470 ;
        RECT 136.330 3021.690 137.510 3022.870 ;
        RECT 137.930 3021.690 139.110 3022.870 ;
        RECT 136.330 2843.290 137.510 2844.470 ;
        RECT 137.930 2843.290 139.110 2844.470 ;
        RECT 136.330 2841.690 137.510 2842.870 ;
        RECT 137.930 2841.690 139.110 2842.870 ;
        RECT 136.330 2663.290 137.510 2664.470 ;
        RECT 137.930 2663.290 139.110 2664.470 ;
        RECT 136.330 2661.690 137.510 2662.870 ;
        RECT 137.930 2661.690 139.110 2662.870 ;
        RECT 136.330 2483.290 137.510 2484.470 ;
        RECT 137.930 2483.290 139.110 2484.470 ;
        RECT 136.330 2481.690 137.510 2482.870 ;
        RECT 137.930 2481.690 139.110 2482.870 ;
        RECT 136.330 2303.290 137.510 2304.470 ;
        RECT 137.930 2303.290 139.110 2304.470 ;
        RECT 136.330 2301.690 137.510 2302.870 ;
        RECT 137.930 2301.690 139.110 2302.870 ;
        RECT 136.330 2123.290 137.510 2124.470 ;
        RECT 137.930 2123.290 139.110 2124.470 ;
        RECT 136.330 2121.690 137.510 2122.870 ;
        RECT 137.930 2121.690 139.110 2122.870 ;
        RECT 136.330 1943.290 137.510 1944.470 ;
        RECT 137.930 1943.290 139.110 1944.470 ;
        RECT 136.330 1941.690 137.510 1942.870 ;
        RECT 137.930 1941.690 139.110 1942.870 ;
        RECT 136.330 1763.290 137.510 1764.470 ;
        RECT 137.930 1763.290 139.110 1764.470 ;
        RECT 136.330 1761.690 137.510 1762.870 ;
        RECT 137.930 1761.690 139.110 1762.870 ;
        RECT 136.330 1583.290 137.510 1584.470 ;
        RECT 137.930 1583.290 139.110 1584.470 ;
        RECT 136.330 1581.690 137.510 1582.870 ;
        RECT 137.930 1581.690 139.110 1582.870 ;
        RECT 136.330 1403.290 137.510 1404.470 ;
        RECT 137.930 1403.290 139.110 1404.470 ;
        RECT 136.330 1401.690 137.510 1402.870 ;
        RECT 137.930 1401.690 139.110 1402.870 ;
        RECT 136.330 1223.290 137.510 1224.470 ;
        RECT 137.930 1223.290 139.110 1224.470 ;
        RECT 136.330 1221.690 137.510 1222.870 ;
        RECT 137.930 1221.690 139.110 1222.870 ;
        RECT 136.330 1043.290 137.510 1044.470 ;
        RECT 137.930 1043.290 139.110 1044.470 ;
        RECT 136.330 1041.690 137.510 1042.870 ;
        RECT 137.930 1041.690 139.110 1042.870 ;
        RECT 316.330 3547.010 317.510 3548.190 ;
        RECT 317.930 3547.010 319.110 3548.190 ;
        RECT 316.330 3545.410 317.510 3546.590 ;
        RECT 317.930 3545.410 319.110 3546.590 ;
        RECT 316.330 3383.290 317.510 3384.470 ;
        RECT 317.930 3383.290 319.110 3384.470 ;
        RECT 316.330 3381.690 317.510 3382.870 ;
        RECT 317.930 3381.690 319.110 3382.870 ;
        RECT 316.330 3203.290 317.510 3204.470 ;
        RECT 317.930 3203.290 319.110 3204.470 ;
        RECT 316.330 3201.690 317.510 3202.870 ;
        RECT 317.930 3201.690 319.110 3202.870 ;
        RECT 316.330 3023.290 317.510 3024.470 ;
        RECT 317.930 3023.290 319.110 3024.470 ;
        RECT 316.330 3021.690 317.510 3022.870 ;
        RECT 317.930 3021.690 319.110 3022.870 ;
        RECT 316.330 2843.290 317.510 2844.470 ;
        RECT 317.930 2843.290 319.110 2844.470 ;
        RECT 316.330 2841.690 317.510 2842.870 ;
        RECT 317.930 2841.690 319.110 2842.870 ;
        RECT 316.330 2663.290 317.510 2664.470 ;
        RECT 317.930 2663.290 319.110 2664.470 ;
        RECT 316.330 2661.690 317.510 2662.870 ;
        RECT 317.930 2661.690 319.110 2662.870 ;
        RECT 316.330 2483.290 317.510 2484.470 ;
        RECT 317.930 2483.290 319.110 2484.470 ;
        RECT 316.330 2481.690 317.510 2482.870 ;
        RECT 317.930 2481.690 319.110 2482.870 ;
        RECT 316.330 2303.290 317.510 2304.470 ;
        RECT 317.930 2303.290 319.110 2304.470 ;
        RECT 316.330 2301.690 317.510 2302.870 ;
        RECT 317.930 2301.690 319.110 2302.870 ;
        RECT 316.330 2123.290 317.510 2124.470 ;
        RECT 317.930 2123.290 319.110 2124.470 ;
        RECT 316.330 2121.690 317.510 2122.870 ;
        RECT 317.930 2121.690 319.110 2122.870 ;
        RECT 316.330 1943.290 317.510 1944.470 ;
        RECT 317.930 1943.290 319.110 1944.470 ;
        RECT 316.330 1941.690 317.510 1942.870 ;
        RECT 317.930 1941.690 319.110 1942.870 ;
        RECT 316.330 1763.290 317.510 1764.470 ;
        RECT 317.930 1763.290 319.110 1764.470 ;
        RECT 316.330 1761.690 317.510 1762.870 ;
        RECT 317.930 1761.690 319.110 1762.870 ;
        RECT 316.330 1583.290 317.510 1584.470 ;
        RECT 317.930 1583.290 319.110 1584.470 ;
        RECT 316.330 1581.690 317.510 1582.870 ;
        RECT 317.930 1581.690 319.110 1582.870 ;
        RECT 316.330 1403.290 317.510 1404.470 ;
        RECT 317.930 1403.290 319.110 1404.470 ;
        RECT 316.330 1401.690 317.510 1402.870 ;
        RECT 317.930 1401.690 319.110 1402.870 ;
        RECT 316.330 1223.290 317.510 1224.470 ;
        RECT 317.930 1223.290 319.110 1224.470 ;
        RECT 316.330 1221.690 317.510 1222.870 ;
        RECT 317.930 1221.690 319.110 1222.870 ;
        RECT 316.330 1043.290 317.510 1044.470 ;
        RECT 317.930 1043.290 319.110 1044.470 ;
        RECT 316.330 1041.690 317.510 1042.870 ;
        RECT 317.930 1041.690 319.110 1042.870 ;
        RECT 496.330 3547.010 497.510 3548.190 ;
        RECT 497.930 3547.010 499.110 3548.190 ;
        RECT 496.330 3545.410 497.510 3546.590 ;
        RECT 497.930 3545.410 499.110 3546.590 ;
        RECT 496.330 3383.290 497.510 3384.470 ;
        RECT 497.930 3383.290 499.110 3384.470 ;
        RECT 496.330 3381.690 497.510 3382.870 ;
        RECT 497.930 3381.690 499.110 3382.870 ;
        RECT 496.330 3203.290 497.510 3204.470 ;
        RECT 497.930 3203.290 499.110 3204.470 ;
        RECT 496.330 3201.690 497.510 3202.870 ;
        RECT 497.930 3201.690 499.110 3202.870 ;
        RECT 496.330 3023.290 497.510 3024.470 ;
        RECT 497.930 3023.290 499.110 3024.470 ;
        RECT 496.330 3021.690 497.510 3022.870 ;
        RECT 497.930 3021.690 499.110 3022.870 ;
        RECT 496.330 2843.290 497.510 2844.470 ;
        RECT 497.930 2843.290 499.110 2844.470 ;
        RECT 496.330 2841.690 497.510 2842.870 ;
        RECT 497.930 2841.690 499.110 2842.870 ;
        RECT 496.330 2663.290 497.510 2664.470 ;
        RECT 497.930 2663.290 499.110 2664.470 ;
        RECT 496.330 2661.690 497.510 2662.870 ;
        RECT 497.930 2661.690 499.110 2662.870 ;
        RECT 496.330 2483.290 497.510 2484.470 ;
        RECT 497.930 2483.290 499.110 2484.470 ;
        RECT 496.330 2481.690 497.510 2482.870 ;
        RECT 497.930 2481.690 499.110 2482.870 ;
        RECT 496.330 2303.290 497.510 2304.470 ;
        RECT 497.930 2303.290 499.110 2304.470 ;
        RECT 496.330 2301.690 497.510 2302.870 ;
        RECT 497.930 2301.690 499.110 2302.870 ;
        RECT 496.330 2123.290 497.510 2124.470 ;
        RECT 497.930 2123.290 499.110 2124.470 ;
        RECT 496.330 2121.690 497.510 2122.870 ;
        RECT 497.930 2121.690 499.110 2122.870 ;
        RECT 496.330 1943.290 497.510 1944.470 ;
        RECT 497.930 1943.290 499.110 1944.470 ;
        RECT 496.330 1941.690 497.510 1942.870 ;
        RECT 497.930 1941.690 499.110 1942.870 ;
        RECT 496.330 1763.290 497.510 1764.470 ;
        RECT 497.930 1763.290 499.110 1764.470 ;
        RECT 496.330 1761.690 497.510 1762.870 ;
        RECT 497.930 1761.690 499.110 1762.870 ;
        RECT 496.330 1583.290 497.510 1584.470 ;
        RECT 497.930 1583.290 499.110 1584.470 ;
        RECT 496.330 1581.690 497.510 1582.870 ;
        RECT 497.930 1581.690 499.110 1582.870 ;
        RECT 496.330 1403.290 497.510 1404.470 ;
        RECT 497.930 1403.290 499.110 1404.470 ;
        RECT 496.330 1401.690 497.510 1402.870 ;
        RECT 497.930 1401.690 499.110 1402.870 ;
        RECT 496.330 1223.290 497.510 1224.470 ;
        RECT 497.930 1223.290 499.110 1224.470 ;
        RECT 496.330 1221.690 497.510 1222.870 ;
        RECT 497.930 1221.690 499.110 1222.870 ;
        RECT 496.330 1043.290 497.510 1044.470 ;
        RECT 497.930 1043.290 499.110 1044.470 ;
        RECT 496.330 1041.690 497.510 1042.870 ;
        RECT 497.930 1041.690 499.110 1042.870 ;
        RECT 676.330 3547.010 677.510 3548.190 ;
        RECT 677.930 3547.010 679.110 3548.190 ;
        RECT 676.330 3545.410 677.510 3546.590 ;
        RECT 677.930 3545.410 679.110 3546.590 ;
        RECT 676.330 3383.290 677.510 3384.470 ;
        RECT 677.930 3383.290 679.110 3384.470 ;
        RECT 676.330 3381.690 677.510 3382.870 ;
        RECT 677.930 3381.690 679.110 3382.870 ;
        RECT 676.330 3203.290 677.510 3204.470 ;
        RECT 677.930 3203.290 679.110 3204.470 ;
        RECT 676.330 3201.690 677.510 3202.870 ;
        RECT 677.930 3201.690 679.110 3202.870 ;
        RECT 676.330 3023.290 677.510 3024.470 ;
        RECT 677.930 3023.290 679.110 3024.470 ;
        RECT 676.330 3021.690 677.510 3022.870 ;
        RECT 677.930 3021.690 679.110 3022.870 ;
        RECT 676.330 2843.290 677.510 2844.470 ;
        RECT 677.930 2843.290 679.110 2844.470 ;
        RECT 676.330 2841.690 677.510 2842.870 ;
        RECT 677.930 2841.690 679.110 2842.870 ;
        RECT 676.330 2663.290 677.510 2664.470 ;
        RECT 677.930 2663.290 679.110 2664.470 ;
        RECT 676.330 2661.690 677.510 2662.870 ;
        RECT 677.930 2661.690 679.110 2662.870 ;
        RECT 676.330 2483.290 677.510 2484.470 ;
        RECT 677.930 2483.290 679.110 2484.470 ;
        RECT 676.330 2481.690 677.510 2482.870 ;
        RECT 677.930 2481.690 679.110 2482.870 ;
        RECT 676.330 2303.290 677.510 2304.470 ;
        RECT 677.930 2303.290 679.110 2304.470 ;
        RECT 676.330 2301.690 677.510 2302.870 ;
        RECT 677.930 2301.690 679.110 2302.870 ;
        RECT 676.330 2123.290 677.510 2124.470 ;
        RECT 677.930 2123.290 679.110 2124.470 ;
        RECT 676.330 2121.690 677.510 2122.870 ;
        RECT 677.930 2121.690 679.110 2122.870 ;
        RECT 676.330 1943.290 677.510 1944.470 ;
        RECT 677.930 1943.290 679.110 1944.470 ;
        RECT 676.330 1941.690 677.510 1942.870 ;
        RECT 677.930 1941.690 679.110 1942.870 ;
        RECT 676.330 1763.290 677.510 1764.470 ;
        RECT 677.930 1763.290 679.110 1764.470 ;
        RECT 676.330 1761.690 677.510 1762.870 ;
        RECT 677.930 1761.690 679.110 1762.870 ;
        RECT 676.330 1583.290 677.510 1584.470 ;
        RECT 677.930 1583.290 679.110 1584.470 ;
        RECT 676.330 1581.690 677.510 1582.870 ;
        RECT 677.930 1581.690 679.110 1582.870 ;
        RECT 676.330 1403.290 677.510 1404.470 ;
        RECT 677.930 1403.290 679.110 1404.470 ;
        RECT 676.330 1401.690 677.510 1402.870 ;
        RECT 677.930 1401.690 679.110 1402.870 ;
        RECT 676.330 1223.290 677.510 1224.470 ;
        RECT 677.930 1223.290 679.110 1224.470 ;
        RECT 676.330 1221.690 677.510 1222.870 ;
        RECT 677.930 1221.690 679.110 1222.870 ;
        RECT 676.330 1043.290 677.510 1044.470 ;
        RECT 677.930 1043.290 679.110 1044.470 ;
        RECT 676.330 1041.690 677.510 1042.870 ;
        RECT 677.930 1041.690 679.110 1042.870 ;
        RECT 856.330 3547.010 857.510 3548.190 ;
        RECT 857.930 3547.010 859.110 3548.190 ;
        RECT 856.330 3545.410 857.510 3546.590 ;
        RECT 857.930 3545.410 859.110 3546.590 ;
        RECT 856.330 3383.290 857.510 3384.470 ;
        RECT 857.930 3383.290 859.110 3384.470 ;
        RECT 856.330 3381.690 857.510 3382.870 ;
        RECT 857.930 3381.690 859.110 3382.870 ;
        RECT 856.330 3203.290 857.510 3204.470 ;
        RECT 857.930 3203.290 859.110 3204.470 ;
        RECT 856.330 3201.690 857.510 3202.870 ;
        RECT 857.930 3201.690 859.110 3202.870 ;
        RECT 856.330 3023.290 857.510 3024.470 ;
        RECT 857.930 3023.290 859.110 3024.470 ;
        RECT 856.330 3021.690 857.510 3022.870 ;
        RECT 857.930 3021.690 859.110 3022.870 ;
        RECT 856.330 2843.290 857.510 2844.470 ;
        RECT 857.930 2843.290 859.110 2844.470 ;
        RECT 856.330 2841.690 857.510 2842.870 ;
        RECT 857.930 2841.690 859.110 2842.870 ;
        RECT 856.330 2663.290 857.510 2664.470 ;
        RECT 857.930 2663.290 859.110 2664.470 ;
        RECT 856.330 2661.690 857.510 2662.870 ;
        RECT 857.930 2661.690 859.110 2662.870 ;
        RECT 856.330 2483.290 857.510 2484.470 ;
        RECT 857.930 2483.290 859.110 2484.470 ;
        RECT 856.330 2481.690 857.510 2482.870 ;
        RECT 857.930 2481.690 859.110 2482.870 ;
        RECT 856.330 2303.290 857.510 2304.470 ;
        RECT 857.930 2303.290 859.110 2304.470 ;
        RECT 856.330 2301.690 857.510 2302.870 ;
        RECT 857.930 2301.690 859.110 2302.870 ;
        RECT 856.330 2123.290 857.510 2124.470 ;
        RECT 857.930 2123.290 859.110 2124.470 ;
        RECT 856.330 2121.690 857.510 2122.870 ;
        RECT 857.930 2121.690 859.110 2122.870 ;
        RECT 856.330 1943.290 857.510 1944.470 ;
        RECT 857.930 1943.290 859.110 1944.470 ;
        RECT 856.330 1941.690 857.510 1942.870 ;
        RECT 857.930 1941.690 859.110 1942.870 ;
        RECT 856.330 1763.290 857.510 1764.470 ;
        RECT 857.930 1763.290 859.110 1764.470 ;
        RECT 856.330 1761.690 857.510 1762.870 ;
        RECT 857.930 1761.690 859.110 1762.870 ;
        RECT 856.330 1583.290 857.510 1584.470 ;
        RECT 857.930 1583.290 859.110 1584.470 ;
        RECT 856.330 1581.690 857.510 1582.870 ;
        RECT 857.930 1581.690 859.110 1582.870 ;
        RECT 856.330 1403.290 857.510 1404.470 ;
        RECT 857.930 1403.290 859.110 1404.470 ;
        RECT 856.330 1401.690 857.510 1402.870 ;
        RECT 857.930 1401.690 859.110 1402.870 ;
        RECT 856.330 1223.290 857.510 1224.470 ;
        RECT 857.930 1223.290 859.110 1224.470 ;
        RECT 856.330 1221.690 857.510 1222.870 ;
        RECT 857.930 1221.690 859.110 1222.870 ;
        RECT 856.330 1043.290 857.510 1044.470 ;
        RECT 857.930 1043.290 859.110 1044.470 ;
        RECT 856.330 1041.690 857.510 1042.870 ;
        RECT 857.930 1041.690 859.110 1042.870 ;
        RECT 1036.330 3547.010 1037.510 3548.190 ;
        RECT 1037.930 3547.010 1039.110 3548.190 ;
        RECT 1036.330 3545.410 1037.510 3546.590 ;
        RECT 1037.930 3545.410 1039.110 3546.590 ;
        RECT 1036.330 3383.290 1037.510 3384.470 ;
        RECT 1037.930 3383.290 1039.110 3384.470 ;
        RECT 1036.330 3381.690 1037.510 3382.870 ;
        RECT 1037.930 3381.690 1039.110 3382.870 ;
        RECT 1036.330 3203.290 1037.510 3204.470 ;
        RECT 1037.930 3203.290 1039.110 3204.470 ;
        RECT 1036.330 3201.690 1037.510 3202.870 ;
        RECT 1037.930 3201.690 1039.110 3202.870 ;
        RECT 1036.330 3023.290 1037.510 3024.470 ;
        RECT 1037.930 3023.290 1039.110 3024.470 ;
        RECT 1036.330 3021.690 1037.510 3022.870 ;
        RECT 1037.930 3021.690 1039.110 3022.870 ;
        RECT 1036.330 2843.290 1037.510 2844.470 ;
        RECT 1037.930 2843.290 1039.110 2844.470 ;
        RECT 1036.330 2841.690 1037.510 2842.870 ;
        RECT 1037.930 2841.690 1039.110 2842.870 ;
        RECT 1036.330 2663.290 1037.510 2664.470 ;
        RECT 1037.930 2663.290 1039.110 2664.470 ;
        RECT 1036.330 2661.690 1037.510 2662.870 ;
        RECT 1037.930 2661.690 1039.110 2662.870 ;
        RECT 1036.330 2483.290 1037.510 2484.470 ;
        RECT 1037.930 2483.290 1039.110 2484.470 ;
        RECT 1036.330 2481.690 1037.510 2482.870 ;
        RECT 1037.930 2481.690 1039.110 2482.870 ;
        RECT 1036.330 2303.290 1037.510 2304.470 ;
        RECT 1037.930 2303.290 1039.110 2304.470 ;
        RECT 1036.330 2301.690 1037.510 2302.870 ;
        RECT 1037.930 2301.690 1039.110 2302.870 ;
        RECT 1036.330 2123.290 1037.510 2124.470 ;
        RECT 1037.930 2123.290 1039.110 2124.470 ;
        RECT 1036.330 2121.690 1037.510 2122.870 ;
        RECT 1037.930 2121.690 1039.110 2122.870 ;
        RECT 1036.330 1943.290 1037.510 1944.470 ;
        RECT 1037.930 1943.290 1039.110 1944.470 ;
        RECT 1036.330 1941.690 1037.510 1942.870 ;
        RECT 1037.930 1941.690 1039.110 1942.870 ;
        RECT 1036.330 1763.290 1037.510 1764.470 ;
        RECT 1037.930 1763.290 1039.110 1764.470 ;
        RECT 1036.330 1761.690 1037.510 1762.870 ;
        RECT 1037.930 1761.690 1039.110 1762.870 ;
        RECT 1036.330 1583.290 1037.510 1584.470 ;
        RECT 1037.930 1583.290 1039.110 1584.470 ;
        RECT 1036.330 1581.690 1037.510 1582.870 ;
        RECT 1037.930 1581.690 1039.110 1582.870 ;
        RECT 1036.330 1403.290 1037.510 1404.470 ;
        RECT 1037.930 1403.290 1039.110 1404.470 ;
        RECT 1036.330 1401.690 1037.510 1402.870 ;
        RECT 1037.930 1401.690 1039.110 1402.870 ;
        RECT 1036.330 1223.290 1037.510 1224.470 ;
        RECT 1037.930 1223.290 1039.110 1224.470 ;
        RECT 1036.330 1221.690 1037.510 1222.870 ;
        RECT 1037.930 1221.690 1039.110 1222.870 ;
        RECT 1036.330 1043.290 1037.510 1044.470 ;
        RECT 1037.930 1043.290 1039.110 1044.470 ;
        RECT 1036.330 1041.690 1037.510 1042.870 ;
        RECT 1037.930 1041.690 1039.110 1042.870 ;
        RECT 1216.330 3547.010 1217.510 3548.190 ;
        RECT 1217.930 3547.010 1219.110 3548.190 ;
        RECT 1216.330 3545.410 1217.510 3546.590 ;
        RECT 1217.930 3545.410 1219.110 3546.590 ;
        RECT 1216.330 3383.290 1217.510 3384.470 ;
        RECT 1217.930 3383.290 1219.110 3384.470 ;
        RECT 1216.330 3381.690 1217.510 3382.870 ;
        RECT 1217.930 3381.690 1219.110 3382.870 ;
        RECT 1216.330 3203.290 1217.510 3204.470 ;
        RECT 1217.930 3203.290 1219.110 3204.470 ;
        RECT 1216.330 3201.690 1217.510 3202.870 ;
        RECT 1217.930 3201.690 1219.110 3202.870 ;
        RECT 1216.330 3023.290 1217.510 3024.470 ;
        RECT 1217.930 3023.290 1219.110 3024.470 ;
        RECT 1216.330 3021.690 1217.510 3022.870 ;
        RECT 1217.930 3021.690 1219.110 3022.870 ;
        RECT 1216.330 2843.290 1217.510 2844.470 ;
        RECT 1217.930 2843.290 1219.110 2844.470 ;
        RECT 1216.330 2841.690 1217.510 2842.870 ;
        RECT 1217.930 2841.690 1219.110 2842.870 ;
        RECT 1216.330 2663.290 1217.510 2664.470 ;
        RECT 1217.930 2663.290 1219.110 2664.470 ;
        RECT 1216.330 2661.690 1217.510 2662.870 ;
        RECT 1217.930 2661.690 1219.110 2662.870 ;
        RECT 1216.330 2483.290 1217.510 2484.470 ;
        RECT 1217.930 2483.290 1219.110 2484.470 ;
        RECT 1216.330 2481.690 1217.510 2482.870 ;
        RECT 1217.930 2481.690 1219.110 2482.870 ;
        RECT 1216.330 2303.290 1217.510 2304.470 ;
        RECT 1217.930 2303.290 1219.110 2304.470 ;
        RECT 1216.330 2301.690 1217.510 2302.870 ;
        RECT 1217.930 2301.690 1219.110 2302.870 ;
        RECT 1216.330 2123.290 1217.510 2124.470 ;
        RECT 1217.930 2123.290 1219.110 2124.470 ;
        RECT 1216.330 2121.690 1217.510 2122.870 ;
        RECT 1217.930 2121.690 1219.110 2122.870 ;
        RECT 1216.330 1943.290 1217.510 1944.470 ;
        RECT 1217.930 1943.290 1219.110 1944.470 ;
        RECT 1216.330 1941.690 1217.510 1942.870 ;
        RECT 1217.930 1941.690 1219.110 1942.870 ;
        RECT 1216.330 1763.290 1217.510 1764.470 ;
        RECT 1217.930 1763.290 1219.110 1764.470 ;
        RECT 1216.330 1761.690 1217.510 1762.870 ;
        RECT 1217.930 1761.690 1219.110 1762.870 ;
        RECT 1216.330 1583.290 1217.510 1584.470 ;
        RECT 1217.930 1583.290 1219.110 1584.470 ;
        RECT 1216.330 1581.690 1217.510 1582.870 ;
        RECT 1217.930 1581.690 1219.110 1582.870 ;
        RECT 1216.330 1403.290 1217.510 1404.470 ;
        RECT 1217.930 1403.290 1219.110 1404.470 ;
        RECT 1216.330 1401.690 1217.510 1402.870 ;
        RECT 1217.930 1401.690 1219.110 1402.870 ;
        RECT 1216.330 1223.290 1217.510 1224.470 ;
        RECT 1217.930 1223.290 1219.110 1224.470 ;
        RECT 1216.330 1221.690 1217.510 1222.870 ;
        RECT 1217.930 1221.690 1219.110 1222.870 ;
        RECT 1216.330 1043.290 1217.510 1044.470 ;
        RECT 1217.930 1043.290 1219.110 1044.470 ;
        RECT 1216.330 1041.690 1217.510 1042.870 ;
        RECT 1217.930 1041.690 1219.110 1042.870 ;
        RECT 136.330 863.290 137.510 864.470 ;
        RECT 137.930 863.290 139.110 864.470 ;
        RECT 136.330 861.690 137.510 862.870 ;
        RECT 137.930 861.690 139.110 862.870 ;
        RECT 136.330 683.290 137.510 684.470 ;
        RECT 137.930 683.290 139.110 684.470 ;
        RECT 136.330 681.690 137.510 682.870 ;
        RECT 137.930 681.690 139.110 682.870 ;
        RECT 136.330 503.290 137.510 504.470 ;
        RECT 137.930 503.290 139.110 504.470 ;
        RECT 136.330 501.690 137.510 502.870 ;
        RECT 137.930 501.690 139.110 502.870 ;
        RECT 1216.330 863.290 1217.510 864.470 ;
        RECT 1217.930 863.290 1219.110 864.470 ;
        RECT 1216.330 861.690 1217.510 862.870 ;
        RECT 1217.930 861.690 1219.110 862.870 ;
        RECT 1216.330 683.290 1217.510 684.470 ;
        RECT 1217.930 683.290 1219.110 684.470 ;
        RECT 1216.330 681.690 1217.510 682.870 ;
        RECT 1217.930 681.690 1219.110 682.870 ;
        RECT 1216.330 503.290 1217.510 504.470 ;
        RECT 1217.930 503.290 1219.110 504.470 ;
        RECT 1216.330 501.690 1217.510 502.870 ;
        RECT 1217.930 501.690 1219.110 502.870 ;
        RECT 136.330 323.290 137.510 324.470 ;
        RECT 137.930 323.290 139.110 324.470 ;
        RECT 136.330 321.690 137.510 322.870 ;
        RECT 137.930 321.690 139.110 322.870 ;
        RECT 136.330 143.290 137.510 144.470 ;
        RECT 137.930 143.290 139.110 144.470 ;
        RECT 136.330 141.690 137.510 142.870 ;
        RECT 137.930 141.690 139.110 142.870 ;
        RECT 136.330 -26.910 137.510 -25.730 ;
        RECT 137.930 -26.910 139.110 -25.730 ;
        RECT 136.330 -28.510 137.510 -27.330 ;
        RECT 137.930 -28.510 139.110 -27.330 ;
        RECT 316.330 323.290 317.510 324.470 ;
        RECT 317.930 323.290 319.110 324.470 ;
        RECT 316.330 321.690 317.510 322.870 ;
        RECT 317.930 321.690 319.110 322.870 ;
        RECT 316.330 143.290 317.510 144.470 ;
        RECT 317.930 143.290 319.110 144.470 ;
        RECT 316.330 141.690 317.510 142.870 ;
        RECT 317.930 141.690 319.110 142.870 ;
        RECT 316.330 -26.910 317.510 -25.730 ;
        RECT 317.930 -26.910 319.110 -25.730 ;
        RECT 316.330 -28.510 317.510 -27.330 ;
        RECT 317.930 -28.510 319.110 -27.330 ;
        RECT 496.330 323.290 497.510 324.470 ;
        RECT 497.930 323.290 499.110 324.470 ;
        RECT 496.330 321.690 497.510 322.870 ;
        RECT 497.930 321.690 499.110 322.870 ;
        RECT 496.330 143.290 497.510 144.470 ;
        RECT 497.930 143.290 499.110 144.470 ;
        RECT 496.330 141.690 497.510 142.870 ;
        RECT 497.930 141.690 499.110 142.870 ;
        RECT 496.330 -26.910 497.510 -25.730 ;
        RECT 497.930 -26.910 499.110 -25.730 ;
        RECT 496.330 -28.510 497.510 -27.330 ;
        RECT 497.930 -28.510 499.110 -27.330 ;
        RECT 676.330 323.290 677.510 324.470 ;
        RECT 677.930 323.290 679.110 324.470 ;
        RECT 676.330 321.690 677.510 322.870 ;
        RECT 677.930 321.690 679.110 322.870 ;
        RECT 676.330 143.290 677.510 144.470 ;
        RECT 677.930 143.290 679.110 144.470 ;
        RECT 676.330 141.690 677.510 142.870 ;
        RECT 677.930 141.690 679.110 142.870 ;
        RECT 676.330 -26.910 677.510 -25.730 ;
        RECT 677.930 -26.910 679.110 -25.730 ;
        RECT 676.330 -28.510 677.510 -27.330 ;
        RECT 677.930 -28.510 679.110 -27.330 ;
        RECT 856.330 323.290 857.510 324.470 ;
        RECT 857.930 323.290 859.110 324.470 ;
        RECT 856.330 321.690 857.510 322.870 ;
        RECT 857.930 321.690 859.110 322.870 ;
        RECT 856.330 143.290 857.510 144.470 ;
        RECT 857.930 143.290 859.110 144.470 ;
        RECT 856.330 141.690 857.510 142.870 ;
        RECT 857.930 141.690 859.110 142.870 ;
        RECT 856.330 -26.910 857.510 -25.730 ;
        RECT 857.930 -26.910 859.110 -25.730 ;
        RECT 856.330 -28.510 857.510 -27.330 ;
        RECT 857.930 -28.510 859.110 -27.330 ;
        RECT 1036.330 323.290 1037.510 324.470 ;
        RECT 1037.930 323.290 1039.110 324.470 ;
        RECT 1036.330 321.690 1037.510 322.870 ;
        RECT 1037.930 321.690 1039.110 322.870 ;
        RECT 1036.330 143.290 1037.510 144.470 ;
        RECT 1037.930 143.290 1039.110 144.470 ;
        RECT 1036.330 141.690 1037.510 142.870 ;
        RECT 1037.930 141.690 1039.110 142.870 ;
        RECT 1036.330 -26.910 1037.510 -25.730 ;
        RECT 1037.930 -26.910 1039.110 -25.730 ;
        RECT 1036.330 -28.510 1037.510 -27.330 ;
        RECT 1037.930 -28.510 1039.110 -27.330 ;
        RECT 1216.330 323.290 1217.510 324.470 ;
        RECT 1217.930 323.290 1219.110 324.470 ;
        RECT 1216.330 321.690 1217.510 322.870 ;
        RECT 1217.930 321.690 1219.110 322.870 ;
        RECT 1216.330 143.290 1217.510 144.470 ;
        RECT 1217.930 143.290 1219.110 144.470 ;
        RECT 1216.330 141.690 1217.510 142.870 ;
        RECT 1217.930 141.690 1219.110 142.870 ;
        RECT 1216.330 -26.910 1217.510 -25.730 ;
        RECT 1217.930 -26.910 1219.110 -25.730 ;
        RECT 1216.330 -28.510 1217.510 -27.330 ;
        RECT 1217.930 -28.510 1219.110 -27.330 ;
        RECT 1396.330 3547.010 1397.510 3548.190 ;
        RECT 1397.930 3547.010 1399.110 3548.190 ;
        RECT 1396.330 3545.410 1397.510 3546.590 ;
        RECT 1397.930 3545.410 1399.110 3546.590 ;
        RECT 1396.330 3383.290 1397.510 3384.470 ;
        RECT 1397.930 3383.290 1399.110 3384.470 ;
        RECT 1396.330 3381.690 1397.510 3382.870 ;
        RECT 1397.930 3381.690 1399.110 3382.870 ;
        RECT 1396.330 3203.290 1397.510 3204.470 ;
        RECT 1397.930 3203.290 1399.110 3204.470 ;
        RECT 1396.330 3201.690 1397.510 3202.870 ;
        RECT 1397.930 3201.690 1399.110 3202.870 ;
        RECT 1396.330 3023.290 1397.510 3024.470 ;
        RECT 1397.930 3023.290 1399.110 3024.470 ;
        RECT 1396.330 3021.690 1397.510 3022.870 ;
        RECT 1397.930 3021.690 1399.110 3022.870 ;
        RECT 1396.330 2843.290 1397.510 2844.470 ;
        RECT 1397.930 2843.290 1399.110 2844.470 ;
        RECT 1396.330 2841.690 1397.510 2842.870 ;
        RECT 1397.930 2841.690 1399.110 2842.870 ;
        RECT 1396.330 2663.290 1397.510 2664.470 ;
        RECT 1397.930 2663.290 1399.110 2664.470 ;
        RECT 1396.330 2661.690 1397.510 2662.870 ;
        RECT 1397.930 2661.690 1399.110 2662.870 ;
        RECT 1396.330 2483.290 1397.510 2484.470 ;
        RECT 1397.930 2483.290 1399.110 2484.470 ;
        RECT 1396.330 2481.690 1397.510 2482.870 ;
        RECT 1397.930 2481.690 1399.110 2482.870 ;
        RECT 1396.330 2303.290 1397.510 2304.470 ;
        RECT 1397.930 2303.290 1399.110 2304.470 ;
        RECT 1396.330 2301.690 1397.510 2302.870 ;
        RECT 1397.930 2301.690 1399.110 2302.870 ;
        RECT 1396.330 2123.290 1397.510 2124.470 ;
        RECT 1397.930 2123.290 1399.110 2124.470 ;
        RECT 1396.330 2121.690 1397.510 2122.870 ;
        RECT 1397.930 2121.690 1399.110 2122.870 ;
        RECT 1396.330 1943.290 1397.510 1944.470 ;
        RECT 1397.930 1943.290 1399.110 1944.470 ;
        RECT 1396.330 1941.690 1397.510 1942.870 ;
        RECT 1397.930 1941.690 1399.110 1942.870 ;
        RECT 1396.330 1763.290 1397.510 1764.470 ;
        RECT 1397.930 1763.290 1399.110 1764.470 ;
        RECT 1396.330 1761.690 1397.510 1762.870 ;
        RECT 1397.930 1761.690 1399.110 1762.870 ;
        RECT 1396.330 1583.290 1397.510 1584.470 ;
        RECT 1397.930 1583.290 1399.110 1584.470 ;
        RECT 1396.330 1581.690 1397.510 1582.870 ;
        RECT 1397.930 1581.690 1399.110 1582.870 ;
        RECT 1396.330 1403.290 1397.510 1404.470 ;
        RECT 1397.930 1403.290 1399.110 1404.470 ;
        RECT 1396.330 1401.690 1397.510 1402.870 ;
        RECT 1397.930 1401.690 1399.110 1402.870 ;
        RECT 1396.330 1223.290 1397.510 1224.470 ;
        RECT 1397.930 1223.290 1399.110 1224.470 ;
        RECT 1396.330 1221.690 1397.510 1222.870 ;
        RECT 1397.930 1221.690 1399.110 1222.870 ;
        RECT 1396.330 1043.290 1397.510 1044.470 ;
        RECT 1397.930 1043.290 1399.110 1044.470 ;
        RECT 1396.330 1041.690 1397.510 1042.870 ;
        RECT 1397.930 1041.690 1399.110 1042.870 ;
        RECT 1396.330 863.290 1397.510 864.470 ;
        RECT 1397.930 863.290 1399.110 864.470 ;
        RECT 1396.330 861.690 1397.510 862.870 ;
        RECT 1397.930 861.690 1399.110 862.870 ;
        RECT 1396.330 683.290 1397.510 684.470 ;
        RECT 1397.930 683.290 1399.110 684.470 ;
        RECT 1396.330 681.690 1397.510 682.870 ;
        RECT 1397.930 681.690 1399.110 682.870 ;
        RECT 1396.330 503.290 1397.510 504.470 ;
        RECT 1397.930 503.290 1399.110 504.470 ;
        RECT 1396.330 501.690 1397.510 502.870 ;
        RECT 1397.930 501.690 1399.110 502.870 ;
        RECT 1396.330 323.290 1397.510 324.470 ;
        RECT 1397.930 323.290 1399.110 324.470 ;
        RECT 1396.330 321.690 1397.510 322.870 ;
        RECT 1397.930 321.690 1399.110 322.870 ;
        RECT 1396.330 143.290 1397.510 144.470 ;
        RECT 1397.930 143.290 1399.110 144.470 ;
        RECT 1396.330 141.690 1397.510 142.870 ;
        RECT 1397.930 141.690 1399.110 142.870 ;
        RECT 1396.330 -26.910 1397.510 -25.730 ;
        RECT 1397.930 -26.910 1399.110 -25.730 ;
        RECT 1396.330 -28.510 1397.510 -27.330 ;
        RECT 1397.930 -28.510 1399.110 -27.330 ;
        RECT 1576.330 3547.010 1577.510 3548.190 ;
        RECT 1577.930 3547.010 1579.110 3548.190 ;
        RECT 1576.330 3545.410 1577.510 3546.590 ;
        RECT 1577.930 3545.410 1579.110 3546.590 ;
        RECT 1576.330 3383.290 1577.510 3384.470 ;
        RECT 1577.930 3383.290 1579.110 3384.470 ;
        RECT 1576.330 3381.690 1577.510 3382.870 ;
        RECT 1577.930 3381.690 1579.110 3382.870 ;
        RECT 1576.330 3203.290 1577.510 3204.470 ;
        RECT 1577.930 3203.290 1579.110 3204.470 ;
        RECT 1576.330 3201.690 1577.510 3202.870 ;
        RECT 1577.930 3201.690 1579.110 3202.870 ;
        RECT 1576.330 3023.290 1577.510 3024.470 ;
        RECT 1577.930 3023.290 1579.110 3024.470 ;
        RECT 1576.330 3021.690 1577.510 3022.870 ;
        RECT 1577.930 3021.690 1579.110 3022.870 ;
        RECT 1576.330 2843.290 1577.510 2844.470 ;
        RECT 1577.930 2843.290 1579.110 2844.470 ;
        RECT 1576.330 2841.690 1577.510 2842.870 ;
        RECT 1577.930 2841.690 1579.110 2842.870 ;
        RECT 1576.330 2663.290 1577.510 2664.470 ;
        RECT 1577.930 2663.290 1579.110 2664.470 ;
        RECT 1576.330 2661.690 1577.510 2662.870 ;
        RECT 1577.930 2661.690 1579.110 2662.870 ;
        RECT 1576.330 2483.290 1577.510 2484.470 ;
        RECT 1577.930 2483.290 1579.110 2484.470 ;
        RECT 1576.330 2481.690 1577.510 2482.870 ;
        RECT 1577.930 2481.690 1579.110 2482.870 ;
        RECT 1576.330 2303.290 1577.510 2304.470 ;
        RECT 1577.930 2303.290 1579.110 2304.470 ;
        RECT 1576.330 2301.690 1577.510 2302.870 ;
        RECT 1577.930 2301.690 1579.110 2302.870 ;
        RECT 1576.330 2123.290 1577.510 2124.470 ;
        RECT 1577.930 2123.290 1579.110 2124.470 ;
        RECT 1576.330 2121.690 1577.510 2122.870 ;
        RECT 1577.930 2121.690 1579.110 2122.870 ;
        RECT 1576.330 1943.290 1577.510 1944.470 ;
        RECT 1577.930 1943.290 1579.110 1944.470 ;
        RECT 1576.330 1941.690 1577.510 1942.870 ;
        RECT 1577.930 1941.690 1579.110 1942.870 ;
        RECT 1576.330 1763.290 1577.510 1764.470 ;
        RECT 1577.930 1763.290 1579.110 1764.470 ;
        RECT 1576.330 1761.690 1577.510 1762.870 ;
        RECT 1577.930 1761.690 1579.110 1762.870 ;
        RECT 1576.330 1583.290 1577.510 1584.470 ;
        RECT 1577.930 1583.290 1579.110 1584.470 ;
        RECT 1576.330 1581.690 1577.510 1582.870 ;
        RECT 1577.930 1581.690 1579.110 1582.870 ;
        RECT 1576.330 1403.290 1577.510 1404.470 ;
        RECT 1577.930 1403.290 1579.110 1404.470 ;
        RECT 1576.330 1401.690 1577.510 1402.870 ;
        RECT 1577.930 1401.690 1579.110 1402.870 ;
        RECT 1576.330 1223.290 1577.510 1224.470 ;
        RECT 1577.930 1223.290 1579.110 1224.470 ;
        RECT 1576.330 1221.690 1577.510 1222.870 ;
        RECT 1577.930 1221.690 1579.110 1222.870 ;
        RECT 1576.330 1043.290 1577.510 1044.470 ;
        RECT 1577.930 1043.290 1579.110 1044.470 ;
        RECT 1576.330 1041.690 1577.510 1042.870 ;
        RECT 1577.930 1041.690 1579.110 1042.870 ;
        RECT 1576.330 863.290 1577.510 864.470 ;
        RECT 1577.930 863.290 1579.110 864.470 ;
        RECT 1576.330 861.690 1577.510 862.870 ;
        RECT 1577.930 861.690 1579.110 862.870 ;
        RECT 1576.330 683.290 1577.510 684.470 ;
        RECT 1577.930 683.290 1579.110 684.470 ;
        RECT 1576.330 681.690 1577.510 682.870 ;
        RECT 1577.930 681.690 1579.110 682.870 ;
        RECT 1576.330 503.290 1577.510 504.470 ;
        RECT 1577.930 503.290 1579.110 504.470 ;
        RECT 1576.330 501.690 1577.510 502.870 ;
        RECT 1577.930 501.690 1579.110 502.870 ;
        RECT 1576.330 323.290 1577.510 324.470 ;
        RECT 1577.930 323.290 1579.110 324.470 ;
        RECT 1576.330 321.690 1577.510 322.870 ;
        RECT 1577.930 321.690 1579.110 322.870 ;
        RECT 1576.330 143.290 1577.510 144.470 ;
        RECT 1577.930 143.290 1579.110 144.470 ;
        RECT 1576.330 141.690 1577.510 142.870 ;
        RECT 1577.930 141.690 1579.110 142.870 ;
        RECT 1576.330 -26.910 1577.510 -25.730 ;
        RECT 1577.930 -26.910 1579.110 -25.730 ;
        RECT 1576.330 -28.510 1577.510 -27.330 ;
        RECT 1577.930 -28.510 1579.110 -27.330 ;
        RECT 1756.330 3547.010 1757.510 3548.190 ;
        RECT 1757.930 3547.010 1759.110 3548.190 ;
        RECT 1756.330 3545.410 1757.510 3546.590 ;
        RECT 1757.930 3545.410 1759.110 3546.590 ;
        RECT 1756.330 3383.290 1757.510 3384.470 ;
        RECT 1757.930 3383.290 1759.110 3384.470 ;
        RECT 1756.330 3381.690 1757.510 3382.870 ;
        RECT 1757.930 3381.690 1759.110 3382.870 ;
        RECT 1756.330 3203.290 1757.510 3204.470 ;
        RECT 1757.930 3203.290 1759.110 3204.470 ;
        RECT 1756.330 3201.690 1757.510 3202.870 ;
        RECT 1757.930 3201.690 1759.110 3202.870 ;
        RECT 1756.330 3023.290 1757.510 3024.470 ;
        RECT 1757.930 3023.290 1759.110 3024.470 ;
        RECT 1756.330 3021.690 1757.510 3022.870 ;
        RECT 1757.930 3021.690 1759.110 3022.870 ;
        RECT 1756.330 2843.290 1757.510 2844.470 ;
        RECT 1757.930 2843.290 1759.110 2844.470 ;
        RECT 1756.330 2841.690 1757.510 2842.870 ;
        RECT 1757.930 2841.690 1759.110 2842.870 ;
        RECT 1756.330 2663.290 1757.510 2664.470 ;
        RECT 1757.930 2663.290 1759.110 2664.470 ;
        RECT 1756.330 2661.690 1757.510 2662.870 ;
        RECT 1757.930 2661.690 1759.110 2662.870 ;
        RECT 1756.330 2483.290 1757.510 2484.470 ;
        RECT 1757.930 2483.290 1759.110 2484.470 ;
        RECT 1756.330 2481.690 1757.510 2482.870 ;
        RECT 1757.930 2481.690 1759.110 2482.870 ;
        RECT 1756.330 2303.290 1757.510 2304.470 ;
        RECT 1757.930 2303.290 1759.110 2304.470 ;
        RECT 1756.330 2301.690 1757.510 2302.870 ;
        RECT 1757.930 2301.690 1759.110 2302.870 ;
        RECT 1756.330 2123.290 1757.510 2124.470 ;
        RECT 1757.930 2123.290 1759.110 2124.470 ;
        RECT 1756.330 2121.690 1757.510 2122.870 ;
        RECT 1757.930 2121.690 1759.110 2122.870 ;
        RECT 1756.330 1943.290 1757.510 1944.470 ;
        RECT 1757.930 1943.290 1759.110 1944.470 ;
        RECT 1756.330 1941.690 1757.510 1942.870 ;
        RECT 1757.930 1941.690 1759.110 1942.870 ;
        RECT 1756.330 1763.290 1757.510 1764.470 ;
        RECT 1757.930 1763.290 1759.110 1764.470 ;
        RECT 1756.330 1761.690 1757.510 1762.870 ;
        RECT 1757.930 1761.690 1759.110 1762.870 ;
        RECT 1756.330 1583.290 1757.510 1584.470 ;
        RECT 1757.930 1583.290 1759.110 1584.470 ;
        RECT 1756.330 1581.690 1757.510 1582.870 ;
        RECT 1757.930 1581.690 1759.110 1582.870 ;
        RECT 1756.330 1403.290 1757.510 1404.470 ;
        RECT 1757.930 1403.290 1759.110 1404.470 ;
        RECT 1756.330 1401.690 1757.510 1402.870 ;
        RECT 1757.930 1401.690 1759.110 1402.870 ;
        RECT 1756.330 1223.290 1757.510 1224.470 ;
        RECT 1757.930 1223.290 1759.110 1224.470 ;
        RECT 1756.330 1221.690 1757.510 1222.870 ;
        RECT 1757.930 1221.690 1759.110 1222.870 ;
        RECT 1756.330 1043.290 1757.510 1044.470 ;
        RECT 1757.930 1043.290 1759.110 1044.470 ;
        RECT 1756.330 1041.690 1757.510 1042.870 ;
        RECT 1757.930 1041.690 1759.110 1042.870 ;
        RECT 1756.330 863.290 1757.510 864.470 ;
        RECT 1757.930 863.290 1759.110 864.470 ;
        RECT 1756.330 861.690 1757.510 862.870 ;
        RECT 1757.930 861.690 1759.110 862.870 ;
        RECT 1756.330 683.290 1757.510 684.470 ;
        RECT 1757.930 683.290 1759.110 684.470 ;
        RECT 1756.330 681.690 1757.510 682.870 ;
        RECT 1757.930 681.690 1759.110 682.870 ;
        RECT 1756.330 503.290 1757.510 504.470 ;
        RECT 1757.930 503.290 1759.110 504.470 ;
        RECT 1756.330 501.690 1757.510 502.870 ;
        RECT 1757.930 501.690 1759.110 502.870 ;
        RECT 1756.330 323.290 1757.510 324.470 ;
        RECT 1757.930 323.290 1759.110 324.470 ;
        RECT 1756.330 321.690 1757.510 322.870 ;
        RECT 1757.930 321.690 1759.110 322.870 ;
        RECT 1756.330 143.290 1757.510 144.470 ;
        RECT 1757.930 143.290 1759.110 144.470 ;
        RECT 1756.330 141.690 1757.510 142.870 ;
        RECT 1757.930 141.690 1759.110 142.870 ;
        RECT 1756.330 -26.910 1757.510 -25.730 ;
        RECT 1757.930 -26.910 1759.110 -25.730 ;
        RECT 1756.330 -28.510 1757.510 -27.330 ;
        RECT 1757.930 -28.510 1759.110 -27.330 ;
        RECT 1936.330 3547.010 1937.510 3548.190 ;
        RECT 1937.930 3547.010 1939.110 3548.190 ;
        RECT 1936.330 3545.410 1937.510 3546.590 ;
        RECT 1937.930 3545.410 1939.110 3546.590 ;
        RECT 1936.330 3383.290 1937.510 3384.470 ;
        RECT 1937.930 3383.290 1939.110 3384.470 ;
        RECT 1936.330 3381.690 1937.510 3382.870 ;
        RECT 1937.930 3381.690 1939.110 3382.870 ;
        RECT 1936.330 3203.290 1937.510 3204.470 ;
        RECT 1937.930 3203.290 1939.110 3204.470 ;
        RECT 1936.330 3201.690 1937.510 3202.870 ;
        RECT 1937.930 3201.690 1939.110 3202.870 ;
        RECT 1936.330 3023.290 1937.510 3024.470 ;
        RECT 1937.930 3023.290 1939.110 3024.470 ;
        RECT 1936.330 3021.690 1937.510 3022.870 ;
        RECT 1937.930 3021.690 1939.110 3022.870 ;
        RECT 1936.330 2843.290 1937.510 2844.470 ;
        RECT 1937.930 2843.290 1939.110 2844.470 ;
        RECT 1936.330 2841.690 1937.510 2842.870 ;
        RECT 1937.930 2841.690 1939.110 2842.870 ;
        RECT 1936.330 2663.290 1937.510 2664.470 ;
        RECT 1937.930 2663.290 1939.110 2664.470 ;
        RECT 1936.330 2661.690 1937.510 2662.870 ;
        RECT 1937.930 2661.690 1939.110 2662.870 ;
        RECT 1936.330 2483.290 1937.510 2484.470 ;
        RECT 1937.930 2483.290 1939.110 2484.470 ;
        RECT 1936.330 2481.690 1937.510 2482.870 ;
        RECT 1937.930 2481.690 1939.110 2482.870 ;
        RECT 1936.330 2303.290 1937.510 2304.470 ;
        RECT 1937.930 2303.290 1939.110 2304.470 ;
        RECT 1936.330 2301.690 1937.510 2302.870 ;
        RECT 1937.930 2301.690 1939.110 2302.870 ;
        RECT 1936.330 2123.290 1937.510 2124.470 ;
        RECT 1937.930 2123.290 1939.110 2124.470 ;
        RECT 1936.330 2121.690 1937.510 2122.870 ;
        RECT 1937.930 2121.690 1939.110 2122.870 ;
        RECT 1936.330 1943.290 1937.510 1944.470 ;
        RECT 1937.930 1943.290 1939.110 1944.470 ;
        RECT 1936.330 1941.690 1937.510 1942.870 ;
        RECT 1937.930 1941.690 1939.110 1942.870 ;
        RECT 1936.330 1763.290 1937.510 1764.470 ;
        RECT 1937.930 1763.290 1939.110 1764.470 ;
        RECT 1936.330 1761.690 1937.510 1762.870 ;
        RECT 1937.930 1761.690 1939.110 1762.870 ;
        RECT 1936.330 1583.290 1937.510 1584.470 ;
        RECT 1937.930 1583.290 1939.110 1584.470 ;
        RECT 1936.330 1581.690 1937.510 1582.870 ;
        RECT 1937.930 1581.690 1939.110 1582.870 ;
        RECT 1936.330 1403.290 1937.510 1404.470 ;
        RECT 1937.930 1403.290 1939.110 1404.470 ;
        RECT 1936.330 1401.690 1937.510 1402.870 ;
        RECT 1937.930 1401.690 1939.110 1402.870 ;
        RECT 1936.330 1223.290 1937.510 1224.470 ;
        RECT 1937.930 1223.290 1939.110 1224.470 ;
        RECT 1936.330 1221.690 1937.510 1222.870 ;
        RECT 1937.930 1221.690 1939.110 1222.870 ;
        RECT 1936.330 1043.290 1937.510 1044.470 ;
        RECT 1937.930 1043.290 1939.110 1044.470 ;
        RECT 1936.330 1041.690 1937.510 1042.870 ;
        RECT 1937.930 1041.690 1939.110 1042.870 ;
        RECT 1936.330 863.290 1937.510 864.470 ;
        RECT 1937.930 863.290 1939.110 864.470 ;
        RECT 1936.330 861.690 1937.510 862.870 ;
        RECT 1937.930 861.690 1939.110 862.870 ;
        RECT 1936.330 683.290 1937.510 684.470 ;
        RECT 1937.930 683.290 1939.110 684.470 ;
        RECT 1936.330 681.690 1937.510 682.870 ;
        RECT 1937.930 681.690 1939.110 682.870 ;
        RECT 1936.330 503.290 1937.510 504.470 ;
        RECT 1937.930 503.290 1939.110 504.470 ;
        RECT 1936.330 501.690 1937.510 502.870 ;
        RECT 1937.930 501.690 1939.110 502.870 ;
        RECT 1936.330 323.290 1937.510 324.470 ;
        RECT 1937.930 323.290 1939.110 324.470 ;
        RECT 1936.330 321.690 1937.510 322.870 ;
        RECT 1937.930 321.690 1939.110 322.870 ;
        RECT 1936.330 143.290 1937.510 144.470 ;
        RECT 1937.930 143.290 1939.110 144.470 ;
        RECT 1936.330 141.690 1937.510 142.870 ;
        RECT 1937.930 141.690 1939.110 142.870 ;
        RECT 1936.330 -26.910 1937.510 -25.730 ;
        RECT 1937.930 -26.910 1939.110 -25.730 ;
        RECT 1936.330 -28.510 1937.510 -27.330 ;
        RECT 1937.930 -28.510 1939.110 -27.330 ;
        RECT 2116.330 3547.010 2117.510 3548.190 ;
        RECT 2117.930 3547.010 2119.110 3548.190 ;
        RECT 2116.330 3545.410 2117.510 3546.590 ;
        RECT 2117.930 3545.410 2119.110 3546.590 ;
        RECT 2116.330 3383.290 2117.510 3384.470 ;
        RECT 2117.930 3383.290 2119.110 3384.470 ;
        RECT 2116.330 3381.690 2117.510 3382.870 ;
        RECT 2117.930 3381.690 2119.110 3382.870 ;
        RECT 2116.330 3203.290 2117.510 3204.470 ;
        RECT 2117.930 3203.290 2119.110 3204.470 ;
        RECT 2116.330 3201.690 2117.510 3202.870 ;
        RECT 2117.930 3201.690 2119.110 3202.870 ;
        RECT 2116.330 3023.290 2117.510 3024.470 ;
        RECT 2117.930 3023.290 2119.110 3024.470 ;
        RECT 2116.330 3021.690 2117.510 3022.870 ;
        RECT 2117.930 3021.690 2119.110 3022.870 ;
        RECT 2116.330 2843.290 2117.510 2844.470 ;
        RECT 2117.930 2843.290 2119.110 2844.470 ;
        RECT 2116.330 2841.690 2117.510 2842.870 ;
        RECT 2117.930 2841.690 2119.110 2842.870 ;
        RECT 2116.330 2663.290 2117.510 2664.470 ;
        RECT 2117.930 2663.290 2119.110 2664.470 ;
        RECT 2116.330 2661.690 2117.510 2662.870 ;
        RECT 2117.930 2661.690 2119.110 2662.870 ;
        RECT 2116.330 2483.290 2117.510 2484.470 ;
        RECT 2117.930 2483.290 2119.110 2484.470 ;
        RECT 2116.330 2481.690 2117.510 2482.870 ;
        RECT 2117.930 2481.690 2119.110 2482.870 ;
        RECT 2116.330 2303.290 2117.510 2304.470 ;
        RECT 2117.930 2303.290 2119.110 2304.470 ;
        RECT 2116.330 2301.690 2117.510 2302.870 ;
        RECT 2117.930 2301.690 2119.110 2302.870 ;
        RECT 2116.330 2123.290 2117.510 2124.470 ;
        RECT 2117.930 2123.290 2119.110 2124.470 ;
        RECT 2116.330 2121.690 2117.510 2122.870 ;
        RECT 2117.930 2121.690 2119.110 2122.870 ;
        RECT 2116.330 1943.290 2117.510 1944.470 ;
        RECT 2117.930 1943.290 2119.110 1944.470 ;
        RECT 2116.330 1941.690 2117.510 1942.870 ;
        RECT 2117.930 1941.690 2119.110 1942.870 ;
        RECT 2116.330 1763.290 2117.510 1764.470 ;
        RECT 2117.930 1763.290 2119.110 1764.470 ;
        RECT 2116.330 1761.690 2117.510 1762.870 ;
        RECT 2117.930 1761.690 2119.110 1762.870 ;
        RECT 2116.330 1583.290 2117.510 1584.470 ;
        RECT 2117.930 1583.290 2119.110 1584.470 ;
        RECT 2116.330 1581.690 2117.510 1582.870 ;
        RECT 2117.930 1581.690 2119.110 1582.870 ;
        RECT 2116.330 1403.290 2117.510 1404.470 ;
        RECT 2117.930 1403.290 2119.110 1404.470 ;
        RECT 2116.330 1401.690 2117.510 1402.870 ;
        RECT 2117.930 1401.690 2119.110 1402.870 ;
        RECT 2116.330 1223.290 2117.510 1224.470 ;
        RECT 2117.930 1223.290 2119.110 1224.470 ;
        RECT 2116.330 1221.690 2117.510 1222.870 ;
        RECT 2117.930 1221.690 2119.110 1222.870 ;
        RECT 2116.330 1043.290 2117.510 1044.470 ;
        RECT 2117.930 1043.290 2119.110 1044.470 ;
        RECT 2116.330 1041.690 2117.510 1042.870 ;
        RECT 2117.930 1041.690 2119.110 1042.870 ;
        RECT 2116.330 863.290 2117.510 864.470 ;
        RECT 2117.930 863.290 2119.110 864.470 ;
        RECT 2116.330 861.690 2117.510 862.870 ;
        RECT 2117.930 861.690 2119.110 862.870 ;
        RECT 2116.330 683.290 2117.510 684.470 ;
        RECT 2117.930 683.290 2119.110 684.470 ;
        RECT 2116.330 681.690 2117.510 682.870 ;
        RECT 2117.930 681.690 2119.110 682.870 ;
        RECT 2116.330 503.290 2117.510 504.470 ;
        RECT 2117.930 503.290 2119.110 504.470 ;
        RECT 2116.330 501.690 2117.510 502.870 ;
        RECT 2117.930 501.690 2119.110 502.870 ;
        RECT 2116.330 323.290 2117.510 324.470 ;
        RECT 2117.930 323.290 2119.110 324.470 ;
        RECT 2116.330 321.690 2117.510 322.870 ;
        RECT 2117.930 321.690 2119.110 322.870 ;
        RECT 2116.330 143.290 2117.510 144.470 ;
        RECT 2117.930 143.290 2119.110 144.470 ;
        RECT 2116.330 141.690 2117.510 142.870 ;
        RECT 2117.930 141.690 2119.110 142.870 ;
        RECT 2116.330 -26.910 2117.510 -25.730 ;
        RECT 2117.930 -26.910 2119.110 -25.730 ;
        RECT 2116.330 -28.510 2117.510 -27.330 ;
        RECT 2117.930 -28.510 2119.110 -27.330 ;
        RECT 2296.330 3547.010 2297.510 3548.190 ;
        RECT 2297.930 3547.010 2299.110 3548.190 ;
        RECT 2296.330 3545.410 2297.510 3546.590 ;
        RECT 2297.930 3545.410 2299.110 3546.590 ;
        RECT 2296.330 3383.290 2297.510 3384.470 ;
        RECT 2297.930 3383.290 2299.110 3384.470 ;
        RECT 2296.330 3381.690 2297.510 3382.870 ;
        RECT 2297.930 3381.690 2299.110 3382.870 ;
        RECT 2296.330 3203.290 2297.510 3204.470 ;
        RECT 2297.930 3203.290 2299.110 3204.470 ;
        RECT 2296.330 3201.690 2297.510 3202.870 ;
        RECT 2297.930 3201.690 2299.110 3202.870 ;
        RECT 2296.330 3023.290 2297.510 3024.470 ;
        RECT 2297.930 3023.290 2299.110 3024.470 ;
        RECT 2296.330 3021.690 2297.510 3022.870 ;
        RECT 2297.930 3021.690 2299.110 3022.870 ;
        RECT 2296.330 2843.290 2297.510 2844.470 ;
        RECT 2297.930 2843.290 2299.110 2844.470 ;
        RECT 2296.330 2841.690 2297.510 2842.870 ;
        RECT 2297.930 2841.690 2299.110 2842.870 ;
        RECT 2296.330 2663.290 2297.510 2664.470 ;
        RECT 2297.930 2663.290 2299.110 2664.470 ;
        RECT 2296.330 2661.690 2297.510 2662.870 ;
        RECT 2297.930 2661.690 2299.110 2662.870 ;
        RECT 2296.330 2483.290 2297.510 2484.470 ;
        RECT 2297.930 2483.290 2299.110 2484.470 ;
        RECT 2296.330 2481.690 2297.510 2482.870 ;
        RECT 2297.930 2481.690 2299.110 2482.870 ;
        RECT 2296.330 2303.290 2297.510 2304.470 ;
        RECT 2297.930 2303.290 2299.110 2304.470 ;
        RECT 2296.330 2301.690 2297.510 2302.870 ;
        RECT 2297.930 2301.690 2299.110 2302.870 ;
        RECT 2296.330 2123.290 2297.510 2124.470 ;
        RECT 2297.930 2123.290 2299.110 2124.470 ;
        RECT 2296.330 2121.690 2297.510 2122.870 ;
        RECT 2297.930 2121.690 2299.110 2122.870 ;
        RECT 2296.330 1943.290 2297.510 1944.470 ;
        RECT 2297.930 1943.290 2299.110 1944.470 ;
        RECT 2296.330 1941.690 2297.510 1942.870 ;
        RECT 2297.930 1941.690 2299.110 1942.870 ;
        RECT 2296.330 1763.290 2297.510 1764.470 ;
        RECT 2297.930 1763.290 2299.110 1764.470 ;
        RECT 2296.330 1761.690 2297.510 1762.870 ;
        RECT 2297.930 1761.690 2299.110 1762.870 ;
        RECT 2296.330 1583.290 2297.510 1584.470 ;
        RECT 2297.930 1583.290 2299.110 1584.470 ;
        RECT 2296.330 1581.690 2297.510 1582.870 ;
        RECT 2297.930 1581.690 2299.110 1582.870 ;
        RECT 2296.330 1403.290 2297.510 1404.470 ;
        RECT 2297.930 1403.290 2299.110 1404.470 ;
        RECT 2296.330 1401.690 2297.510 1402.870 ;
        RECT 2297.930 1401.690 2299.110 1402.870 ;
        RECT 2296.330 1223.290 2297.510 1224.470 ;
        RECT 2297.930 1223.290 2299.110 1224.470 ;
        RECT 2296.330 1221.690 2297.510 1222.870 ;
        RECT 2297.930 1221.690 2299.110 1222.870 ;
        RECT 2296.330 1043.290 2297.510 1044.470 ;
        RECT 2297.930 1043.290 2299.110 1044.470 ;
        RECT 2296.330 1041.690 2297.510 1042.870 ;
        RECT 2297.930 1041.690 2299.110 1042.870 ;
        RECT 2296.330 863.290 2297.510 864.470 ;
        RECT 2297.930 863.290 2299.110 864.470 ;
        RECT 2296.330 861.690 2297.510 862.870 ;
        RECT 2297.930 861.690 2299.110 862.870 ;
        RECT 2296.330 683.290 2297.510 684.470 ;
        RECT 2297.930 683.290 2299.110 684.470 ;
        RECT 2296.330 681.690 2297.510 682.870 ;
        RECT 2297.930 681.690 2299.110 682.870 ;
        RECT 2296.330 503.290 2297.510 504.470 ;
        RECT 2297.930 503.290 2299.110 504.470 ;
        RECT 2296.330 501.690 2297.510 502.870 ;
        RECT 2297.930 501.690 2299.110 502.870 ;
        RECT 2296.330 323.290 2297.510 324.470 ;
        RECT 2297.930 323.290 2299.110 324.470 ;
        RECT 2296.330 321.690 2297.510 322.870 ;
        RECT 2297.930 321.690 2299.110 322.870 ;
        RECT 2296.330 143.290 2297.510 144.470 ;
        RECT 2297.930 143.290 2299.110 144.470 ;
        RECT 2296.330 141.690 2297.510 142.870 ;
        RECT 2297.930 141.690 2299.110 142.870 ;
        RECT 2296.330 -26.910 2297.510 -25.730 ;
        RECT 2297.930 -26.910 2299.110 -25.730 ;
        RECT 2296.330 -28.510 2297.510 -27.330 ;
        RECT 2297.930 -28.510 2299.110 -27.330 ;
        RECT 2476.330 3547.010 2477.510 3548.190 ;
        RECT 2477.930 3547.010 2479.110 3548.190 ;
        RECT 2476.330 3545.410 2477.510 3546.590 ;
        RECT 2477.930 3545.410 2479.110 3546.590 ;
        RECT 2476.330 3383.290 2477.510 3384.470 ;
        RECT 2477.930 3383.290 2479.110 3384.470 ;
        RECT 2476.330 3381.690 2477.510 3382.870 ;
        RECT 2477.930 3381.690 2479.110 3382.870 ;
        RECT 2476.330 3203.290 2477.510 3204.470 ;
        RECT 2477.930 3203.290 2479.110 3204.470 ;
        RECT 2476.330 3201.690 2477.510 3202.870 ;
        RECT 2477.930 3201.690 2479.110 3202.870 ;
        RECT 2476.330 3023.290 2477.510 3024.470 ;
        RECT 2477.930 3023.290 2479.110 3024.470 ;
        RECT 2476.330 3021.690 2477.510 3022.870 ;
        RECT 2477.930 3021.690 2479.110 3022.870 ;
        RECT 2476.330 2843.290 2477.510 2844.470 ;
        RECT 2477.930 2843.290 2479.110 2844.470 ;
        RECT 2476.330 2841.690 2477.510 2842.870 ;
        RECT 2477.930 2841.690 2479.110 2842.870 ;
        RECT 2476.330 2663.290 2477.510 2664.470 ;
        RECT 2477.930 2663.290 2479.110 2664.470 ;
        RECT 2476.330 2661.690 2477.510 2662.870 ;
        RECT 2477.930 2661.690 2479.110 2662.870 ;
        RECT 2476.330 2483.290 2477.510 2484.470 ;
        RECT 2477.930 2483.290 2479.110 2484.470 ;
        RECT 2476.330 2481.690 2477.510 2482.870 ;
        RECT 2477.930 2481.690 2479.110 2482.870 ;
        RECT 2476.330 2303.290 2477.510 2304.470 ;
        RECT 2477.930 2303.290 2479.110 2304.470 ;
        RECT 2476.330 2301.690 2477.510 2302.870 ;
        RECT 2477.930 2301.690 2479.110 2302.870 ;
        RECT 2476.330 2123.290 2477.510 2124.470 ;
        RECT 2477.930 2123.290 2479.110 2124.470 ;
        RECT 2476.330 2121.690 2477.510 2122.870 ;
        RECT 2477.930 2121.690 2479.110 2122.870 ;
        RECT 2476.330 1943.290 2477.510 1944.470 ;
        RECT 2477.930 1943.290 2479.110 1944.470 ;
        RECT 2476.330 1941.690 2477.510 1942.870 ;
        RECT 2477.930 1941.690 2479.110 1942.870 ;
        RECT 2476.330 1763.290 2477.510 1764.470 ;
        RECT 2477.930 1763.290 2479.110 1764.470 ;
        RECT 2476.330 1761.690 2477.510 1762.870 ;
        RECT 2477.930 1761.690 2479.110 1762.870 ;
        RECT 2476.330 1583.290 2477.510 1584.470 ;
        RECT 2477.930 1583.290 2479.110 1584.470 ;
        RECT 2476.330 1581.690 2477.510 1582.870 ;
        RECT 2477.930 1581.690 2479.110 1582.870 ;
        RECT 2476.330 1403.290 2477.510 1404.470 ;
        RECT 2477.930 1403.290 2479.110 1404.470 ;
        RECT 2476.330 1401.690 2477.510 1402.870 ;
        RECT 2477.930 1401.690 2479.110 1402.870 ;
        RECT 2476.330 1223.290 2477.510 1224.470 ;
        RECT 2477.930 1223.290 2479.110 1224.470 ;
        RECT 2476.330 1221.690 2477.510 1222.870 ;
        RECT 2477.930 1221.690 2479.110 1222.870 ;
        RECT 2476.330 1043.290 2477.510 1044.470 ;
        RECT 2477.930 1043.290 2479.110 1044.470 ;
        RECT 2476.330 1041.690 2477.510 1042.870 ;
        RECT 2477.930 1041.690 2479.110 1042.870 ;
        RECT 2476.330 863.290 2477.510 864.470 ;
        RECT 2477.930 863.290 2479.110 864.470 ;
        RECT 2476.330 861.690 2477.510 862.870 ;
        RECT 2477.930 861.690 2479.110 862.870 ;
        RECT 2476.330 683.290 2477.510 684.470 ;
        RECT 2477.930 683.290 2479.110 684.470 ;
        RECT 2476.330 681.690 2477.510 682.870 ;
        RECT 2477.930 681.690 2479.110 682.870 ;
        RECT 2476.330 503.290 2477.510 504.470 ;
        RECT 2477.930 503.290 2479.110 504.470 ;
        RECT 2476.330 501.690 2477.510 502.870 ;
        RECT 2477.930 501.690 2479.110 502.870 ;
        RECT 2476.330 323.290 2477.510 324.470 ;
        RECT 2477.930 323.290 2479.110 324.470 ;
        RECT 2476.330 321.690 2477.510 322.870 ;
        RECT 2477.930 321.690 2479.110 322.870 ;
        RECT 2476.330 143.290 2477.510 144.470 ;
        RECT 2477.930 143.290 2479.110 144.470 ;
        RECT 2476.330 141.690 2477.510 142.870 ;
        RECT 2477.930 141.690 2479.110 142.870 ;
        RECT 2476.330 -26.910 2477.510 -25.730 ;
        RECT 2477.930 -26.910 2479.110 -25.730 ;
        RECT 2476.330 -28.510 2477.510 -27.330 ;
        RECT 2477.930 -28.510 2479.110 -27.330 ;
        RECT 2656.330 3547.010 2657.510 3548.190 ;
        RECT 2657.930 3547.010 2659.110 3548.190 ;
        RECT 2656.330 3545.410 2657.510 3546.590 ;
        RECT 2657.930 3545.410 2659.110 3546.590 ;
        RECT 2656.330 3383.290 2657.510 3384.470 ;
        RECT 2657.930 3383.290 2659.110 3384.470 ;
        RECT 2656.330 3381.690 2657.510 3382.870 ;
        RECT 2657.930 3381.690 2659.110 3382.870 ;
        RECT 2656.330 3203.290 2657.510 3204.470 ;
        RECT 2657.930 3203.290 2659.110 3204.470 ;
        RECT 2656.330 3201.690 2657.510 3202.870 ;
        RECT 2657.930 3201.690 2659.110 3202.870 ;
        RECT 2656.330 3023.290 2657.510 3024.470 ;
        RECT 2657.930 3023.290 2659.110 3024.470 ;
        RECT 2656.330 3021.690 2657.510 3022.870 ;
        RECT 2657.930 3021.690 2659.110 3022.870 ;
        RECT 2656.330 2843.290 2657.510 2844.470 ;
        RECT 2657.930 2843.290 2659.110 2844.470 ;
        RECT 2656.330 2841.690 2657.510 2842.870 ;
        RECT 2657.930 2841.690 2659.110 2842.870 ;
        RECT 2656.330 2663.290 2657.510 2664.470 ;
        RECT 2657.930 2663.290 2659.110 2664.470 ;
        RECT 2656.330 2661.690 2657.510 2662.870 ;
        RECT 2657.930 2661.690 2659.110 2662.870 ;
        RECT 2656.330 2483.290 2657.510 2484.470 ;
        RECT 2657.930 2483.290 2659.110 2484.470 ;
        RECT 2656.330 2481.690 2657.510 2482.870 ;
        RECT 2657.930 2481.690 2659.110 2482.870 ;
        RECT 2656.330 2303.290 2657.510 2304.470 ;
        RECT 2657.930 2303.290 2659.110 2304.470 ;
        RECT 2656.330 2301.690 2657.510 2302.870 ;
        RECT 2657.930 2301.690 2659.110 2302.870 ;
        RECT 2656.330 2123.290 2657.510 2124.470 ;
        RECT 2657.930 2123.290 2659.110 2124.470 ;
        RECT 2656.330 2121.690 2657.510 2122.870 ;
        RECT 2657.930 2121.690 2659.110 2122.870 ;
        RECT 2656.330 1943.290 2657.510 1944.470 ;
        RECT 2657.930 1943.290 2659.110 1944.470 ;
        RECT 2656.330 1941.690 2657.510 1942.870 ;
        RECT 2657.930 1941.690 2659.110 1942.870 ;
        RECT 2656.330 1763.290 2657.510 1764.470 ;
        RECT 2657.930 1763.290 2659.110 1764.470 ;
        RECT 2656.330 1761.690 2657.510 1762.870 ;
        RECT 2657.930 1761.690 2659.110 1762.870 ;
        RECT 2656.330 1583.290 2657.510 1584.470 ;
        RECT 2657.930 1583.290 2659.110 1584.470 ;
        RECT 2656.330 1581.690 2657.510 1582.870 ;
        RECT 2657.930 1581.690 2659.110 1582.870 ;
        RECT 2656.330 1403.290 2657.510 1404.470 ;
        RECT 2657.930 1403.290 2659.110 1404.470 ;
        RECT 2656.330 1401.690 2657.510 1402.870 ;
        RECT 2657.930 1401.690 2659.110 1402.870 ;
        RECT 2656.330 1223.290 2657.510 1224.470 ;
        RECT 2657.930 1223.290 2659.110 1224.470 ;
        RECT 2656.330 1221.690 2657.510 1222.870 ;
        RECT 2657.930 1221.690 2659.110 1222.870 ;
        RECT 2656.330 1043.290 2657.510 1044.470 ;
        RECT 2657.930 1043.290 2659.110 1044.470 ;
        RECT 2656.330 1041.690 2657.510 1042.870 ;
        RECT 2657.930 1041.690 2659.110 1042.870 ;
        RECT 2656.330 863.290 2657.510 864.470 ;
        RECT 2657.930 863.290 2659.110 864.470 ;
        RECT 2656.330 861.690 2657.510 862.870 ;
        RECT 2657.930 861.690 2659.110 862.870 ;
        RECT 2656.330 683.290 2657.510 684.470 ;
        RECT 2657.930 683.290 2659.110 684.470 ;
        RECT 2656.330 681.690 2657.510 682.870 ;
        RECT 2657.930 681.690 2659.110 682.870 ;
        RECT 2656.330 503.290 2657.510 504.470 ;
        RECT 2657.930 503.290 2659.110 504.470 ;
        RECT 2656.330 501.690 2657.510 502.870 ;
        RECT 2657.930 501.690 2659.110 502.870 ;
        RECT 2656.330 323.290 2657.510 324.470 ;
        RECT 2657.930 323.290 2659.110 324.470 ;
        RECT 2656.330 321.690 2657.510 322.870 ;
        RECT 2657.930 321.690 2659.110 322.870 ;
        RECT 2656.330 143.290 2657.510 144.470 ;
        RECT 2657.930 143.290 2659.110 144.470 ;
        RECT 2656.330 141.690 2657.510 142.870 ;
        RECT 2657.930 141.690 2659.110 142.870 ;
        RECT 2656.330 -26.910 2657.510 -25.730 ;
        RECT 2657.930 -26.910 2659.110 -25.730 ;
        RECT 2656.330 -28.510 2657.510 -27.330 ;
        RECT 2657.930 -28.510 2659.110 -27.330 ;
        RECT 2836.330 3547.010 2837.510 3548.190 ;
        RECT 2837.930 3547.010 2839.110 3548.190 ;
        RECT 2836.330 3545.410 2837.510 3546.590 ;
        RECT 2837.930 3545.410 2839.110 3546.590 ;
        RECT 2836.330 3383.290 2837.510 3384.470 ;
        RECT 2837.930 3383.290 2839.110 3384.470 ;
        RECT 2836.330 3381.690 2837.510 3382.870 ;
        RECT 2837.930 3381.690 2839.110 3382.870 ;
        RECT 2836.330 3203.290 2837.510 3204.470 ;
        RECT 2837.930 3203.290 2839.110 3204.470 ;
        RECT 2836.330 3201.690 2837.510 3202.870 ;
        RECT 2837.930 3201.690 2839.110 3202.870 ;
        RECT 2836.330 3023.290 2837.510 3024.470 ;
        RECT 2837.930 3023.290 2839.110 3024.470 ;
        RECT 2836.330 3021.690 2837.510 3022.870 ;
        RECT 2837.930 3021.690 2839.110 3022.870 ;
        RECT 2836.330 2843.290 2837.510 2844.470 ;
        RECT 2837.930 2843.290 2839.110 2844.470 ;
        RECT 2836.330 2841.690 2837.510 2842.870 ;
        RECT 2837.930 2841.690 2839.110 2842.870 ;
        RECT 2836.330 2663.290 2837.510 2664.470 ;
        RECT 2837.930 2663.290 2839.110 2664.470 ;
        RECT 2836.330 2661.690 2837.510 2662.870 ;
        RECT 2837.930 2661.690 2839.110 2662.870 ;
        RECT 2836.330 2483.290 2837.510 2484.470 ;
        RECT 2837.930 2483.290 2839.110 2484.470 ;
        RECT 2836.330 2481.690 2837.510 2482.870 ;
        RECT 2837.930 2481.690 2839.110 2482.870 ;
        RECT 2836.330 2303.290 2837.510 2304.470 ;
        RECT 2837.930 2303.290 2839.110 2304.470 ;
        RECT 2836.330 2301.690 2837.510 2302.870 ;
        RECT 2837.930 2301.690 2839.110 2302.870 ;
        RECT 2836.330 2123.290 2837.510 2124.470 ;
        RECT 2837.930 2123.290 2839.110 2124.470 ;
        RECT 2836.330 2121.690 2837.510 2122.870 ;
        RECT 2837.930 2121.690 2839.110 2122.870 ;
        RECT 2836.330 1943.290 2837.510 1944.470 ;
        RECT 2837.930 1943.290 2839.110 1944.470 ;
        RECT 2836.330 1941.690 2837.510 1942.870 ;
        RECT 2837.930 1941.690 2839.110 1942.870 ;
        RECT 2836.330 1763.290 2837.510 1764.470 ;
        RECT 2837.930 1763.290 2839.110 1764.470 ;
        RECT 2836.330 1761.690 2837.510 1762.870 ;
        RECT 2837.930 1761.690 2839.110 1762.870 ;
        RECT 2836.330 1583.290 2837.510 1584.470 ;
        RECT 2837.930 1583.290 2839.110 1584.470 ;
        RECT 2836.330 1581.690 2837.510 1582.870 ;
        RECT 2837.930 1581.690 2839.110 1582.870 ;
        RECT 2836.330 1403.290 2837.510 1404.470 ;
        RECT 2837.930 1403.290 2839.110 1404.470 ;
        RECT 2836.330 1401.690 2837.510 1402.870 ;
        RECT 2837.930 1401.690 2839.110 1402.870 ;
        RECT 2836.330 1223.290 2837.510 1224.470 ;
        RECT 2837.930 1223.290 2839.110 1224.470 ;
        RECT 2836.330 1221.690 2837.510 1222.870 ;
        RECT 2837.930 1221.690 2839.110 1222.870 ;
        RECT 2836.330 1043.290 2837.510 1044.470 ;
        RECT 2837.930 1043.290 2839.110 1044.470 ;
        RECT 2836.330 1041.690 2837.510 1042.870 ;
        RECT 2837.930 1041.690 2839.110 1042.870 ;
        RECT 2836.330 863.290 2837.510 864.470 ;
        RECT 2837.930 863.290 2839.110 864.470 ;
        RECT 2836.330 861.690 2837.510 862.870 ;
        RECT 2837.930 861.690 2839.110 862.870 ;
        RECT 2836.330 683.290 2837.510 684.470 ;
        RECT 2837.930 683.290 2839.110 684.470 ;
        RECT 2836.330 681.690 2837.510 682.870 ;
        RECT 2837.930 681.690 2839.110 682.870 ;
        RECT 2836.330 503.290 2837.510 504.470 ;
        RECT 2837.930 503.290 2839.110 504.470 ;
        RECT 2836.330 501.690 2837.510 502.870 ;
        RECT 2837.930 501.690 2839.110 502.870 ;
        RECT 2836.330 323.290 2837.510 324.470 ;
        RECT 2837.930 323.290 2839.110 324.470 ;
        RECT 2836.330 321.690 2837.510 322.870 ;
        RECT 2837.930 321.690 2839.110 322.870 ;
        RECT 2836.330 143.290 2837.510 144.470 ;
        RECT 2837.930 143.290 2839.110 144.470 ;
        RECT 2836.330 141.690 2837.510 142.870 ;
        RECT 2837.930 141.690 2839.110 142.870 ;
        RECT 2836.330 -26.910 2837.510 -25.730 ;
        RECT 2837.930 -26.910 2839.110 -25.730 ;
        RECT 2836.330 -28.510 2837.510 -27.330 ;
        RECT 2837.930 -28.510 2839.110 -27.330 ;
        RECT 2950.710 3547.010 2951.890 3548.190 ;
        RECT 2952.310 3547.010 2953.490 3548.190 ;
        RECT 2950.710 3545.410 2951.890 3546.590 ;
        RECT 2952.310 3545.410 2953.490 3546.590 ;
        RECT 2950.710 3383.290 2951.890 3384.470 ;
        RECT 2952.310 3383.290 2953.490 3384.470 ;
        RECT 2950.710 3381.690 2951.890 3382.870 ;
        RECT 2952.310 3381.690 2953.490 3382.870 ;
        RECT 2950.710 3203.290 2951.890 3204.470 ;
        RECT 2952.310 3203.290 2953.490 3204.470 ;
        RECT 2950.710 3201.690 2951.890 3202.870 ;
        RECT 2952.310 3201.690 2953.490 3202.870 ;
        RECT 2950.710 3023.290 2951.890 3024.470 ;
        RECT 2952.310 3023.290 2953.490 3024.470 ;
        RECT 2950.710 3021.690 2951.890 3022.870 ;
        RECT 2952.310 3021.690 2953.490 3022.870 ;
        RECT 2950.710 2843.290 2951.890 2844.470 ;
        RECT 2952.310 2843.290 2953.490 2844.470 ;
        RECT 2950.710 2841.690 2951.890 2842.870 ;
        RECT 2952.310 2841.690 2953.490 2842.870 ;
        RECT 2950.710 2663.290 2951.890 2664.470 ;
        RECT 2952.310 2663.290 2953.490 2664.470 ;
        RECT 2950.710 2661.690 2951.890 2662.870 ;
        RECT 2952.310 2661.690 2953.490 2662.870 ;
        RECT 2950.710 2483.290 2951.890 2484.470 ;
        RECT 2952.310 2483.290 2953.490 2484.470 ;
        RECT 2950.710 2481.690 2951.890 2482.870 ;
        RECT 2952.310 2481.690 2953.490 2482.870 ;
        RECT 2950.710 2303.290 2951.890 2304.470 ;
        RECT 2952.310 2303.290 2953.490 2304.470 ;
        RECT 2950.710 2301.690 2951.890 2302.870 ;
        RECT 2952.310 2301.690 2953.490 2302.870 ;
        RECT 2950.710 2123.290 2951.890 2124.470 ;
        RECT 2952.310 2123.290 2953.490 2124.470 ;
        RECT 2950.710 2121.690 2951.890 2122.870 ;
        RECT 2952.310 2121.690 2953.490 2122.870 ;
        RECT 2950.710 1943.290 2951.890 1944.470 ;
        RECT 2952.310 1943.290 2953.490 1944.470 ;
        RECT 2950.710 1941.690 2951.890 1942.870 ;
        RECT 2952.310 1941.690 2953.490 1942.870 ;
        RECT 2950.710 1763.290 2951.890 1764.470 ;
        RECT 2952.310 1763.290 2953.490 1764.470 ;
        RECT 2950.710 1761.690 2951.890 1762.870 ;
        RECT 2952.310 1761.690 2953.490 1762.870 ;
        RECT 2950.710 1583.290 2951.890 1584.470 ;
        RECT 2952.310 1583.290 2953.490 1584.470 ;
        RECT 2950.710 1581.690 2951.890 1582.870 ;
        RECT 2952.310 1581.690 2953.490 1582.870 ;
        RECT 2950.710 1403.290 2951.890 1404.470 ;
        RECT 2952.310 1403.290 2953.490 1404.470 ;
        RECT 2950.710 1401.690 2951.890 1402.870 ;
        RECT 2952.310 1401.690 2953.490 1402.870 ;
        RECT 2950.710 1223.290 2951.890 1224.470 ;
        RECT 2952.310 1223.290 2953.490 1224.470 ;
        RECT 2950.710 1221.690 2951.890 1222.870 ;
        RECT 2952.310 1221.690 2953.490 1222.870 ;
        RECT 2950.710 1043.290 2951.890 1044.470 ;
        RECT 2952.310 1043.290 2953.490 1044.470 ;
        RECT 2950.710 1041.690 2951.890 1042.870 ;
        RECT 2952.310 1041.690 2953.490 1042.870 ;
        RECT 2950.710 863.290 2951.890 864.470 ;
        RECT 2952.310 863.290 2953.490 864.470 ;
        RECT 2950.710 861.690 2951.890 862.870 ;
        RECT 2952.310 861.690 2953.490 862.870 ;
        RECT 2950.710 683.290 2951.890 684.470 ;
        RECT 2952.310 683.290 2953.490 684.470 ;
        RECT 2950.710 681.690 2951.890 682.870 ;
        RECT 2952.310 681.690 2953.490 682.870 ;
        RECT 2950.710 503.290 2951.890 504.470 ;
        RECT 2952.310 503.290 2953.490 504.470 ;
        RECT 2950.710 501.690 2951.890 502.870 ;
        RECT 2952.310 501.690 2953.490 502.870 ;
        RECT 2950.710 323.290 2951.890 324.470 ;
        RECT 2952.310 323.290 2953.490 324.470 ;
        RECT 2950.710 321.690 2951.890 322.870 ;
        RECT 2952.310 321.690 2953.490 322.870 ;
        RECT 2950.710 143.290 2951.890 144.470 ;
        RECT 2952.310 143.290 2953.490 144.470 ;
        RECT 2950.710 141.690 2951.890 142.870 ;
        RECT 2952.310 141.690 2953.490 142.870 ;
        RECT 2950.710 -26.910 2951.890 -25.730 ;
        RECT 2952.310 -26.910 2953.490 -25.730 ;
        RECT 2950.710 -28.510 2951.890 -27.330 ;
        RECT 2952.310 -28.510 2953.490 -27.330 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
        RECT -34.030 861.530 2953.650 864.630 ;
        RECT -34.030 681.530 2953.650 684.630 ;
        RECT -34.030 501.530 2953.650 504.630 ;
        RECT -34.030 321.530 2953.650 324.630 ;
        RECT -34.030 141.530 2953.650 144.630 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
        RECT 334.770 1010.000 337.870 3557.950 ;
        RECT 514.770 1010.000 517.870 3557.950 ;
        RECT 694.770 1010.000 697.870 3557.950 ;
        RECT 874.770 1010.000 877.870 3557.950 ;
        RECT 1054.770 1010.000 1057.870 3557.950 ;
        RECT 334.770 -38.270 337.870 390.000 ;
        RECT 514.770 -38.270 517.870 390.000 ;
        RECT 694.770 -38.270 697.870 390.000 ;
        RECT 874.770 -38.270 877.870 390.000 ;
        RECT 1054.770 -38.270 1057.870 390.000 ;
        RECT 1234.770 -38.270 1237.870 3557.950 ;
        RECT 1414.770 -38.270 1417.870 3557.950 ;
        RECT 1594.770 -38.270 1597.870 3557.950 ;
        RECT 1774.770 -38.270 1777.870 3557.950 ;
        RECT 1954.770 -38.270 1957.870 3557.950 ;
        RECT 2134.770 -38.270 2137.870 3557.950 ;
        RECT 2314.770 -38.270 2317.870 3557.950 ;
        RECT 2494.770 -38.270 2497.870 3557.950 ;
        RECT 2674.770 -38.270 2677.870 3557.950 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER via4 ;
        RECT -43.470 3556.610 -42.290 3557.790 ;
        RECT -41.870 3556.610 -40.690 3557.790 ;
        RECT -43.470 3555.010 -42.290 3556.190 ;
        RECT -41.870 3555.010 -40.690 3556.190 ;
        RECT -43.470 3401.890 -42.290 3403.070 ;
        RECT -41.870 3401.890 -40.690 3403.070 ;
        RECT -43.470 3400.290 -42.290 3401.470 ;
        RECT -41.870 3400.290 -40.690 3401.470 ;
        RECT -43.470 3221.890 -42.290 3223.070 ;
        RECT -41.870 3221.890 -40.690 3223.070 ;
        RECT -43.470 3220.290 -42.290 3221.470 ;
        RECT -41.870 3220.290 -40.690 3221.470 ;
        RECT -43.470 3041.890 -42.290 3043.070 ;
        RECT -41.870 3041.890 -40.690 3043.070 ;
        RECT -43.470 3040.290 -42.290 3041.470 ;
        RECT -41.870 3040.290 -40.690 3041.470 ;
        RECT -43.470 2861.890 -42.290 2863.070 ;
        RECT -41.870 2861.890 -40.690 2863.070 ;
        RECT -43.470 2860.290 -42.290 2861.470 ;
        RECT -41.870 2860.290 -40.690 2861.470 ;
        RECT -43.470 2681.890 -42.290 2683.070 ;
        RECT -41.870 2681.890 -40.690 2683.070 ;
        RECT -43.470 2680.290 -42.290 2681.470 ;
        RECT -41.870 2680.290 -40.690 2681.470 ;
        RECT -43.470 2501.890 -42.290 2503.070 ;
        RECT -41.870 2501.890 -40.690 2503.070 ;
        RECT -43.470 2500.290 -42.290 2501.470 ;
        RECT -41.870 2500.290 -40.690 2501.470 ;
        RECT -43.470 2321.890 -42.290 2323.070 ;
        RECT -41.870 2321.890 -40.690 2323.070 ;
        RECT -43.470 2320.290 -42.290 2321.470 ;
        RECT -41.870 2320.290 -40.690 2321.470 ;
        RECT -43.470 2141.890 -42.290 2143.070 ;
        RECT -41.870 2141.890 -40.690 2143.070 ;
        RECT -43.470 2140.290 -42.290 2141.470 ;
        RECT -41.870 2140.290 -40.690 2141.470 ;
        RECT -43.470 1961.890 -42.290 1963.070 ;
        RECT -41.870 1961.890 -40.690 1963.070 ;
        RECT -43.470 1960.290 -42.290 1961.470 ;
        RECT -41.870 1960.290 -40.690 1961.470 ;
        RECT -43.470 1781.890 -42.290 1783.070 ;
        RECT -41.870 1781.890 -40.690 1783.070 ;
        RECT -43.470 1780.290 -42.290 1781.470 ;
        RECT -41.870 1780.290 -40.690 1781.470 ;
        RECT -43.470 1601.890 -42.290 1603.070 ;
        RECT -41.870 1601.890 -40.690 1603.070 ;
        RECT -43.470 1600.290 -42.290 1601.470 ;
        RECT -41.870 1600.290 -40.690 1601.470 ;
        RECT -43.470 1421.890 -42.290 1423.070 ;
        RECT -41.870 1421.890 -40.690 1423.070 ;
        RECT -43.470 1420.290 -42.290 1421.470 ;
        RECT -41.870 1420.290 -40.690 1421.470 ;
        RECT -43.470 1241.890 -42.290 1243.070 ;
        RECT -41.870 1241.890 -40.690 1243.070 ;
        RECT -43.470 1240.290 -42.290 1241.470 ;
        RECT -41.870 1240.290 -40.690 1241.470 ;
        RECT -43.470 1061.890 -42.290 1063.070 ;
        RECT -41.870 1061.890 -40.690 1063.070 ;
        RECT -43.470 1060.290 -42.290 1061.470 ;
        RECT -41.870 1060.290 -40.690 1061.470 ;
        RECT -43.470 881.890 -42.290 883.070 ;
        RECT -41.870 881.890 -40.690 883.070 ;
        RECT -43.470 880.290 -42.290 881.470 ;
        RECT -41.870 880.290 -40.690 881.470 ;
        RECT -43.470 701.890 -42.290 703.070 ;
        RECT -41.870 701.890 -40.690 703.070 ;
        RECT -43.470 700.290 -42.290 701.470 ;
        RECT -41.870 700.290 -40.690 701.470 ;
        RECT -43.470 521.890 -42.290 523.070 ;
        RECT -41.870 521.890 -40.690 523.070 ;
        RECT -43.470 520.290 -42.290 521.470 ;
        RECT -41.870 520.290 -40.690 521.470 ;
        RECT -43.470 341.890 -42.290 343.070 ;
        RECT -41.870 341.890 -40.690 343.070 ;
        RECT -43.470 340.290 -42.290 341.470 ;
        RECT -41.870 340.290 -40.690 341.470 ;
        RECT -43.470 161.890 -42.290 163.070 ;
        RECT -41.870 161.890 -40.690 163.070 ;
        RECT -43.470 160.290 -42.290 161.470 ;
        RECT -41.870 160.290 -40.690 161.470 ;
        RECT -43.470 -36.510 -42.290 -35.330 ;
        RECT -41.870 -36.510 -40.690 -35.330 ;
        RECT -43.470 -38.110 -42.290 -36.930 ;
        RECT -41.870 -38.110 -40.690 -36.930 ;
        RECT 154.930 3556.610 156.110 3557.790 ;
        RECT 156.530 3556.610 157.710 3557.790 ;
        RECT 154.930 3555.010 156.110 3556.190 ;
        RECT 156.530 3555.010 157.710 3556.190 ;
        RECT 154.930 3401.890 156.110 3403.070 ;
        RECT 156.530 3401.890 157.710 3403.070 ;
        RECT 154.930 3400.290 156.110 3401.470 ;
        RECT 156.530 3400.290 157.710 3401.470 ;
        RECT 154.930 3221.890 156.110 3223.070 ;
        RECT 156.530 3221.890 157.710 3223.070 ;
        RECT 154.930 3220.290 156.110 3221.470 ;
        RECT 156.530 3220.290 157.710 3221.470 ;
        RECT 154.930 3041.890 156.110 3043.070 ;
        RECT 156.530 3041.890 157.710 3043.070 ;
        RECT 154.930 3040.290 156.110 3041.470 ;
        RECT 156.530 3040.290 157.710 3041.470 ;
        RECT 154.930 2861.890 156.110 2863.070 ;
        RECT 156.530 2861.890 157.710 2863.070 ;
        RECT 154.930 2860.290 156.110 2861.470 ;
        RECT 156.530 2860.290 157.710 2861.470 ;
        RECT 154.930 2681.890 156.110 2683.070 ;
        RECT 156.530 2681.890 157.710 2683.070 ;
        RECT 154.930 2680.290 156.110 2681.470 ;
        RECT 156.530 2680.290 157.710 2681.470 ;
        RECT 154.930 2501.890 156.110 2503.070 ;
        RECT 156.530 2501.890 157.710 2503.070 ;
        RECT 154.930 2500.290 156.110 2501.470 ;
        RECT 156.530 2500.290 157.710 2501.470 ;
        RECT 154.930 2321.890 156.110 2323.070 ;
        RECT 156.530 2321.890 157.710 2323.070 ;
        RECT 154.930 2320.290 156.110 2321.470 ;
        RECT 156.530 2320.290 157.710 2321.470 ;
        RECT 154.930 2141.890 156.110 2143.070 ;
        RECT 156.530 2141.890 157.710 2143.070 ;
        RECT 154.930 2140.290 156.110 2141.470 ;
        RECT 156.530 2140.290 157.710 2141.470 ;
        RECT 154.930 1961.890 156.110 1963.070 ;
        RECT 156.530 1961.890 157.710 1963.070 ;
        RECT 154.930 1960.290 156.110 1961.470 ;
        RECT 156.530 1960.290 157.710 1961.470 ;
        RECT 154.930 1781.890 156.110 1783.070 ;
        RECT 156.530 1781.890 157.710 1783.070 ;
        RECT 154.930 1780.290 156.110 1781.470 ;
        RECT 156.530 1780.290 157.710 1781.470 ;
        RECT 154.930 1601.890 156.110 1603.070 ;
        RECT 156.530 1601.890 157.710 1603.070 ;
        RECT 154.930 1600.290 156.110 1601.470 ;
        RECT 156.530 1600.290 157.710 1601.470 ;
        RECT 154.930 1421.890 156.110 1423.070 ;
        RECT 156.530 1421.890 157.710 1423.070 ;
        RECT 154.930 1420.290 156.110 1421.470 ;
        RECT 156.530 1420.290 157.710 1421.470 ;
        RECT 154.930 1241.890 156.110 1243.070 ;
        RECT 156.530 1241.890 157.710 1243.070 ;
        RECT 154.930 1240.290 156.110 1241.470 ;
        RECT 156.530 1240.290 157.710 1241.470 ;
        RECT 154.930 1061.890 156.110 1063.070 ;
        RECT 156.530 1061.890 157.710 1063.070 ;
        RECT 154.930 1060.290 156.110 1061.470 ;
        RECT 156.530 1060.290 157.710 1061.470 ;
        RECT 334.930 3556.610 336.110 3557.790 ;
        RECT 336.530 3556.610 337.710 3557.790 ;
        RECT 334.930 3555.010 336.110 3556.190 ;
        RECT 336.530 3555.010 337.710 3556.190 ;
        RECT 334.930 3401.890 336.110 3403.070 ;
        RECT 336.530 3401.890 337.710 3403.070 ;
        RECT 334.930 3400.290 336.110 3401.470 ;
        RECT 336.530 3400.290 337.710 3401.470 ;
        RECT 334.930 3221.890 336.110 3223.070 ;
        RECT 336.530 3221.890 337.710 3223.070 ;
        RECT 334.930 3220.290 336.110 3221.470 ;
        RECT 336.530 3220.290 337.710 3221.470 ;
        RECT 334.930 3041.890 336.110 3043.070 ;
        RECT 336.530 3041.890 337.710 3043.070 ;
        RECT 334.930 3040.290 336.110 3041.470 ;
        RECT 336.530 3040.290 337.710 3041.470 ;
        RECT 334.930 2861.890 336.110 2863.070 ;
        RECT 336.530 2861.890 337.710 2863.070 ;
        RECT 334.930 2860.290 336.110 2861.470 ;
        RECT 336.530 2860.290 337.710 2861.470 ;
        RECT 334.930 2681.890 336.110 2683.070 ;
        RECT 336.530 2681.890 337.710 2683.070 ;
        RECT 334.930 2680.290 336.110 2681.470 ;
        RECT 336.530 2680.290 337.710 2681.470 ;
        RECT 334.930 2501.890 336.110 2503.070 ;
        RECT 336.530 2501.890 337.710 2503.070 ;
        RECT 334.930 2500.290 336.110 2501.470 ;
        RECT 336.530 2500.290 337.710 2501.470 ;
        RECT 334.930 2321.890 336.110 2323.070 ;
        RECT 336.530 2321.890 337.710 2323.070 ;
        RECT 334.930 2320.290 336.110 2321.470 ;
        RECT 336.530 2320.290 337.710 2321.470 ;
        RECT 334.930 2141.890 336.110 2143.070 ;
        RECT 336.530 2141.890 337.710 2143.070 ;
        RECT 334.930 2140.290 336.110 2141.470 ;
        RECT 336.530 2140.290 337.710 2141.470 ;
        RECT 334.930 1961.890 336.110 1963.070 ;
        RECT 336.530 1961.890 337.710 1963.070 ;
        RECT 334.930 1960.290 336.110 1961.470 ;
        RECT 336.530 1960.290 337.710 1961.470 ;
        RECT 334.930 1781.890 336.110 1783.070 ;
        RECT 336.530 1781.890 337.710 1783.070 ;
        RECT 334.930 1780.290 336.110 1781.470 ;
        RECT 336.530 1780.290 337.710 1781.470 ;
        RECT 334.930 1601.890 336.110 1603.070 ;
        RECT 336.530 1601.890 337.710 1603.070 ;
        RECT 334.930 1600.290 336.110 1601.470 ;
        RECT 336.530 1600.290 337.710 1601.470 ;
        RECT 334.930 1421.890 336.110 1423.070 ;
        RECT 336.530 1421.890 337.710 1423.070 ;
        RECT 334.930 1420.290 336.110 1421.470 ;
        RECT 336.530 1420.290 337.710 1421.470 ;
        RECT 334.930 1241.890 336.110 1243.070 ;
        RECT 336.530 1241.890 337.710 1243.070 ;
        RECT 334.930 1240.290 336.110 1241.470 ;
        RECT 336.530 1240.290 337.710 1241.470 ;
        RECT 334.930 1061.890 336.110 1063.070 ;
        RECT 336.530 1061.890 337.710 1063.070 ;
        RECT 334.930 1060.290 336.110 1061.470 ;
        RECT 336.530 1060.290 337.710 1061.470 ;
        RECT 514.930 3556.610 516.110 3557.790 ;
        RECT 516.530 3556.610 517.710 3557.790 ;
        RECT 514.930 3555.010 516.110 3556.190 ;
        RECT 516.530 3555.010 517.710 3556.190 ;
        RECT 514.930 3401.890 516.110 3403.070 ;
        RECT 516.530 3401.890 517.710 3403.070 ;
        RECT 514.930 3400.290 516.110 3401.470 ;
        RECT 516.530 3400.290 517.710 3401.470 ;
        RECT 514.930 3221.890 516.110 3223.070 ;
        RECT 516.530 3221.890 517.710 3223.070 ;
        RECT 514.930 3220.290 516.110 3221.470 ;
        RECT 516.530 3220.290 517.710 3221.470 ;
        RECT 514.930 3041.890 516.110 3043.070 ;
        RECT 516.530 3041.890 517.710 3043.070 ;
        RECT 514.930 3040.290 516.110 3041.470 ;
        RECT 516.530 3040.290 517.710 3041.470 ;
        RECT 514.930 2861.890 516.110 2863.070 ;
        RECT 516.530 2861.890 517.710 2863.070 ;
        RECT 514.930 2860.290 516.110 2861.470 ;
        RECT 516.530 2860.290 517.710 2861.470 ;
        RECT 514.930 2681.890 516.110 2683.070 ;
        RECT 516.530 2681.890 517.710 2683.070 ;
        RECT 514.930 2680.290 516.110 2681.470 ;
        RECT 516.530 2680.290 517.710 2681.470 ;
        RECT 514.930 2501.890 516.110 2503.070 ;
        RECT 516.530 2501.890 517.710 2503.070 ;
        RECT 514.930 2500.290 516.110 2501.470 ;
        RECT 516.530 2500.290 517.710 2501.470 ;
        RECT 514.930 2321.890 516.110 2323.070 ;
        RECT 516.530 2321.890 517.710 2323.070 ;
        RECT 514.930 2320.290 516.110 2321.470 ;
        RECT 516.530 2320.290 517.710 2321.470 ;
        RECT 514.930 2141.890 516.110 2143.070 ;
        RECT 516.530 2141.890 517.710 2143.070 ;
        RECT 514.930 2140.290 516.110 2141.470 ;
        RECT 516.530 2140.290 517.710 2141.470 ;
        RECT 514.930 1961.890 516.110 1963.070 ;
        RECT 516.530 1961.890 517.710 1963.070 ;
        RECT 514.930 1960.290 516.110 1961.470 ;
        RECT 516.530 1960.290 517.710 1961.470 ;
        RECT 514.930 1781.890 516.110 1783.070 ;
        RECT 516.530 1781.890 517.710 1783.070 ;
        RECT 514.930 1780.290 516.110 1781.470 ;
        RECT 516.530 1780.290 517.710 1781.470 ;
        RECT 514.930 1601.890 516.110 1603.070 ;
        RECT 516.530 1601.890 517.710 1603.070 ;
        RECT 514.930 1600.290 516.110 1601.470 ;
        RECT 516.530 1600.290 517.710 1601.470 ;
        RECT 514.930 1421.890 516.110 1423.070 ;
        RECT 516.530 1421.890 517.710 1423.070 ;
        RECT 514.930 1420.290 516.110 1421.470 ;
        RECT 516.530 1420.290 517.710 1421.470 ;
        RECT 514.930 1241.890 516.110 1243.070 ;
        RECT 516.530 1241.890 517.710 1243.070 ;
        RECT 514.930 1240.290 516.110 1241.470 ;
        RECT 516.530 1240.290 517.710 1241.470 ;
        RECT 514.930 1061.890 516.110 1063.070 ;
        RECT 516.530 1061.890 517.710 1063.070 ;
        RECT 514.930 1060.290 516.110 1061.470 ;
        RECT 516.530 1060.290 517.710 1061.470 ;
        RECT 694.930 3556.610 696.110 3557.790 ;
        RECT 696.530 3556.610 697.710 3557.790 ;
        RECT 694.930 3555.010 696.110 3556.190 ;
        RECT 696.530 3555.010 697.710 3556.190 ;
        RECT 694.930 3401.890 696.110 3403.070 ;
        RECT 696.530 3401.890 697.710 3403.070 ;
        RECT 694.930 3400.290 696.110 3401.470 ;
        RECT 696.530 3400.290 697.710 3401.470 ;
        RECT 694.930 3221.890 696.110 3223.070 ;
        RECT 696.530 3221.890 697.710 3223.070 ;
        RECT 694.930 3220.290 696.110 3221.470 ;
        RECT 696.530 3220.290 697.710 3221.470 ;
        RECT 694.930 3041.890 696.110 3043.070 ;
        RECT 696.530 3041.890 697.710 3043.070 ;
        RECT 694.930 3040.290 696.110 3041.470 ;
        RECT 696.530 3040.290 697.710 3041.470 ;
        RECT 694.930 2861.890 696.110 2863.070 ;
        RECT 696.530 2861.890 697.710 2863.070 ;
        RECT 694.930 2860.290 696.110 2861.470 ;
        RECT 696.530 2860.290 697.710 2861.470 ;
        RECT 694.930 2681.890 696.110 2683.070 ;
        RECT 696.530 2681.890 697.710 2683.070 ;
        RECT 694.930 2680.290 696.110 2681.470 ;
        RECT 696.530 2680.290 697.710 2681.470 ;
        RECT 694.930 2501.890 696.110 2503.070 ;
        RECT 696.530 2501.890 697.710 2503.070 ;
        RECT 694.930 2500.290 696.110 2501.470 ;
        RECT 696.530 2500.290 697.710 2501.470 ;
        RECT 694.930 2321.890 696.110 2323.070 ;
        RECT 696.530 2321.890 697.710 2323.070 ;
        RECT 694.930 2320.290 696.110 2321.470 ;
        RECT 696.530 2320.290 697.710 2321.470 ;
        RECT 694.930 2141.890 696.110 2143.070 ;
        RECT 696.530 2141.890 697.710 2143.070 ;
        RECT 694.930 2140.290 696.110 2141.470 ;
        RECT 696.530 2140.290 697.710 2141.470 ;
        RECT 694.930 1961.890 696.110 1963.070 ;
        RECT 696.530 1961.890 697.710 1963.070 ;
        RECT 694.930 1960.290 696.110 1961.470 ;
        RECT 696.530 1960.290 697.710 1961.470 ;
        RECT 694.930 1781.890 696.110 1783.070 ;
        RECT 696.530 1781.890 697.710 1783.070 ;
        RECT 694.930 1780.290 696.110 1781.470 ;
        RECT 696.530 1780.290 697.710 1781.470 ;
        RECT 694.930 1601.890 696.110 1603.070 ;
        RECT 696.530 1601.890 697.710 1603.070 ;
        RECT 694.930 1600.290 696.110 1601.470 ;
        RECT 696.530 1600.290 697.710 1601.470 ;
        RECT 694.930 1421.890 696.110 1423.070 ;
        RECT 696.530 1421.890 697.710 1423.070 ;
        RECT 694.930 1420.290 696.110 1421.470 ;
        RECT 696.530 1420.290 697.710 1421.470 ;
        RECT 694.930 1241.890 696.110 1243.070 ;
        RECT 696.530 1241.890 697.710 1243.070 ;
        RECT 694.930 1240.290 696.110 1241.470 ;
        RECT 696.530 1240.290 697.710 1241.470 ;
        RECT 694.930 1061.890 696.110 1063.070 ;
        RECT 696.530 1061.890 697.710 1063.070 ;
        RECT 694.930 1060.290 696.110 1061.470 ;
        RECT 696.530 1060.290 697.710 1061.470 ;
        RECT 874.930 3556.610 876.110 3557.790 ;
        RECT 876.530 3556.610 877.710 3557.790 ;
        RECT 874.930 3555.010 876.110 3556.190 ;
        RECT 876.530 3555.010 877.710 3556.190 ;
        RECT 874.930 3401.890 876.110 3403.070 ;
        RECT 876.530 3401.890 877.710 3403.070 ;
        RECT 874.930 3400.290 876.110 3401.470 ;
        RECT 876.530 3400.290 877.710 3401.470 ;
        RECT 874.930 3221.890 876.110 3223.070 ;
        RECT 876.530 3221.890 877.710 3223.070 ;
        RECT 874.930 3220.290 876.110 3221.470 ;
        RECT 876.530 3220.290 877.710 3221.470 ;
        RECT 874.930 3041.890 876.110 3043.070 ;
        RECT 876.530 3041.890 877.710 3043.070 ;
        RECT 874.930 3040.290 876.110 3041.470 ;
        RECT 876.530 3040.290 877.710 3041.470 ;
        RECT 874.930 2861.890 876.110 2863.070 ;
        RECT 876.530 2861.890 877.710 2863.070 ;
        RECT 874.930 2860.290 876.110 2861.470 ;
        RECT 876.530 2860.290 877.710 2861.470 ;
        RECT 874.930 2681.890 876.110 2683.070 ;
        RECT 876.530 2681.890 877.710 2683.070 ;
        RECT 874.930 2680.290 876.110 2681.470 ;
        RECT 876.530 2680.290 877.710 2681.470 ;
        RECT 874.930 2501.890 876.110 2503.070 ;
        RECT 876.530 2501.890 877.710 2503.070 ;
        RECT 874.930 2500.290 876.110 2501.470 ;
        RECT 876.530 2500.290 877.710 2501.470 ;
        RECT 874.930 2321.890 876.110 2323.070 ;
        RECT 876.530 2321.890 877.710 2323.070 ;
        RECT 874.930 2320.290 876.110 2321.470 ;
        RECT 876.530 2320.290 877.710 2321.470 ;
        RECT 874.930 2141.890 876.110 2143.070 ;
        RECT 876.530 2141.890 877.710 2143.070 ;
        RECT 874.930 2140.290 876.110 2141.470 ;
        RECT 876.530 2140.290 877.710 2141.470 ;
        RECT 874.930 1961.890 876.110 1963.070 ;
        RECT 876.530 1961.890 877.710 1963.070 ;
        RECT 874.930 1960.290 876.110 1961.470 ;
        RECT 876.530 1960.290 877.710 1961.470 ;
        RECT 874.930 1781.890 876.110 1783.070 ;
        RECT 876.530 1781.890 877.710 1783.070 ;
        RECT 874.930 1780.290 876.110 1781.470 ;
        RECT 876.530 1780.290 877.710 1781.470 ;
        RECT 874.930 1601.890 876.110 1603.070 ;
        RECT 876.530 1601.890 877.710 1603.070 ;
        RECT 874.930 1600.290 876.110 1601.470 ;
        RECT 876.530 1600.290 877.710 1601.470 ;
        RECT 874.930 1421.890 876.110 1423.070 ;
        RECT 876.530 1421.890 877.710 1423.070 ;
        RECT 874.930 1420.290 876.110 1421.470 ;
        RECT 876.530 1420.290 877.710 1421.470 ;
        RECT 874.930 1241.890 876.110 1243.070 ;
        RECT 876.530 1241.890 877.710 1243.070 ;
        RECT 874.930 1240.290 876.110 1241.470 ;
        RECT 876.530 1240.290 877.710 1241.470 ;
        RECT 874.930 1061.890 876.110 1063.070 ;
        RECT 876.530 1061.890 877.710 1063.070 ;
        RECT 874.930 1060.290 876.110 1061.470 ;
        RECT 876.530 1060.290 877.710 1061.470 ;
        RECT 1054.930 3556.610 1056.110 3557.790 ;
        RECT 1056.530 3556.610 1057.710 3557.790 ;
        RECT 1054.930 3555.010 1056.110 3556.190 ;
        RECT 1056.530 3555.010 1057.710 3556.190 ;
        RECT 1054.930 3401.890 1056.110 3403.070 ;
        RECT 1056.530 3401.890 1057.710 3403.070 ;
        RECT 1054.930 3400.290 1056.110 3401.470 ;
        RECT 1056.530 3400.290 1057.710 3401.470 ;
        RECT 1054.930 3221.890 1056.110 3223.070 ;
        RECT 1056.530 3221.890 1057.710 3223.070 ;
        RECT 1054.930 3220.290 1056.110 3221.470 ;
        RECT 1056.530 3220.290 1057.710 3221.470 ;
        RECT 1054.930 3041.890 1056.110 3043.070 ;
        RECT 1056.530 3041.890 1057.710 3043.070 ;
        RECT 1054.930 3040.290 1056.110 3041.470 ;
        RECT 1056.530 3040.290 1057.710 3041.470 ;
        RECT 1054.930 2861.890 1056.110 2863.070 ;
        RECT 1056.530 2861.890 1057.710 2863.070 ;
        RECT 1054.930 2860.290 1056.110 2861.470 ;
        RECT 1056.530 2860.290 1057.710 2861.470 ;
        RECT 1054.930 2681.890 1056.110 2683.070 ;
        RECT 1056.530 2681.890 1057.710 2683.070 ;
        RECT 1054.930 2680.290 1056.110 2681.470 ;
        RECT 1056.530 2680.290 1057.710 2681.470 ;
        RECT 1054.930 2501.890 1056.110 2503.070 ;
        RECT 1056.530 2501.890 1057.710 2503.070 ;
        RECT 1054.930 2500.290 1056.110 2501.470 ;
        RECT 1056.530 2500.290 1057.710 2501.470 ;
        RECT 1054.930 2321.890 1056.110 2323.070 ;
        RECT 1056.530 2321.890 1057.710 2323.070 ;
        RECT 1054.930 2320.290 1056.110 2321.470 ;
        RECT 1056.530 2320.290 1057.710 2321.470 ;
        RECT 1054.930 2141.890 1056.110 2143.070 ;
        RECT 1056.530 2141.890 1057.710 2143.070 ;
        RECT 1054.930 2140.290 1056.110 2141.470 ;
        RECT 1056.530 2140.290 1057.710 2141.470 ;
        RECT 1054.930 1961.890 1056.110 1963.070 ;
        RECT 1056.530 1961.890 1057.710 1963.070 ;
        RECT 1054.930 1960.290 1056.110 1961.470 ;
        RECT 1056.530 1960.290 1057.710 1961.470 ;
        RECT 1054.930 1781.890 1056.110 1783.070 ;
        RECT 1056.530 1781.890 1057.710 1783.070 ;
        RECT 1054.930 1780.290 1056.110 1781.470 ;
        RECT 1056.530 1780.290 1057.710 1781.470 ;
        RECT 1054.930 1601.890 1056.110 1603.070 ;
        RECT 1056.530 1601.890 1057.710 1603.070 ;
        RECT 1054.930 1600.290 1056.110 1601.470 ;
        RECT 1056.530 1600.290 1057.710 1601.470 ;
        RECT 1054.930 1421.890 1056.110 1423.070 ;
        RECT 1056.530 1421.890 1057.710 1423.070 ;
        RECT 1054.930 1420.290 1056.110 1421.470 ;
        RECT 1056.530 1420.290 1057.710 1421.470 ;
        RECT 1054.930 1241.890 1056.110 1243.070 ;
        RECT 1056.530 1241.890 1057.710 1243.070 ;
        RECT 1054.930 1240.290 1056.110 1241.470 ;
        RECT 1056.530 1240.290 1057.710 1241.470 ;
        RECT 1054.930 1061.890 1056.110 1063.070 ;
        RECT 1056.530 1061.890 1057.710 1063.070 ;
        RECT 1054.930 1060.290 1056.110 1061.470 ;
        RECT 1056.530 1060.290 1057.710 1061.470 ;
        RECT 1234.930 3556.610 1236.110 3557.790 ;
        RECT 1236.530 3556.610 1237.710 3557.790 ;
        RECT 1234.930 3555.010 1236.110 3556.190 ;
        RECT 1236.530 3555.010 1237.710 3556.190 ;
        RECT 1234.930 3401.890 1236.110 3403.070 ;
        RECT 1236.530 3401.890 1237.710 3403.070 ;
        RECT 1234.930 3400.290 1236.110 3401.470 ;
        RECT 1236.530 3400.290 1237.710 3401.470 ;
        RECT 1234.930 3221.890 1236.110 3223.070 ;
        RECT 1236.530 3221.890 1237.710 3223.070 ;
        RECT 1234.930 3220.290 1236.110 3221.470 ;
        RECT 1236.530 3220.290 1237.710 3221.470 ;
        RECT 1234.930 3041.890 1236.110 3043.070 ;
        RECT 1236.530 3041.890 1237.710 3043.070 ;
        RECT 1234.930 3040.290 1236.110 3041.470 ;
        RECT 1236.530 3040.290 1237.710 3041.470 ;
        RECT 1234.930 2861.890 1236.110 2863.070 ;
        RECT 1236.530 2861.890 1237.710 2863.070 ;
        RECT 1234.930 2860.290 1236.110 2861.470 ;
        RECT 1236.530 2860.290 1237.710 2861.470 ;
        RECT 1234.930 2681.890 1236.110 2683.070 ;
        RECT 1236.530 2681.890 1237.710 2683.070 ;
        RECT 1234.930 2680.290 1236.110 2681.470 ;
        RECT 1236.530 2680.290 1237.710 2681.470 ;
        RECT 1234.930 2501.890 1236.110 2503.070 ;
        RECT 1236.530 2501.890 1237.710 2503.070 ;
        RECT 1234.930 2500.290 1236.110 2501.470 ;
        RECT 1236.530 2500.290 1237.710 2501.470 ;
        RECT 1234.930 2321.890 1236.110 2323.070 ;
        RECT 1236.530 2321.890 1237.710 2323.070 ;
        RECT 1234.930 2320.290 1236.110 2321.470 ;
        RECT 1236.530 2320.290 1237.710 2321.470 ;
        RECT 1234.930 2141.890 1236.110 2143.070 ;
        RECT 1236.530 2141.890 1237.710 2143.070 ;
        RECT 1234.930 2140.290 1236.110 2141.470 ;
        RECT 1236.530 2140.290 1237.710 2141.470 ;
        RECT 1234.930 1961.890 1236.110 1963.070 ;
        RECT 1236.530 1961.890 1237.710 1963.070 ;
        RECT 1234.930 1960.290 1236.110 1961.470 ;
        RECT 1236.530 1960.290 1237.710 1961.470 ;
        RECT 1234.930 1781.890 1236.110 1783.070 ;
        RECT 1236.530 1781.890 1237.710 1783.070 ;
        RECT 1234.930 1780.290 1236.110 1781.470 ;
        RECT 1236.530 1780.290 1237.710 1781.470 ;
        RECT 1234.930 1601.890 1236.110 1603.070 ;
        RECT 1236.530 1601.890 1237.710 1603.070 ;
        RECT 1234.930 1600.290 1236.110 1601.470 ;
        RECT 1236.530 1600.290 1237.710 1601.470 ;
        RECT 1234.930 1421.890 1236.110 1423.070 ;
        RECT 1236.530 1421.890 1237.710 1423.070 ;
        RECT 1234.930 1420.290 1236.110 1421.470 ;
        RECT 1236.530 1420.290 1237.710 1421.470 ;
        RECT 1234.930 1241.890 1236.110 1243.070 ;
        RECT 1236.530 1241.890 1237.710 1243.070 ;
        RECT 1234.930 1240.290 1236.110 1241.470 ;
        RECT 1236.530 1240.290 1237.710 1241.470 ;
        RECT 1234.930 1061.890 1236.110 1063.070 ;
        RECT 1236.530 1061.890 1237.710 1063.070 ;
        RECT 1234.930 1060.290 1236.110 1061.470 ;
        RECT 1236.530 1060.290 1237.710 1061.470 ;
        RECT 154.930 881.890 156.110 883.070 ;
        RECT 156.530 881.890 157.710 883.070 ;
        RECT 154.930 880.290 156.110 881.470 ;
        RECT 156.530 880.290 157.710 881.470 ;
        RECT 154.930 701.890 156.110 703.070 ;
        RECT 156.530 701.890 157.710 703.070 ;
        RECT 154.930 700.290 156.110 701.470 ;
        RECT 156.530 700.290 157.710 701.470 ;
        RECT 154.930 521.890 156.110 523.070 ;
        RECT 156.530 521.890 157.710 523.070 ;
        RECT 154.930 520.290 156.110 521.470 ;
        RECT 156.530 520.290 157.710 521.470 ;
        RECT 1234.930 881.890 1236.110 883.070 ;
        RECT 1236.530 881.890 1237.710 883.070 ;
        RECT 1234.930 880.290 1236.110 881.470 ;
        RECT 1236.530 880.290 1237.710 881.470 ;
        RECT 1234.930 701.890 1236.110 703.070 ;
        RECT 1236.530 701.890 1237.710 703.070 ;
        RECT 1234.930 700.290 1236.110 701.470 ;
        RECT 1236.530 700.290 1237.710 701.470 ;
        RECT 1234.930 521.890 1236.110 523.070 ;
        RECT 1236.530 521.890 1237.710 523.070 ;
        RECT 1234.930 520.290 1236.110 521.470 ;
        RECT 1236.530 520.290 1237.710 521.470 ;
        RECT 154.930 341.890 156.110 343.070 ;
        RECT 156.530 341.890 157.710 343.070 ;
        RECT 154.930 340.290 156.110 341.470 ;
        RECT 156.530 340.290 157.710 341.470 ;
        RECT 154.930 161.890 156.110 163.070 ;
        RECT 156.530 161.890 157.710 163.070 ;
        RECT 154.930 160.290 156.110 161.470 ;
        RECT 156.530 160.290 157.710 161.470 ;
        RECT 154.930 -36.510 156.110 -35.330 ;
        RECT 156.530 -36.510 157.710 -35.330 ;
        RECT 154.930 -38.110 156.110 -36.930 ;
        RECT 156.530 -38.110 157.710 -36.930 ;
        RECT 334.930 341.890 336.110 343.070 ;
        RECT 336.530 341.890 337.710 343.070 ;
        RECT 334.930 340.290 336.110 341.470 ;
        RECT 336.530 340.290 337.710 341.470 ;
        RECT 334.930 161.890 336.110 163.070 ;
        RECT 336.530 161.890 337.710 163.070 ;
        RECT 334.930 160.290 336.110 161.470 ;
        RECT 336.530 160.290 337.710 161.470 ;
        RECT 334.930 -36.510 336.110 -35.330 ;
        RECT 336.530 -36.510 337.710 -35.330 ;
        RECT 334.930 -38.110 336.110 -36.930 ;
        RECT 336.530 -38.110 337.710 -36.930 ;
        RECT 514.930 341.890 516.110 343.070 ;
        RECT 516.530 341.890 517.710 343.070 ;
        RECT 514.930 340.290 516.110 341.470 ;
        RECT 516.530 340.290 517.710 341.470 ;
        RECT 514.930 161.890 516.110 163.070 ;
        RECT 516.530 161.890 517.710 163.070 ;
        RECT 514.930 160.290 516.110 161.470 ;
        RECT 516.530 160.290 517.710 161.470 ;
        RECT 514.930 -36.510 516.110 -35.330 ;
        RECT 516.530 -36.510 517.710 -35.330 ;
        RECT 514.930 -38.110 516.110 -36.930 ;
        RECT 516.530 -38.110 517.710 -36.930 ;
        RECT 694.930 341.890 696.110 343.070 ;
        RECT 696.530 341.890 697.710 343.070 ;
        RECT 694.930 340.290 696.110 341.470 ;
        RECT 696.530 340.290 697.710 341.470 ;
        RECT 694.930 161.890 696.110 163.070 ;
        RECT 696.530 161.890 697.710 163.070 ;
        RECT 694.930 160.290 696.110 161.470 ;
        RECT 696.530 160.290 697.710 161.470 ;
        RECT 694.930 -36.510 696.110 -35.330 ;
        RECT 696.530 -36.510 697.710 -35.330 ;
        RECT 694.930 -38.110 696.110 -36.930 ;
        RECT 696.530 -38.110 697.710 -36.930 ;
        RECT 874.930 341.890 876.110 343.070 ;
        RECT 876.530 341.890 877.710 343.070 ;
        RECT 874.930 340.290 876.110 341.470 ;
        RECT 876.530 340.290 877.710 341.470 ;
        RECT 874.930 161.890 876.110 163.070 ;
        RECT 876.530 161.890 877.710 163.070 ;
        RECT 874.930 160.290 876.110 161.470 ;
        RECT 876.530 160.290 877.710 161.470 ;
        RECT 874.930 -36.510 876.110 -35.330 ;
        RECT 876.530 -36.510 877.710 -35.330 ;
        RECT 874.930 -38.110 876.110 -36.930 ;
        RECT 876.530 -38.110 877.710 -36.930 ;
        RECT 1054.930 341.890 1056.110 343.070 ;
        RECT 1056.530 341.890 1057.710 343.070 ;
        RECT 1054.930 340.290 1056.110 341.470 ;
        RECT 1056.530 340.290 1057.710 341.470 ;
        RECT 1054.930 161.890 1056.110 163.070 ;
        RECT 1056.530 161.890 1057.710 163.070 ;
        RECT 1054.930 160.290 1056.110 161.470 ;
        RECT 1056.530 160.290 1057.710 161.470 ;
        RECT 1054.930 -36.510 1056.110 -35.330 ;
        RECT 1056.530 -36.510 1057.710 -35.330 ;
        RECT 1054.930 -38.110 1056.110 -36.930 ;
        RECT 1056.530 -38.110 1057.710 -36.930 ;
        RECT 1234.930 341.890 1236.110 343.070 ;
        RECT 1236.530 341.890 1237.710 343.070 ;
        RECT 1234.930 340.290 1236.110 341.470 ;
        RECT 1236.530 340.290 1237.710 341.470 ;
        RECT 1234.930 161.890 1236.110 163.070 ;
        RECT 1236.530 161.890 1237.710 163.070 ;
        RECT 1234.930 160.290 1236.110 161.470 ;
        RECT 1236.530 160.290 1237.710 161.470 ;
        RECT 1234.930 -36.510 1236.110 -35.330 ;
        RECT 1236.530 -36.510 1237.710 -35.330 ;
        RECT 1234.930 -38.110 1236.110 -36.930 ;
        RECT 1236.530 -38.110 1237.710 -36.930 ;
        RECT 1414.930 3556.610 1416.110 3557.790 ;
        RECT 1416.530 3556.610 1417.710 3557.790 ;
        RECT 1414.930 3555.010 1416.110 3556.190 ;
        RECT 1416.530 3555.010 1417.710 3556.190 ;
        RECT 1414.930 3401.890 1416.110 3403.070 ;
        RECT 1416.530 3401.890 1417.710 3403.070 ;
        RECT 1414.930 3400.290 1416.110 3401.470 ;
        RECT 1416.530 3400.290 1417.710 3401.470 ;
        RECT 1414.930 3221.890 1416.110 3223.070 ;
        RECT 1416.530 3221.890 1417.710 3223.070 ;
        RECT 1414.930 3220.290 1416.110 3221.470 ;
        RECT 1416.530 3220.290 1417.710 3221.470 ;
        RECT 1414.930 3041.890 1416.110 3043.070 ;
        RECT 1416.530 3041.890 1417.710 3043.070 ;
        RECT 1414.930 3040.290 1416.110 3041.470 ;
        RECT 1416.530 3040.290 1417.710 3041.470 ;
        RECT 1414.930 2861.890 1416.110 2863.070 ;
        RECT 1416.530 2861.890 1417.710 2863.070 ;
        RECT 1414.930 2860.290 1416.110 2861.470 ;
        RECT 1416.530 2860.290 1417.710 2861.470 ;
        RECT 1414.930 2681.890 1416.110 2683.070 ;
        RECT 1416.530 2681.890 1417.710 2683.070 ;
        RECT 1414.930 2680.290 1416.110 2681.470 ;
        RECT 1416.530 2680.290 1417.710 2681.470 ;
        RECT 1414.930 2501.890 1416.110 2503.070 ;
        RECT 1416.530 2501.890 1417.710 2503.070 ;
        RECT 1414.930 2500.290 1416.110 2501.470 ;
        RECT 1416.530 2500.290 1417.710 2501.470 ;
        RECT 1414.930 2321.890 1416.110 2323.070 ;
        RECT 1416.530 2321.890 1417.710 2323.070 ;
        RECT 1414.930 2320.290 1416.110 2321.470 ;
        RECT 1416.530 2320.290 1417.710 2321.470 ;
        RECT 1414.930 2141.890 1416.110 2143.070 ;
        RECT 1416.530 2141.890 1417.710 2143.070 ;
        RECT 1414.930 2140.290 1416.110 2141.470 ;
        RECT 1416.530 2140.290 1417.710 2141.470 ;
        RECT 1414.930 1961.890 1416.110 1963.070 ;
        RECT 1416.530 1961.890 1417.710 1963.070 ;
        RECT 1414.930 1960.290 1416.110 1961.470 ;
        RECT 1416.530 1960.290 1417.710 1961.470 ;
        RECT 1414.930 1781.890 1416.110 1783.070 ;
        RECT 1416.530 1781.890 1417.710 1783.070 ;
        RECT 1414.930 1780.290 1416.110 1781.470 ;
        RECT 1416.530 1780.290 1417.710 1781.470 ;
        RECT 1414.930 1601.890 1416.110 1603.070 ;
        RECT 1416.530 1601.890 1417.710 1603.070 ;
        RECT 1414.930 1600.290 1416.110 1601.470 ;
        RECT 1416.530 1600.290 1417.710 1601.470 ;
        RECT 1414.930 1421.890 1416.110 1423.070 ;
        RECT 1416.530 1421.890 1417.710 1423.070 ;
        RECT 1414.930 1420.290 1416.110 1421.470 ;
        RECT 1416.530 1420.290 1417.710 1421.470 ;
        RECT 1414.930 1241.890 1416.110 1243.070 ;
        RECT 1416.530 1241.890 1417.710 1243.070 ;
        RECT 1414.930 1240.290 1416.110 1241.470 ;
        RECT 1416.530 1240.290 1417.710 1241.470 ;
        RECT 1414.930 1061.890 1416.110 1063.070 ;
        RECT 1416.530 1061.890 1417.710 1063.070 ;
        RECT 1414.930 1060.290 1416.110 1061.470 ;
        RECT 1416.530 1060.290 1417.710 1061.470 ;
        RECT 1414.930 881.890 1416.110 883.070 ;
        RECT 1416.530 881.890 1417.710 883.070 ;
        RECT 1414.930 880.290 1416.110 881.470 ;
        RECT 1416.530 880.290 1417.710 881.470 ;
        RECT 1414.930 701.890 1416.110 703.070 ;
        RECT 1416.530 701.890 1417.710 703.070 ;
        RECT 1414.930 700.290 1416.110 701.470 ;
        RECT 1416.530 700.290 1417.710 701.470 ;
        RECT 1414.930 521.890 1416.110 523.070 ;
        RECT 1416.530 521.890 1417.710 523.070 ;
        RECT 1414.930 520.290 1416.110 521.470 ;
        RECT 1416.530 520.290 1417.710 521.470 ;
        RECT 1414.930 341.890 1416.110 343.070 ;
        RECT 1416.530 341.890 1417.710 343.070 ;
        RECT 1414.930 340.290 1416.110 341.470 ;
        RECT 1416.530 340.290 1417.710 341.470 ;
        RECT 1414.930 161.890 1416.110 163.070 ;
        RECT 1416.530 161.890 1417.710 163.070 ;
        RECT 1414.930 160.290 1416.110 161.470 ;
        RECT 1416.530 160.290 1417.710 161.470 ;
        RECT 1414.930 -36.510 1416.110 -35.330 ;
        RECT 1416.530 -36.510 1417.710 -35.330 ;
        RECT 1414.930 -38.110 1416.110 -36.930 ;
        RECT 1416.530 -38.110 1417.710 -36.930 ;
        RECT 1594.930 3556.610 1596.110 3557.790 ;
        RECT 1596.530 3556.610 1597.710 3557.790 ;
        RECT 1594.930 3555.010 1596.110 3556.190 ;
        RECT 1596.530 3555.010 1597.710 3556.190 ;
        RECT 1594.930 3401.890 1596.110 3403.070 ;
        RECT 1596.530 3401.890 1597.710 3403.070 ;
        RECT 1594.930 3400.290 1596.110 3401.470 ;
        RECT 1596.530 3400.290 1597.710 3401.470 ;
        RECT 1594.930 3221.890 1596.110 3223.070 ;
        RECT 1596.530 3221.890 1597.710 3223.070 ;
        RECT 1594.930 3220.290 1596.110 3221.470 ;
        RECT 1596.530 3220.290 1597.710 3221.470 ;
        RECT 1594.930 3041.890 1596.110 3043.070 ;
        RECT 1596.530 3041.890 1597.710 3043.070 ;
        RECT 1594.930 3040.290 1596.110 3041.470 ;
        RECT 1596.530 3040.290 1597.710 3041.470 ;
        RECT 1594.930 2861.890 1596.110 2863.070 ;
        RECT 1596.530 2861.890 1597.710 2863.070 ;
        RECT 1594.930 2860.290 1596.110 2861.470 ;
        RECT 1596.530 2860.290 1597.710 2861.470 ;
        RECT 1594.930 2681.890 1596.110 2683.070 ;
        RECT 1596.530 2681.890 1597.710 2683.070 ;
        RECT 1594.930 2680.290 1596.110 2681.470 ;
        RECT 1596.530 2680.290 1597.710 2681.470 ;
        RECT 1594.930 2501.890 1596.110 2503.070 ;
        RECT 1596.530 2501.890 1597.710 2503.070 ;
        RECT 1594.930 2500.290 1596.110 2501.470 ;
        RECT 1596.530 2500.290 1597.710 2501.470 ;
        RECT 1594.930 2321.890 1596.110 2323.070 ;
        RECT 1596.530 2321.890 1597.710 2323.070 ;
        RECT 1594.930 2320.290 1596.110 2321.470 ;
        RECT 1596.530 2320.290 1597.710 2321.470 ;
        RECT 1594.930 2141.890 1596.110 2143.070 ;
        RECT 1596.530 2141.890 1597.710 2143.070 ;
        RECT 1594.930 2140.290 1596.110 2141.470 ;
        RECT 1596.530 2140.290 1597.710 2141.470 ;
        RECT 1594.930 1961.890 1596.110 1963.070 ;
        RECT 1596.530 1961.890 1597.710 1963.070 ;
        RECT 1594.930 1960.290 1596.110 1961.470 ;
        RECT 1596.530 1960.290 1597.710 1961.470 ;
        RECT 1594.930 1781.890 1596.110 1783.070 ;
        RECT 1596.530 1781.890 1597.710 1783.070 ;
        RECT 1594.930 1780.290 1596.110 1781.470 ;
        RECT 1596.530 1780.290 1597.710 1781.470 ;
        RECT 1594.930 1601.890 1596.110 1603.070 ;
        RECT 1596.530 1601.890 1597.710 1603.070 ;
        RECT 1594.930 1600.290 1596.110 1601.470 ;
        RECT 1596.530 1600.290 1597.710 1601.470 ;
        RECT 1594.930 1421.890 1596.110 1423.070 ;
        RECT 1596.530 1421.890 1597.710 1423.070 ;
        RECT 1594.930 1420.290 1596.110 1421.470 ;
        RECT 1596.530 1420.290 1597.710 1421.470 ;
        RECT 1594.930 1241.890 1596.110 1243.070 ;
        RECT 1596.530 1241.890 1597.710 1243.070 ;
        RECT 1594.930 1240.290 1596.110 1241.470 ;
        RECT 1596.530 1240.290 1597.710 1241.470 ;
        RECT 1594.930 1061.890 1596.110 1063.070 ;
        RECT 1596.530 1061.890 1597.710 1063.070 ;
        RECT 1594.930 1060.290 1596.110 1061.470 ;
        RECT 1596.530 1060.290 1597.710 1061.470 ;
        RECT 1594.930 881.890 1596.110 883.070 ;
        RECT 1596.530 881.890 1597.710 883.070 ;
        RECT 1594.930 880.290 1596.110 881.470 ;
        RECT 1596.530 880.290 1597.710 881.470 ;
        RECT 1594.930 701.890 1596.110 703.070 ;
        RECT 1596.530 701.890 1597.710 703.070 ;
        RECT 1594.930 700.290 1596.110 701.470 ;
        RECT 1596.530 700.290 1597.710 701.470 ;
        RECT 1594.930 521.890 1596.110 523.070 ;
        RECT 1596.530 521.890 1597.710 523.070 ;
        RECT 1594.930 520.290 1596.110 521.470 ;
        RECT 1596.530 520.290 1597.710 521.470 ;
        RECT 1594.930 341.890 1596.110 343.070 ;
        RECT 1596.530 341.890 1597.710 343.070 ;
        RECT 1594.930 340.290 1596.110 341.470 ;
        RECT 1596.530 340.290 1597.710 341.470 ;
        RECT 1594.930 161.890 1596.110 163.070 ;
        RECT 1596.530 161.890 1597.710 163.070 ;
        RECT 1594.930 160.290 1596.110 161.470 ;
        RECT 1596.530 160.290 1597.710 161.470 ;
        RECT 1594.930 -36.510 1596.110 -35.330 ;
        RECT 1596.530 -36.510 1597.710 -35.330 ;
        RECT 1594.930 -38.110 1596.110 -36.930 ;
        RECT 1596.530 -38.110 1597.710 -36.930 ;
        RECT 1774.930 3556.610 1776.110 3557.790 ;
        RECT 1776.530 3556.610 1777.710 3557.790 ;
        RECT 1774.930 3555.010 1776.110 3556.190 ;
        RECT 1776.530 3555.010 1777.710 3556.190 ;
        RECT 1774.930 3401.890 1776.110 3403.070 ;
        RECT 1776.530 3401.890 1777.710 3403.070 ;
        RECT 1774.930 3400.290 1776.110 3401.470 ;
        RECT 1776.530 3400.290 1777.710 3401.470 ;
        RECT 1774.930 3221.890 1776.110 3223.070 ;
        RECT 1776.530 3221.890 1777.710 3223.070 ;
        RECT 1774.930 3220.290 1776.110 3221.470 ;
        RECT 1776.530 3220.290 1777.710 3221.470 ;
        RECT 1774.930 3041.890 1776.110 3043.070 ;
        RECT 1776.530 3041.890 1777.710 3043.070 ;
        RECT 1774.930 3040.290 1776.110 3041.470 ;
        RECT 1776.530 3040.290 1777.710 3041.470 ;
        RECT 1774.930 2861.890 1776.110 2863.070 ;
        RECT 1776.530 2861.890 1777.710 2863.070 ;
        RECT 1774.930 2860.290 1776.110 2861.470 ;
        RECT 1776.530 2860.290 1777.710 2861.470 ;
        RECT 1774.930 2681.890 1776.110 2683.070 ;
        RECT 1776.530 2681.890 1777.710 2683.070 ;
        RECT 1774.930 2680.290 1776.110 2681.470 ;
        RECT 1776.530 2680.290 1777.710 2681.470 ;
        RECT 1774.930 2501.890 1776.110 2503.070 ;
        RECT 1776.530 2501.890 1777.710 2503.070 ;
        RECT 1774.930 2500.290 1776.110 2501.470 ;
        RECT 1776.530 2500.290 1777.710 2501.470 ;
        RECT 1774.930 2321.890 1776.110 2323.070 ;
        RECT 1776.530 2321.890 1777.710 2323.070 ;
        RECT 1774.930 2320.290 1776.110 2321.470 ;
        RECT 1776.530 2320.290 1777.710 2321.470 ;
        RECT 1774.930 2141.890 1776.110 2143.070 ;
        RECT 1776.530 2141.890 1777.710 2143.070 ;
        RECT 1774.930 2140.290 1776.110 2141.470 ;
        RECT 1776.530 2140.290 1777.710 2141.470 ;
        RECT 1774.930 1961.890 1776.110 1963.070 ;
        RECT 1776.530 1961.890 1777.710 1963.070 ;
        RECT 1774.930 1960.290 1776.110 1961.470 ;
        RECT 1776.530 1960.290 1777.710 1961.470 ;
        RECT 1774.930 1781.890 1776.110 1783.070 ;
        RECT 1776.530 1781.890 1777.710 1783.070 ;
        RECT 1774.930 1780.290 1776.110 1781.470 ;
        RECT 1776.530 1780.290 1777.710 1781.470 ;
        RECT 1774.930 1601.890 1776.110 1603.070 ;
        RECT 1776.530 1601.890 1777.710 1603.070 ;
        RECT 1774.930 1600.290 1776.110 1601.470 ;
        RECT 1776.530 1600.290 1777.710 1601.470 ;
        RECT 1774.930 1421.890 1776.110 1423.070 ;
        RECT 1776.530 1421.890 1777.710 1423.070 ;
        RECT 1774.930 1420.290 1776.110 1421.470 ;
        RECT 1776.530 1420.290 1777.710 1421.470 ;
        RECT 1774.930 1241.890 1776.110 1243.070 ;
        RECT 1776.530 1241.890 1777.710 1243.070 ;
        RECT 1774.930 1240.290 1776.110 1241.470 ;
        RECT 1776.530 1240.290 1777.710 1241.470 ;
        RECT 1774.930 1061.890 1776.110 1063.070 ;
        RECT 1776.530 1061.890 1777.710 1063.070 ;
        RECT 1774.930 1060.290 1776.110 1061.470 ;
        RECT 1776.530 1060.290 1777.710 1061.470 ;
        RECT 1774.930 881.890 1776.110 883.070 ;
        RECT 1776.530 881.890 1777.710 883.070 ;
        RECT 1774.930 880.290 1776.110 881.470 ;
        RECT 1776.530 880.290 1777.710 881.470 ;
        RECT 1774.930 701.890 1776.110 703.070 ;
        RECT 1776.530 701.890 1777.710 703.070 ;
        RECT 1774.930 700.290 1776.110 701.470 ;
        RECT 1776.530 700.290 1777.710 701.470 ;
        RECT 1774.930 521.890 1776.110 523.070 ;
        RECT 1776.530 521.890 1777.710 523.070 ;
        RECT 1774.930 520.290 1776.110 521.470 ;
        RECT 1776.530 520.290 1777.710 521.470 ;
        RECT 1774.930 341.890 1776.110 343.070 ;
        RECT 1776.530 341.890 1777.710 343.070 ;
        RECT 1774.930 340.290 1776.110 341.470 ;
        RECT 1776.530 340.290 1777.710 341.470 ;
        RECT 1774.930 161.890 1776.110 163.070 ;
        RECT 1776.530 161.890 1777.710 163.070 ;
        RECT 1774.930 160.290 1776.110 161.470 ;
        RECT 1776.530 160.290 1777.710 161.470 ;
        RECT 1774.930 -36.510 1776.110 -35.330 ;
        RECT 1776.530 -36.510 1777.710 -35.330 ;
        RECT 1774.930 -38.110 1776.110 -36.930 ;
        RECT 1776.530 -38.110 1777.710 -36.930 ;
        RECT 1954.930 3556.610 1956.110 3557.790 ;
        RECT 1956.530 3556.610 1957.710 3557.790 ;
        RECT 1954.930 3555.010 1956.110 3556.190 ;
        RECT 1956.530 3555.010 1957.710 3556.190 ;
        RECT 1954.930 3401.890 1956.110 3403.070 ;
        RECT 1956.530 3401.890 1957.710 3403.070 ;
        RECT 1954.930 3400.290 1956.110 3401.470 ;
        RECT 1956.530 3400.290 1957.710 3401.470 ;
        RECT 1954.930 3221.890 1956.110 3223.070 ;
        RECT 1956.530 3221.890 1957.710 3223.070 ;
        RECT 1954.930 3220.290 1956.110 3221.470 ;
        RECT 1956.530 3220.290 1957.710 3221.470 ;
        RECT 1954.930 3041.890 1956.110 3043.070 ;
        RECT 1956.530 3041.890 1957.710 3043.070 ;
        RECT 1954.930 3040.290 1956.110 3041.470 ;
        RECT 1956.530 3040.290 1957.710 3041.470 ;
        RECT 1954.930 2861.890 1956.110 2863.070 ;
        RECT 1956.530 2861.890 1957.710 2863.070 ;
        RECT 1954.930 2860.290 1956.110 2861.470 ;
        RECT 1956.530 2860.290 1957.710 2861.470 ;
        RECT 1954.930 2681.890 1956.110 2683.070 ;
        RECT 1956.530 2681.890 1957.710 2683.070 ;
        RECT 1954.930 2680.290 1956.110 2681.470 ;
        RECT 1956.530 2680.290 1957.710 2681.470 ;
        RECT 1954.930 2501.890 1956.110 2503.070 ;
        RECT 1956.530 2501.890 1957.710 2503.070 ;
        RECT 1954.930 2500.290 1956.110 2501.470 ;
        RECT 1956.530 2500.290 1957.710 2501.470 ;
        RECT 1954.930 2321.890 1956.110 2323.070 ;
        RECT 1956.530 2321.890 1957.710 2323.070 ;
        RECT 1954.930 2320.290 1956.110 2321.470 ;
        RECT 1956.530 2320.290 1957.710 2321.470 ;
        RECT 1954.930 2141.890 1956.110 2143.070 ;
        RECT 1956.530 2141.890 1957.710 2143.070 ;
        RECT 1954.930 2140.290 1956.110 2141.470 ;
        RECT 1956.530 2140.290 1957.710 2141.470 ;
        RECT 1954.930 1961.890 1956.110 1963.070 ;
        RECT 1956.530 1961.890 1957.710 1963.070 ;
        RECT 1954.930 1960.290 1956.110 1961.470 ;
        RECT 1956.530 1960.290 1957.710 1961.470 ;
        RECT 1954.930 1781.890 1956.110 1783.070 ;
        RECT 1956.530 1781.890 1957.710 1783.070 ;
        RECT 1954.930 1780.290 1956.110 1781.470 ;
        RECT 1956.530 1780.290 1957.710 1781.470 ;
        RECT 1954.930 1601.890 1956.110 1603.070 ;
        RECT 1956.530 1601.890 1957.710 1603.070 ;
        RECT 1954.930 1600.290 1956.110 1601.470 ;
        RECT 1956.530 1600.290 1957.710 1601.470 ;
        RECT 1954.930 1421.890 1956.110 1423.070 ;
        RECT 1956.530 1421.890 1957.710 1423.070 ;
        RECT 1954.930 1420.290 1956.110 1421.470 ;
        RECT 1956.530 1420.290 1957.710 1421.470 ;
        RECT 1954.930 1241.890 1956.110 1243.070 ;
        RECT 1956.530 1241.890 1957.710 1243.070 ;
        RECT 1954.930 1240.290 1956.110 1241.470 ;
        RECT 1956.530 1240.290 1957.710 1241.470 ;
        RECT 1954.930 1061.890 1956.110 1063.070 ;
        RECT 1956.530 1061.890 1957.710 1063.070 ;
        RECT 1954.930 1060.290 1956.110 1061.470 ;
        RECT 1956.530 1060.290 1957.710 1061.470 ;
        RECT 1954.930 881.890 1956.110 883.070 ;
        RECT 1956.530 881.890 1957.710 883.070 ;
        RECT 1954.930 880.290 1956.110 881.470 ;
        RECT 1956.530 880.290 1957.710 881.470 ;
        RECT 1954.930 701.890 1956.110 703.070 ;
        RECT 1956.530 701.890 1957.710 703.070 ;
        RECT 1954.930 700.290 1956.110 701.470 ;
        RECT 1956.530 700.290 1957.710 701.470 ;
        RECT 1954.930 521.890 1956.110 523.070 ;
        RECT 1956.530 521.890 1957.710 523.070 ;
        RECT 1954.930 520.290 1956.110 521.470 ;
        RECT 1956.530 520.290 1957.710 521.470 ;
        RECT 1954.930 341.890 1956.110 343.070 ;
        RECT 1956.530 341.890 1957.710 343.070 ;
        RECT 1954.930 340.290 1956.110 341.470 ;
        RECT 1956.530 340.290 1957.710 341.470 ;
        RECT 1954.930 161.890 1956.110 163.070 ;
        RECT 1956.530 161.890 1957.710 163.070 ;
        RECT 1954.930 160.290 1956.110 161.470 ;
        RECT 1956.530 160.290 1957.710 161.470 ;
        RECT 1954.930 -36.510 1956.110 -35.330 ;
        RECT 1956.530 -36.510 1957.710 -35.330 ;
        RECT 1954.930 -38.110 1956.110 -36.930 ;
        RECT 1956.530 -38.110 1957.710 -36.930 ;
        RECT 2134.930 3556.610 2136.110 3557.790 ;
        RECT 2136.530 3556.610 2137.710 3557.790 ;
        RECT 2134.930 3555.010 2136.110 3556.190 ;
        RECT 2136.530 3555.010 2137.710 3556.190 ;
        RECT 2134.930 3401.890 2136.110 3403.070 ;
        RECT 2136.530 3401.890 2137.710 3403.070 ;
        RECT 2134.930 3400.290 2136.110 3401.470 ;
        RECT 2136.530 3400.290 2137.710 3401.470 ;
        RECT 2134.930 3221.890 2136.110 3223.070 ;
        RECT 2136.530 3221.890 2137.710 3223.070 ;
        RECT 2134.930 3220.290 2136.110 3221.470 ;
        RECT 2136.530 3220.290 2137.710 3221.470 ;
        RECT 2134.930 3041.890 2136.110 3043.070 ;
        RECT 2136.530 3041.890 2137.710 3043.070 ;
        RECT 2134.930 3040.290 2136.110 3041.470 ;
        RECT 2136.530 3040.290 2137.710 3041.470 ;
        RECT 2134.930 2861.890 2136.110 2863.070 ;
        RECT 2136.530 2861.890 2137.710 2863.070 ;
        RECT 2134.930 2860.290 2136.110 2861.470 ;
        RECT 2136.530 2860.290 2137.710 2861.470 ;
        RECT 2134.930 2681.890 2136.110 2683.070 ;
        RECT 2136.530 2681.890 2137.710 2683.070 ;
        RECT 2134.930 2680.290 2136.110 2681.470 ;
        RECT 2136.530 2680.290 2137.710 2681.470 ;
        RECT 2134.930 2501.890 2136.110 2503.070 ;
        RECT 2136.530 2501.890 2137.710 2503.070 ;
        RECT 2134.930 2500.290 2136.110 2501.470 ;
        RECT 2136.530 2500.290 2137.710 2501.470 ;
        RECT 2134.930 2321.890 2136.110 2323.070 ;
        RECT 2136.530 2321.890 2137.710 2323.070 ;
        RECT 2134.930 2320.290 2136.110 2321.470 ;
        RECT 2136.530 2320.290 2137.710 2321.470 ;
        RECT 2134.930 2141.890 2136.110 2143.070 ;
        RECT 2136.530 2141.890 2137.710 2143.070 ;
        RECT 2134.930 2140.290 2136.110 2141.470 ;
        RECT 2136.530 2140.290 2137.710 2141.470 ;
        RECT 2134.930 1961.890 2136.110 1963.070 ;
        RECT 2136.530 1961.890 2137.710 1963.070 ;
        RECT 2134.930 1960.290 2136.110 1961.470 ;
        RECT 2136.530 1960.290 2137.710 1961.470 ;
        RECT 2134.930 1781.890 2136.110 1783.070 ;
        RECT 2136.530 1781.890 2137.710 1783.070 ;
        RECT 2134.930 1780.290 2136.110 1781.470 ;
        RECT 2136.530 1780.290 2137.710 1781.470 ;
        RECT 2134.930 1601.890 2136.110 1603.070 ;
        RECT 2136.530 1601.890 2137.710 1603.070 ;
        RECT 2134.930 1600.290 2136.110 1601.470 ;
        RECT 2136.530 1600.290 2137.710 1601.470 ;
        RECT 2134.930 1421.890 2136.110 1423.070 ;
        RECT 2136.530 1421.890 2137.710 1423.070 ;
        RECT 2134.930 1420.290 2136.110 1421.470 ;
        RECT 2136.530 1420.290 2137.710 1421.470 ;
        RECT 2134.930 1241.890 2136.110 1243.070 ;
        RECT 2136.530 1241.890 2137.710 1243.070 ;
        RECT 2134.930 1240.290 2136.110 1241.470 ;
        RECT 2136.530 1240.290 2137.710 1241.470 ;
        RECT 2134.930 1061.890 2136.110 1063.070 ;
        RECT 2136.530 1061.890 2137.710 1063.070 ;
        RECT 2134.930 1060.290 2136.110 1061.470 ;
        RECT 2136.530 1060.290 2137.710 1061.470 ;
        RECT 2134.930 881.890 2136.110 883.070 ;
        RECT 2136.530 881.890 2137.710 883.070 ;
        RECT 2134.930 880.290 2136.110 881.470 ;
        RECT 2136.530 880.290 2137.710 881.470 ;
        RECT 2134.930 701.890 2136.110 703.070 ;
        RECT 2136.530 701.890 2137.710 703.070 ;
        RECT 2134.930 700.290 2136.110 701.470 ;
        RECT 2136.530 700.290 2137.710 701.470 ;
        RECT 2134.930 521.890 2136.110 523.070 ;
        RECT 2136.530 521.890 2137.710 523.070 ;
        RECT 2134.930 520.290 2136.110 521.470 ;
        RECT 2136.530 520.290 2137.710 521.470 ;
        RECT 2134.930 341.890 2136.110 343.070 ;
        RECT 2136.530 341.890 2137.710 343.070 ;
        RECT 2134.930 340.290 2136.110 341.470 ;
        RECT 2136.530 340.290 2137.710 341.470 ;
        RECT 2134.930 161.890 2136.110 163.070 ;
        RECT 2136.530 161.890 2137.710 163.070 ;
        RECT 2134.930 160.290 2136.110 161.470 ;
        RECT 2136.530 160.290 2137.710 161.470 ;
        RECT 2134.930 -36.510 2136.110 -35.330 ;
        RECT 2136.530 -36.510 2137.710 -35.330 ;
        RECT 2134.930 -38.110 2136.110 -36.930 ;
        RECT 2136.530 -38.110 2137.710 -36.930 ;
        RECT 2314.930 3556.610 2316.110 3557.790 ;
        RECT 2316.530 3556.610 2317.710 3557.790 ;
        RECT 2314.930 3555.010 2316.110 3556.190 ;
        RECT 2316.530 3555.010 2317.710 3556.190 ;
        RECT 2314.930 3401.890 2316.110 3403.070 ;
        RECT 2316.530 3401.890 2317.710 3403.070 ;
        RECT 2314.930 3400.290 2316.110 3401.470 ;
        RECT 2316.530 3400.290 2317.710 3401.470 ;
        RECT 2314.930 3221.890 2316.110 3223.070 ;
        RECT 2316.530 3221.890 2317.710 3223.070 ;
        RECT 2314.930 3220.290 2316.110 3221.470 ;
        RECT 2316.530 3220.290 2317.710 3221.470 ;
        RECT 2314.930 3041.890 2316.110 3043.070 ;
        RECT 2316.530 3041.890 2317.710 3043.070 ;
        RECT 2314.930 3040.290 2316.110 3041.470 ;
        RECT 2316.530 3040.290 2317.710 3041.470 ;
        RECT 2314.930 2861.890 2316.110 2863.070 ;
        RECT 2316.530 2861.890 2317.710 2863.070 ;
        RECT 2314.930 2860.290 2316.110 2861.470 ;
        RECT 2316.530 2860.290 2317.710 2861.470 ;
        RECT 2314.930 2681.890 2316.110 2683.070 ;
        RECT 2316.530 2681.890 2317.710 2683.070 ;
        RECT 2314.930 2680.290 2316.110 2681.470 ;
        RECT 2316.530 2680.290 2317.710 2681.470 ;
        RECT 2314.930 2501.890 2316.110 2503.070 ;
        RECT 2316.530 2501.890 2317.710 2503.070 ;
        RECT 2314.930 2500.290 2316.110 2501.470 ;
        RECT 2316.530 2500.290 2317.710 2501.470 ;
        RECT 2314.930 2321.890 2316.110 2323.070 ;
        RECT 2316.530 2321.890 2317.710 2323.070 ;
        RECT 2314.930 2320.290 2316.110 2321.470 ;
        RECT 2316.530 2320.290 2317.710 2321.470 ;
        RECT 2314.930 2141.890 2316.110 2143.070 ;
        RECT 2316.530 2141.890 2317.710 2143.070 ;
        RECT 2314.930 2140.290 2316.110 2141.470 ;
        RECT 2316.530 2140.290 2317.710 2141.470 ;
        RECT 2314.930 1961.890 2316.110 1963.070 ;
        RECT 2316.530 1961.890 2317.710 1963.070 ;
        RECT 2314.930 1960.290 2316.110 1961.470 ;
        RECT 2316.530 1960.290 2317.710 1961.470 ;
        RECT 2314.930 1781.890 2316.110 1783.070 ;
        RECT 2316.530 1781.890 2317.710 1783.070 ;
        RECT 2314.930 1780.290 2316.110 1781.470 ;
        RECT 2316.530 1780.290 2317.710 1781.470 ;
        RECT 2314.930 1601.890 2316.110 1603.070 ;
        RECT 2316.530 1601.890 2317.710 1603.070 ;
        RECT 2314.930 1600.290 2316.110 1601.470 ;
        RECT 2316.530 1600.290 2317.710 1601.470 ;
        RECT 2314.930 1421.890 2316.110 1423.070 ;
        RECT 2316.530 1421.890 2317.710 1423.070 ;
        RECT 2314.930 1420.290 2316.110 1421.470 ;
        RECT 2316.530 1420.290 2317.710 1421.470 ;
        RECT 2314.930 1241.890 2316.110 1243.070 ;
        RECT 2316.530 1241.890 2317.710 1243.070 ;
        RECT 2314.930 1240.290 2316.110 1241.470 ;
        RECT 2316.530 1240.290 2317.710 1241.470 ;
        RECT 2314.930 1061.890 2316.110 1063.070 ;
        RECT 2316.530 1061.890 2317.710 1063.070 ;
        RECT 2314.930 1060.290 2316.110 1061.470 ;
        RECT 2316.530 1060.290 2317.710 1061.470 ;
        RECT 2314.930 881.890 2316.110 883.070 ;
        RECT 2316.530 881.890 2317.710 883.070 ;
        RECT 2314.930 880.290 2316.110 881.470 ;
        RECT 2316.530 880.290 2317.710 881.470 ;
        RECT 2314.930 701.890 2316.110 703.070 ;
        RECT 2316.530 701.890 2317.710 703.070 ;
        RECT 2314.930 700.290 2316.110 701.470 ;
        RECT 2316.530 700.290 2317.710 701.470 ;
        RECT 2314.930 521.890 2316.110 523.070 ;
        RECT 2316.530 521.890 2317.710 523.070 ;
        RECT 2314.930 520.290 2316.110 521.470 ;
        RECT 2316.530 520.290 2317.710 521.470 ;
        RECT 2314.930 341.890 2316.110 343.070 ;
        RECT 2316.530 341.890 2317.710 343.070 ;
        RECT 2314.930 340.290 2316.110 341.470 ;
        RECT 2316.530 340.290 2317.710 341.470 ;
        RECT 2314.930 161.890 2316.110 163.070 ;
        RECT 2316.530 161.890 2317.710 163.070 ;
        RECT 2314.930 160.290 2316.110 161.470 ;
        RECT 2316.530 160.290 2317.710 161.470 ;
        RECT 2314.930 -36.510 2316.110 -35.330 ;
        RECT 2316.530 -36.510 2317.710 -35.330 ;
        RECT 2314.930 -38.110 2316.110 -36.930 ;
        RECT 2316.530 -38.110 2317.710 -36.930 ;
        RECT 2494.930 3556.610 2496.110 3557.790 ;
        RECT 2496.530 3556.610 2497.710 3557.790 ;
        RECT 2494.930 3555.010 2496.110 3556.190 ;
        RECT 2496.530 3555.010 2497.710 3556.190 ;
        RECT 2494.930 3401.890 2496.110 3403.070 ;
        RECT 2496.530 3401.890 2497.710 3403.070 ;
        RECT 2494.930 3400.290 2496.110 3401.470 ;
        RECT 2496.530 3400.290 2497.710 3401.470 ;
        RECT 2494.930 3221.890 2496.110 3223.070 ;
        RECT 2496.530 3221.890 2497.710 3223.070 ;
        RECT 2494.930 3220.290 2496.110 3221.470 ;
        RECT 2496.530 3220.290 2497.710 3221.470 ;
        RECT 2494.930 3041.890 2496.110 3043.070 ;
        RECT 2496.530 3041.890 2497.710 3043.070 ;
        RECT 2494.930 3040.290 2496.110 3041.470 ;
        RECT 2496.530 3040.290 2497.710 3041.470 ;
        RECT 2494.930 2861.890 2496.110 2863.070 ;
        RECT 2496.530 2861.890 2497.710 2863.070 ;
        RECT 2494.930 2860.290 2496.110 2861.470 ;
        RECT 2496.530 2860.290 2497.710 2861.470 ;
        RECT 2494.930 2681.890 2496.110 2683.070 ;
        RECT 2496.530 2681.890 2497.710 2683.070 ;
        RECT 2494.930 2680.290 2496.110 2681.470 ;
        RECT 2496.530 2680.290 2497.710 2681.470 ;
        RECT 2494.930 2501.890 2496.110 2503.070 ;
        RECT 2496.530 2501.890 2497.710 2503.070 ;
        RECT 2494.930 2500.290 2496.110 2501.470 ;
        RECT 2496.530 2500.290 2497.710 2501.470 ;
        RECT 2494.930 2321.890 2496.110 2323.070 ;
        RECT 2496.530 2321.890 2497.710 2323.070 ;
        RECT 2494.930 2320.290 2496.110 2321.470 ;
        RECT 2496.530 2320.290 2497.710 2321.470 ;
        RECT 2494.930 2141.890 2496.110 2143.070 ;
        RECT 2496.530 2141.890 2497.710 2143.070 ;
        RECT 2494.930 2140.290 2496.110 2141.470 ;
        RECT 2496.530 2140.290 2497.710 2141.470 ;
        RECT 2494.930 1961.890 2496.110 1963.070 ;
        RECT 2496.530 1961.890 2497.710 1963.070 ;
        RECT 2494.930 1960.290 2496.110 1961.470 ;
        RECT 2496.530 1960.290 2497.710 1961.470 ;
        RECT 2494.930 1781.890 2496.110 1783.070 ;
        RECT 2496.530 1781.890 2497.710 1783.070 ;
        RECT 2494.930 1780.290 2496.110 1781.470 ;
        RECT 2496.530 1780.290 2497.710 1781.470 ;
        RECT 2494.930 1601.890 2496.110 1603.070 ;
        RECT 2496.530 1601.890 2497.710 1603.070 ;
        RECT 2494.930 1600.290 2496.110 1601.470 ;
        RECT 2496.530 1600.290 2497.710 1601.470 ;
        RECT 2494.930 1421.890 2496.110 1423.070 ;
        RECT 2496.530 1421.890 2497.710 1423.070 ;
        RECT 2494.930 1420.290 2496.110 1421.470 ;
        RECT 2496.530 1420.290 2497.710 1421.470 ;
        RECT 2494.930 1241.890 2496.110 1243.070 ;
        RECT 2496.530 1241.890 2497.710 1243.070 ;
        RECT 2494.930 1240.290 2496.110 1241.470 ;
        RECT 2496.530 1240.290 2497.710 1241.470 ;
        RECT 2494.930 1061.890 2496.110 1063.070 ;
        RECT 2496.530 1061.890 2497.710 1063.070 ;
        RECT 2494.930 1060.290 2496.110 1061.470 ;
        RECT 2496.530 1060.290 2497.710 1061.470 ;
        RECT 2494.930 881.890 2496.110 883.070 ;
        RECT 2496.530 881.890 2497.710 883.070 ;
        RECT 2494.930 880.290 2496.110 881.470 ;
        RECT 2496.530 880.290 2497.710 881.470 ;
        RECT 2494.930 701.890 2496.110 703.070 ;
        RECT 2496.530 701.890 2497.710 703.070 ;
        RECT 2494.930 700.290 2496.110 701.470 ;
        RECT 2496.530 700.290 2497.710 701.470 ;
        RECT 2494.930 521.890 2496.110 523.070 ;
        RECT 2496.530 521.890 2497.710 523.070 ;
        RECT 2494.930 520.290 2496.110 521.470 ;
        RECT 2496.530 520.290 2497.710 521.470 ;
        RECT 2494.930 341.890 2496.110 343.070 ;
        RECT 2496.530 341.890 2497.710 343.070 ;
        RECT 2494.930 340.290 2496.110 341.470 ;
        RECT 2496.530 340.290 2497.710 341.470 ;
        RECT 2494.930 161.890 2496.110 163.070 ;
        RECT 2496.530 161.890 2497.710 163.070 ;
        RECT 2494.930 160.290 2496.110 161.470 ;
        RECT 2496.530 160.290 2497.710 161.470 ;
        RECT 2494.930 -36.510 2496.110 -35.330 ;
        RECT 2496.530 -36.510 2497.710 -35.330 ;
        RECT 2494.930 -38.110 2496.110 -36.930 ;
        RECT 2496.530 -38.110 2497.710 -36.930 ;
        RECT 2674.930 3556.610 2676.110 3557.790 ;
        RECT 2676.530 3556.610 2677.710 3557.790 ;
        RECT 2674.930 3555.010 2676.110 3556.190 ;
        RECT 2676.530 3555.010 2677.710 3556.190 ;
        RECT 2674.930 3401.890 2676.110 3403.070 ;
        RECT 2676.530 3401.890 2677.710 3403.070 ;
        RECT 2674.930 3400.290 2676.110 3401.470 ;
        RECT 2676.530 3400.290 2677.710 3401.470 ;
        RECT 2674.930 3221.890 2676.110 3223.070 ;
        RECT 2676.530 3221.890 2677.710 3223.070 ;
        RECT 2674.930 3220.290 2676.110 3221.470 ;
        RECT 2676.530 3220.290 2677.710 3221.470 ;
        RECT 2674.930 3041.890 2676.110 3043.070 ;
        RECT 2676.530 3041.890 2677.710 3043.070 ;
        RECT 2674.930 3040.290 2676.110 3041.470 ;
        RECT 2676.530 3040.290 2677.710 3041.470 ;
        RECT 2674.930 2861.890 2676.110 2863.070 ;
        RECT 2676.530 2861.890 2677.710 2863.070 ;
        RECT 2674.930 2860.290 2676.110 2861.470 ;
        RECT 2676.530 2860.290 2677.710 2861.470 ;
        RECT 2674.930 2681.890 2676.110 2683.070 ;
        RECT 2676.530 2681.890 2677.710 2683.070 ;
        RECT 2674.930 2680.290 2676.110 2681.470 ;
        RECT 2676.530 2680.290 2677.710 2681.470 ;
        RECT 2674.930 2501.890 2676.110 2503.070 ;
        RECT 2676.530 2501.890 2677.710 2503.070 ;
        RECT 2674.930 2500.290 2676.110 2501.470 ;
        RECT 2676.530 2500.290 2677.710 2501.470 ;
        RECT 2674.930 2321.890 2676.110 2323.070 ;
        RECT 2676.530 2321.890 2677.710 2323.070 ;
        RECT 2674.930 2320.290 2676.110 2321.470 ;
        RECT 2676.530 2320.290 2677.710 2321.470 ;
        RECT 2674.930 2141.890 2676.110 2143.070 ;
        RECT 2676.530 2141.890 2677.710 2143.070 ;
        RECT 2674.930 2140.290 2676.110 2141.470 ;
        RECT 2676.530 2140.290 2677.710 2141.470 ;
        RECT 2674.930 1961.890 2676.110 1963.070 ;
        RECT 2676.530 1961.890 2677.710 1963.070 ;
        RECT 2674.930 1960.290 2676.110 1961.470 ;
        RECT 2676.530 1960.290 2677.710 1961.470 ;
        RECT 2674.930 1781.890 2676.110 1783.070 ;
        RECT 2676.530 1781.890 2677.710 1783.070 ;
        RECT 2674.930 1780.290 2676.110 1781.470 ;
        RECT 2676.530 1780.290 2677.710 1781.470 ;
        RECT 2674.930 1601.890 2676.110 1603.070 ;
        RECT 2676.530 1601.890 2677.710 1603.070 ;
        RECT 2674.930 1600.290 2676.110 1601.470 ;
        RECT 2676.530 1600.290 2677.710 1601.470 ;
        RECT 2674.930 1421.890 2676.110 1423.070 ;
        RECT 2676.530 1421.890 2677.710 1423.070 ;
        RECT 2674.930 1420.290 2676.110 1421.470 ;
        RECT 2676.530 1420.290 2677.710 1421.470 ;
        RECT 2674.930 1241.890 2676.110 1243.070 ;
        RECT 2676.530 1241.890 2677.710 1243.070 ;
        RECT 2674.930 1240.290 2676.110 1241.470 ;
        RECT 2676.530 1240.290 2677.710 1241.470 ;
        RECT 2674.930 1061.890 2676.110 1063.070 ;
        RECT 2676.530 1061.890 2677.710 1063.070 ;
        RECT 2674.930 1060.290 2676.110 1061.470 ;
        RECT 2676.530 1060.290 2677.710 1061.470 ;
        RECT 2674.930 881.890 2676.110 883.070 ;
        RECT 2676.530 881.890 2677.710 883.070 ;
        RECT 2674.930 880.290 2676.110 881.470 ;
        RECT 2676.530 880.290 2677.710 881.470 ;
        RECT 2674.930 701.890 2676.110 703.070 ;
        RECT 2676.530 701.890 2677.710 703.070 ;
        RECT 2674.930 700.290 2676.110 701.470 ;
        RECT 2676.530 700.290 2677.710 701.470 ;
        RECT 2674.930 521.890 2676.110 523.070 ;
        RECT 2676.530 521.890 2677.710 523.070 ;
        RECT 2674.930 520.290 2676.110 521.470 ;
        RECT 2676.530 520.290 2677.710 521.470 ;
        RECT 2674.930 341.890 2676.110 343.070 ;
        RECT 2676.530 341.890 2677.710 343.070 ;
        RECT 2674.930 340.290 2676.110 341.470 ;
        RECT 2676.530 340.290 2677.710 341.470 ;
        RECT 2674.930 161.890 2676.110 163.070 ;
        RECT 2676.530 161.890 2677.710 163.070 ;
        RECT 2674.930 160.290 2676.110 161.470 ;
        RECT 2676.530 160.290 2677.710 161.470 ;
        RECT 2674.930 -36.510 2676.110 -35.330 ;
        RECT 2676.530 -36.510 2677.710 -35.330 ;
        RECT 2674.930 -38.110 2676.110 -36.930 ;
        RECT 2676.530 -38.110 2677.710 -36.930 ;
        RECT 2854.930 3556.610 2856.110 3557.790 ;
        RECT 2856.530 3556.610 2857.710 3557.790 ;
        RECT 2854.930 3555.010 2856.110 3556.190 ;
        RECT 2856.530 3555.010 2857.710 3556.190 ;
        RECT 2854.930 3401.890 2856.110 3403.070 ;
        RECT 2856.530 3401.890 2857.710 3403.070 ;
        RECT 2854.930 3400.290 2856.110 3401.470 ;
        RECT 2856.530 3400.290 2857.710 3401.470 ;
        RECT 2854.930 3221.890 2856.110 3223.070 ;
        RECT 2856.530 3221.890 2857.710 3223.070 ;
        RECT 2854.930 3220.290 2856.110 3221.470 ;
        RECT 2856.530 3220.290 2857.710 3221.470 ;
        RECT 2854.930 3041.890 2856.110 3043.070 ;
        RECT 2856.530 3041.890 2857.710 3043.070 ;
        RECT 2854.930 3040.290 2856.110 3041.470 ;
        RECT 2856.530 3040.290 2857.710 3041.470 ;
        RECT 2854.930 2861.890 2856.110 2863.070 ;
        RECT 2856.530 2861.890 2857.710 2863.070 ;
        RECT 2854.930 2860.290 2856.110 2861.470 ;
        RECT 2856.530 2860.290 2857.710 2861.470 ;
        RECT 2854.930 2681.890 2856.110 2683.070 ;
        RECT 2856.530 2681.890 2857.710 2683.070 ;
        RECT 2854.930 2680.290 2856.110 2681.470 ;
        RECT 2856.530 2680.290 2857.710 2681.470 ;
        RECT 2854.930 2501.890 2856.110 2503.070 ;
        RECT 2856.530 2501.890 2857.710 2503.070 ;
        RECT 2854.930 2500.290 2856.110 2501.470 ;
        RECT 2856.530 2500.290 2857.710 2501.470 ;
        RECT 2854.930 2321.890 2856.110 2323.070 ;
        RECT 2856.530 2321.890 2857.710 2323.070 ;
        RECT 2854.930 2320.290 2856.110 2321.470 ;
        RECT 2856.530 2320.290 2857.710 2321.470 ;
        RECT 2854.930 2141.890 2856.110 2143.070 ;
        RECT 2856.530 2141.890 2857.710 2143.070 ;
        RECT 2854.930 2140.290 2856.110 2141.470 ;
        RECT 2856.530 2140.290 2857.710 2141.470 ;
        RECT 2854.930 1961.890 2856.110 1963.070 ;
        RECT 2856.530 1961.890 2857.710 1963.070 ;
        RECT 2854.930 1960.290 2856.110 1961.470 ;
        RECT 2856.530 1960.290 2857.710 1961.470 ;
        RECT 2854.930 1781.890 2856.110 1783.070 ;
        RECT 2856.530 1781.890 2857.710 1783.070 ;
        RECT 2854.930 1780.290 2856.110 1781.470 ;
        RECT 2856.530 1780.290 2857.710 1781.470 ;
        RECT 2854.930 1601.890 2856.110 1603.070 ;
        RECT 2856.530 1601.890 2857.710 1603.070 ;
        RECT 2854.930 1600.290 2856.110 1601.470 ;
        RECT 2856.530 1600.290 2857.710 1601.470 ;
        RECT 2854.930 1421.890 2856.110 1423.070 ;
        RECT 2856.530 1421.890 2857.710 1423.070 ;
        RECT 2854.930 1420.290 2856.110 1421.470 ;
        RECT 2856.530 1420.290 2857.710 1421.470 ;
        RECT 2854.930 1241.890 2856.110 1243.070 ;
        RECT 2856.530 1241.890 2857.710 1243.070 ;
        RECT 2854.930 1240.290 2856.110 1241.470 ;
        RECT 2856.530 1240.290 2857.710 1241.470 ;
        RECT 2854.930 1061.890 2856.110 1063.070 ;
        RECT 2856.530 1061.890 2857.710 1063.070 ;
        RECT 2854.930 1060.290 2856.110 1061.470 ;
        RECT 2856.530 1060.290 2857.710 1061.470 ;
        RECT 2854.930 881.890 2856.110 883.070 ;
        RECT 2856.530 881.890 2857.710 883.070 ;
        RECT 2854.930 880.290 2856.110 881.470 ;
        RECT 2856.530 880.290 2857.710 881.470 ;
        RECT 2854.930 701.890 2856.110 703.070 ;
        RECT 2856.530 701.890 2857.710 703.070 ;
        RECT 2854.930 700.290 2856.110 701.470 ;
        RECT 2856.530 700.290 2857.710 701.470 ;
        RECT 2854.930 521.890 2856.110 523.070 ;
        RECT 2856.530 521.890 2857.710 523.070 ;
        RECT 2854.930 520.290 2856.110 521.470 ;
        RECT 2856.530 520.290 2857.710 521.470 ;
        RECT 2854.930 341.890 2856.110 343.070 ;
        RECT 2856.530 341.890 2857.710 343.070 ;
        RECT 2854.930 340.290 2856.110 341.470 ;
        RECT 2856.530 340.290 2857.710 341.470 ;
        RECT 2854.930 161.890 2856.110 163.070 ;
        RECT 2856.530 161.890 2857.710 163.070 ;
        RECT 2854.930 160.290 2856.110 161.470 ;
        RECT 2856.530 160.290 2857.710 161.470 ;
        RECT 2854.930 -36.510 2856.110 -35.330 ;
        RECT 2856.530 -36.510 2857.710 -35.330 ;
        RECT 2854.930 -38.110 2856.110 -36.930 ;
        RECT 2856.530 -38.110 2857.710 -36.930 ;
        RECT 2960.310 3556.610 2961.490 3557.790 ;
        RECT 2961.910 3556.610 2963.090 3557.790 ;
        RECT 2960.310 3555.010 2961.490 3556.190 ;
        RECT 2961.910 3555.010 2963.090 3556.190 ;
        RECT 2960.310 3401.890 2961.490 3403.070 ;
        RECT 2961.910 3401.890 2963.090 3403.070 ;
        RECT 2960.310 3400.290 2961.490 3401.470 ;
        RECT 2961.910 3400.290 2963.090 3401.470 ;
        RECT 2960.310 3221.890 2961.490 3223.070 ;
        RECT 2961.910 3221.890 2963.090 3223.070 ;
        RECT 2960.310 3220.290 2961.490 3221.470 ;
        RECT 2961.910 3220.290 2963.090 3221.470 ;
        RECT 2960.310 3041.890 2961.490 3043.070 ;
        RECT 2961.910 3041.890 2963.090 3043.070 ;
        RECT 2960.310 3040.290 2961.490 3041.470 ;
        RECT 2961.910 3040.290 2963.090 3041.470 ;
        RECT 2960.310 2861.890 2961.490 2863.070 ;
        RECT 2961.910 2861.890 2963.090 2863.070 ;
        RECT 2960.310 2860.290 2961.490 2861.470 ;
        RECT 2961.910 2860.290 2963.090 2861.470 ;
        RECT 2960.310 2681.890 2961.490 2683.070 ;
        RECT 2961.910 2681.890 2963.090 2683.070 ;
        RECT 2960.310 2680.290 2961.490 2681.470 ;
        RECT 2961.910 2680.290 2963.090 2681.470 ;
        RECT 2960.310 2501.890 2961.490 2503.070 ;
        RECT 2961.910 2501.890 2963.090 2503.070 ;
        RECT 2960.310 2500.290 2961.490 2501.470 ;
        RECT 2961.910 2500.290 2963.090 2501.470 ;
        RECT 2960.310 2321.890 2961.490 2323.070 ;
        RECT 2961.910 2321.890 2963.090 2323.070 ;
        RECT 2960.310 2320.290 2961.490 2321.470 ;
        RECT 2961.910 2320.290 2963.090 2321.470 ;
        RECT 2960.310 2141.890 2961.490 2143.070 ;
        RECT 2961.910 2141.890 2963.090 2143.070 ;
        RECT 2960.310 2140.290 2961.490 2141.470 ;
        RECT 2961.910 2140.290 2963.090 2141.470 ;
        RECT 2960.310 1961.890 2961.490 1963.070 ;
        RECT 2961.910 1961.890 2963.090 1963.070 ;
        RECT 2960.310 1960.290 2961.490 1961.470 ;
        RECT 2961.910 1960.290 2963.090 1961.470 ;
        RECT 2960.310 1781.890 2961.490 1783.070 ;
        RECT 2961.910 1781.890 2963.090 1783.070 ;
        RECT 2960.310 1780.290 2961.490 1781.470 ;
        RECT 2961.910 1780.290 2963.090 1781.470 ;
        RECT 2960.310 1601.890 2961.490 1603.070 ;
        RECT 2961.910 1601.890 2963.090 1603.070 ;
        RECT 2960.310 1600.290 2961.490 1601.470 ;
        RECT 2961.910 1600.290 2963.090 1601.470 ;
        RECT 2960.310 1421.890 2961.490 1423.070 ;
        RECT 2961.910 1421.890 2963.090 1423.070 ;
        RECT 2960.310 1420.290 2961.490 1421.470 ;
        RECT 2961.910 1420.290 2963.090 1421.470 ;
        RECT 2960.310 1241.890 2961.490 1243.070 ;
        RECT 2961.910 1241.890 2963.090 1243.070 ;
        RECT 2960.310 1240.290 2961.490 1241.470 ;
        RECT 2961.910 1240.290 2963.090 1241.470 ;
        RECT 2960.310 1061.890 2961.490 1063.070 ;
        RECT 2961.910 1061.890 2963.090 1063.070 ;
        RECT 2960.310 1060.290 2961.490 1061.470 ;
        RECT 2961.910 1060.290 2963.090 1061.470 ;
        RECT 2960.310 881.890 2961.490 883.070 ;
        RECT 2961.910 881.890 2963.090 883.070 ;
        RECT 2960.310 880.290 2961.490 881.470 ;
        RECT 2961.910 880.290 2963.090 881.470 ;
        RECT 2960.310 701.890 2961.490 703.070 ;
        RECT 2961.910 701.890 2963.090 703.070 ;
        RECT 2960.310 700.290 2961.490 701.470 ;
        RECT 2961.910 700.290 2963.090 701.470 ;
        RECT 2960.310 521.890 2961.490 523.070 ;
        RECT 2961.910 521.890 2963.090 523.070 ;
        RECT 2960.310 520.290 2961.490 521.470 ;
        RECT 2961.910 520.290 2963.090 521.470 ;
        RECT 2960.310 341.890 2961.490 343.070 ;
        RECT 2961.910 341.890 2963.090 343.070 ;
        RECT 2960.310 340.290 2961.490 341.470 ;
        RECT 2961.910 340.290 2963.090 341.470 ;
        RECT 2960.310 161.890 2961.490 163.070 ;
        RECT 2961.910 161.890 2963.090 163.070 ;
        RECT 2960.310 160.290 2961.490 161.470 ;
        RECT 2961.910 160.290 2963.090 161.470 ;
        RECT 2960.310 -36.510 2961.490 -35.330 ;
        RECT 2961.910 -36.510 2963.090 -35.330 ;
        RECT 2960.310 -38.110 2961.490 -36.930 ;
        RECT 2961.910 -38.110 2963.090 -36.930 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
        RECT -43.630 880.130 2963.250 883.230 ;
        RECT -43.630 700.130 2963.250 703.230 ;
        RECT -43.630 520.130 2963.250 523.230 ;
        RECT -43.630 340.130 2963.250 343.230 ;
        RECT -43.630 160.130 2963.250 163.230 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
        RECT 278.970 1010.000 282.070 3529.150 ;
        RECT 458.970 1010.000 462.070 3529.150 ;
        RECT 638.970 1010.000 642.070 3529.150 ;
        RECT 818.970 1010.000 822.070 3529.150 ;
        RECT 998.970 1010.000 1002.070 3529.150 ;
        RECT 297.840 410.640 299.440 987.760 ;
        RECT 451.440 410.640 453.040 987.760 ;
        RECT 605.040 410.640 606.640 987.760 ;
        RECT 758.640 410.640 760.240 987.760 ;
        RECT 912.240 410.640 913.840 987.760 ;
        RECT 1065.840 410.640 1067.440 987.760 ;
        RECT 278.970 -9.470 282.070 390.000 ;
        RECT 458.970 -9.470 462.070 390.000 ;
        RECT 638.970 -9.470 642.070 390.000 ;
        RECT 818.970 -9.470 822.070 390.000 ;
        RECT 998.970 -9.470 1002.070 390.000 ;
        RECT 1178.970 -9.470 1182.070 3529.150 ;
        RECT 1358.970 -9.470 1362.070 3529.150 ;
        RECT 1538.970 -9.470 1542.070 3529.150 ;
        RECT 1718.970 -9.470 1722.070 3529.150 ;
        RECT 1898.970 -9.470 1902.070 3529.150 ;
        RECT 2078.970 -9.470 2082.070 3529.150 ;
        RECT 2258.970 -9.470 2262.070 3529.150 ;
        RECT 2438.970 -9.470 2442.070 3529.150 ;
        RECT 2618.970 -9.470 2622.070 3529.150 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER via4 ;
        RECT -14.670 3527.810 -13.490 3528.990 ;
        RECT -13.070 3527.810 -11.890 3528.990 ;
        RECT -14.670 3526.210 -13.490 3527.390 ;
        RECT -13.070 3526.210 -11.890 3527.390 ;
        RECT -14.670 3346.090 -13.490 3347.270 ;
        RECT -13.070 3346.090 -11.890 3347.270 ;
        RECT -14.670 3344.490 -13.490 3345.670 ;
        RECT -13.070 3344.490 -11.890 3345.670 ;
        RECT -14.670 3166.090 -13.490 3167.270 ;
        RECT -13.070 3166.090 -11.890 3167.270 ;
        RECT -14.670 3164.490 -13.490 3165.670 ;
        RECT -13.070 3164.490 -11.890 3165.670 ;
        RECT -14.670 2986.090 -13.490 2987.270 ;
        RECT -13.070 2986.090 -11.890 2987.270 ;
        RECT -14.670 2984.490 -13.490 2985.670 ;
        RECT -13.070 2984.490 -11.890 2985.670 ;
        RECT -14.670 2806.090 -13.490 2807.270 ;
        RECT -13.070 2806.090 -11.890 2807.270 ;
        RECT -14.670 2804.490 -13.490 2805.670 ;
        RECT -13.070 2804.490 -11.890 2805.670 ;
        RECT -14.670 2626.090 -13.490 2627.270 ;
        RECT -13.070 2626.090 -11.890 2627.270 ;
        RECT -14.670 2624.490 -13.490 2625.670 ;
        RECT -13.070 2624.490 -11.890 2625.670 ;
        RECT -14.670 2446.090 -13.490 2447.270 ;
        RECT -13.070 2446.090 -11.890 2447.270 ;
        RECT -14.670 2444.490 -13.490 2445.670 ;
        RECT -13.070 2444.490 -11.890 2445.670 ;
        RECT -14.670 2266.090 -13.490 2267.270 ;
        RECT -13.070 2266.090 -11.890 2267.270 ;
        RECT -14.670 2264.490 -13.490 2265.670 ;
        RECT -13.070 2264.490 -11.890 2265.670 ;
        RECT -14.670 2086.090 -13.490 2087.270 ;
        RECT -13.070 2086.090 -11.890 2087.270 ;
        RECT -14.670 2084.490 -13.490 2085.670 ;
        RECT -13.070 2084.490 -11.890 2085.670 ;
        RECT -14.670 1906.090 -13.490 1907.270 ;
        RECT -13.070 1906.090 -11.890 1907.270 ;
        RECT -14.670 1904.490 -13.490 1905.670 ;
        RECT -13.070 1904.490 -11.890 1905.670 ;
        RECT -14.670 1726.090 -13.490 1727.270 ;
        RECT -13.070 1726.090 -11.890 1727.270 ;
        RECT -14.670 1724.490 -13.490 1725.670 ;
        RECT -13.070 1724.490 -11.890 1725.670 ;
        RECT -14.670 1546.090 -13.490 1547.270 ;
        RECT -13.070 1546.090 -11.890 1547.270 ;
        RECT -14.670 1544.490 -13.490 1545.670 ;
        RECT -13.070 1544.490 -11.890 1545.670 ;
        RECT -14.670 1366.090 -13.490 1367.270 ;
        RECT -13.070 1366.090 -11.890 1367.270 ;
        RECT -14.670 1364.490 -13.490 1365.670 ;
        RECT -13.070 1364.490 -11.890 1365.670 ;
        RECT -14.670 1186.090 -13.490 1187.270 ;
        RECT -13.070 1186.090 -11.890 1187.270 ;
        RECT -14.670 1184.490 -13.490 1185.670 ;
        RECT -13.070 1184.490 -11.890 1185.670 ;
        RECT -14.670 1006.090 -13.490 1007.270 ;
        RECT -13.070 1006.090 -11.890 1007.270 ;
        RECT -14.670 1004.490 -13.490 1005.670 ;
        RECT -13.070 1004.490 -11.890 1005.670 ;
        RECT -14.670 826.090 -13.490 827.270 ;
        RECT -13.070 826.090 -11.890 827.270 ;
        RECT -14.670 824.490 -13.490 825.670 ;
        RECT -13.070 824.490 -11.890 825.670 ;
        RECT -14.670 646.090 -13.490 647.270 ;
        RECT -13.070 646.090 -11.890 647.270 ;
        RECT -14.670 644.490 -13.490 645.670 ;
        RECT -13.070 644.490 -11.890 645.670 ;
        RECT -14.670 466.090 -13.490 467.270 ;
        RECT -13.070 466.090 -11.890 467.270 ;
        RECT -14.670 464.490 -13.490 465.670 ;
        RECT -13.070 464.490 -11.890 465.670 ;
        RECT -14.670 286.090 -13.490 287.270 ;
        RECT -13.070 286.090 -11.890 287.270 ;
        RECT -14.670 284.490 -13.490 285.670 ;
        RECT -13.070 284.490 -11.890 285.670 ;
        RECT -14.670 106.090 -13.490 107.270 ;
        RECT -13.070 106.090 -11.890 107.270 ;
        RECT -14.670 104.490 -13.490 105.670 ;
        RECT -13.070 104.490 -11.890 105.670 ;
        RECT -14.670 -7.710 -13.490 -6.530 ;
        RECT -13.070 -7.710 -11.890 -6.530 ;
        RECT -14.670 -9.310 -13.490 -8.130 ;
        RECT -13.070 -9.310 -11.890 -8.130 ;
        RECT 99.130 3527.810 100.310 3528.990 ;
        RECT 100.730 3527.810 101.910 3528.990 ;
        RECT 99.130 3526.210 100.310 3527.390 ;
        RECT 100.730 3526.210 101.910 3527.390 ;
        RECT 99.130 3346.090 100.310 3347.270 ;
        RECT 100.730 3346.090 101.910 3347.270 ;
        RECT 99.130 3344.490 100.310 3345.670 ;
        RECT 100.730 3344.490 101.910 3345.670 ;
        RECT 99.130 3166.090 100.310 3167.270 ;
        RECT 100.730 3166.090 101.910 3167.270 ;
        RECT 99.130 3164.490 100.310 3165.670 ;
        RECT 100.730 3164.490 101.910 3165.670 ;
        RECT 99.130 2986.090 100.310 2987.270 ;
        RECT 100.730 2986.090 101.910 2987.270 ;
        RECT 99.130 2984.490 100.310 2985.670 ;
        RECT 100.730 2984.490 101.910 2985.670 ;
        RECT 99.130 2806.090 100.310 2807.270 ;
        RECT 100.730 2806.090 101.910 2807.270 ;
        RECT 99.130 2804.490 100.310 2805.670 ;
        RECT 100.730 2804.490 101.910 2805.670 ;
        RECT 99.130 2626.090 100.310 2627.270 ;
        RECT 100.730 2626.090 101.910 2627.270 ;
        RECT 99.130 2624.490 100.310 2625.670 ;
        RECT 100.730 2624.490 101.910 2625.670 ;
        RECT 99.130 2446.090 100.310 2447.270 ;
        RECT 100.730 2446.090 101.910 2447.270 ;
        RECT 99.130 2444.490 100.310 2445.670 ;
        RECT 100.730 2444.490 101.910 2445.670 ;
        RECT 99.130 2266.090 100.310 2267.270 ;
        RECT 100.730 2266.090 101.910 2267.270 ;
        RECT 99.130 2264.490 100.310 2265.670 ;
        RECT 100.730 2264.490 101.910 2265.670 ;
        RECT 99.130 2086.090 100.310 2087.270 ;
        RECT 100.730 2086.090 101.910 2087.270 ;
        RECT 99.130 2084.490 100.310 2085.670 ;
        RECT 100.730 2084.490 101.910 2085.670 ;
        RECT 99.130 1906.090 100.310 1907.270 ;
        RECT 100.730 1906.090 101.910 1907.270 ;
        RECT 99.130 1904.490 100.310 1905.670 ;
        RECT 100.730 1904.490 101.910 1905.670 ;
        RECT 99.130 1726.090 100.310 1727.270 ;
        RECT 100.730 1726.090 101.910 1727.270 ;
        RECT 99.130 1724.490 100.310 1725.670 ;
        RECT 100.730 1724.490 101.910 1725.670 ;
        RECT 99.130 1546.090 100.310 1547.270 ;
        RECT 100.730 1546.090 101.910 1547.270 ;
        RECT 99.130 1544.490 100.310 1545.670 ;
        RECT 100.730 1544.490 101.910 1545.670 ;
        RECT 99.130 1366.090 100.310 1367.270 ;
        RECT 100.730 1366.090 101.910 1367.270 ;
        RECT 99.130 1364.490 100.310 1365.670 ;
        RECT 100.730 1364.490 101.910 1365.670 ;
        RECT 99.130 1186.090 100.310 1187.270 ;
        RECT 100.730 1186.090 101.910 1187.270 ;
        RECT 99.130 1184.490 100.310 1185.670 ;
        RECT 100.730 1184.490 101.910 1185.670 ;
        RECT 279.130 3527.810 280.310 3528.990 ;
        RECT 280.730 3527.810 281.910 3528.990 ;
        RECT 279.130 3526.210 280.310 3527.390 ;
        RECT 280.730 3526.210 281.910 3527.390 ;
        RECT 279.130 3346.090 280.310 3347.270 ;
        RECT 280.730 3346.090 281.910 3347.270 ;
        RECT 279.130 3344.490 280.310 3345.670 ;
        RECT 280.730 3344.490 281.910 3345.670 ;
        RECT 279.130 3166.090 280.310 3167.270 ;
        RECT 280.730 3166.090 281.910 3167.270 ;
        RECT 279.130 3164.490 280.310 3165.670 ;
        RECT 280.730 3164.490 281.910 3165.670 ;
        RECT 279.130 2986.090 280.310 2987.270 ;
        RECT 280.730 2986.090 281.910 2987.270 ;
        RECT 279.130 2984.490 280.310 2985.670 ;
        RECT 280.730 2984.490 281.910 2985.670 ;
        RECT 279.130 2806.090 280.310 2807.270 ;
        RECT 280.730 2806.090 281.910 2807.270 ;
        RECT 279.130 2804.490 280.310 2805.670 ;
        RECT 280.730 2804.490 281.910 2805.670 ;
        RECT 279.130 2626.090 280.310 2627.270 ;
        RECT 280.730 2626.090 281.910 2627.270 ;
        RECT 279.130 2624.490 280.310 2625.670 ;
        RECT 280.730 2624.490 281.910 2625.670 ;
        RECT 279.130 2446.090 280.310 2447.270 ;
        RECT 280.730 2446.090 281.910 2447.270 ;
        RECT 279.130 2444.490 280.310 2445.670 ;
        RECT 280.730 2444.490 281.910 2445.670 ;
        RECT 279.130 2266.090 280.310 2267.270 ;
        RECT 280.730 2266.090 281.910 2267.270 ;
        RECT 279.130 2264.490 280.310 2265.670 ;
        RECT 280.730 2264.490 281.910 2265.670 ;
        RECT 279.130 2086.090 280.310 2087.270 ;
        RECT 280.730 2086.090 281.910 2087.270 ;
        RECT 279.130 2084.490 280.310 2085.670 ;
        RECT 280.730 2084.490 281.910 2085.670 ;
        RECT 279.130 1906.090 280.310 1907.270 ;
        RECT 280.730 1906.090 281.910 1907.270 ;
        RECT 279.130 1904.490 280.310 1905.670 ;
        RECT 280.730 1904.490 281.910 1905.670 ;
        RECT 279.130 1726.090 280.310 1727.270 ;
        RECT 280.730 1726.090 281.910 1727.270 ;
        RECT 279.130 1724.490 280.310 1725.670 ;
        RECT 280.730 1724.490 281.910 1725.670 ;
        RECT 279.130 1546.090 280.310 1547.270 ;
        RECT 280.730 1546.090 281.910 1547.270 ;
        RECT 279.130 1544.490 280.310 1545.670 ;
        RECT 280.730 1544.490 281.910 1545.670 ;
        RECT 279.130 1366.090 280.310 1367.270 ;
        RECT 280.730 1366.090 281.910 1367.270 ;
        RECT 279.130 1364.490 280.310 1365.670 ;
        RECT 280.730 1364.490 281.910 1365.670 ;
        RECT 279.130 1186.090 280.310 1187.270 ;
        RECT 280.730 1186.090 281.910 1187.270 ;
        RECT 279.130 1184.490 280.310 1185.670 ;
        RECT 280.730 1184.490 281.910 1185.670 ;
        RECT 459.130 3527.810 460.310 3528.990 ;
        RECT 460.730 3527.810 461.910 3528.990 ;
        RECT 459.130 3526.210 460.310 3527.390 ;
        RECT 460.730 3526.210 461.910 3527.390 ;
        RECT 459.130 3346.090 460.310 3347.270 ;
        RECT 460.730 3346.090 461.910 3347.270 ;
        RECT 459.130 3344.490 460.310 3345.670 ;
        RECT 460.730 3344.490 461.910 3345.670 ;
        RECT 459.130 3166.090 460.310 3167.270 ;
        RECT 460.730 3166.090 461.910 3167.270 ;
        RECT 459.130 3164.490 460.310 3165.670 ;
        RECT 460.730 3164.490 461.910 3165.670 ;
        RECT 459.130 2986.090 460.310 2987.270 ;
        RECT 460.730 2986.090 461.910 2987.270 ;
        RECT 459.130 2984.490 460.310 2985.670 ;
        RECT 460.730 2984.490 461.910 2985.670 ;
        RECT 459.130 2806.090 460.310 2807.270 ;
        RECT 460.730 2806.090 461.910 2807.270 ;
        RECT 459.130 2804.490 460.310 2805.670 ;
        RECT 460.730 2804.490 461.910 2805.670 ;
        RECT 459.130 2626.090 460.310 2627.270 ;
        RECT 460.730 2626.090 461.910 2627.270 ;
        RECT 459.130 2624.490 460.310 2625.670 ;
        RECT 460.730 2624.490 461.910 2625.670 ;
        RECT 459.130 2446.090 460.310 2447.270 ;
        RECT 460.730 2446.090 461.910 2447.270 ;
        RECT 459.130 2444.490 460.310 2445.670 ;
        RECT 460.730 2444.490 461.910 2445.670 ;
        RECT 459.130 2266.090 460.310 2267.270 ;
        RECT 460.730 2266.090 461.910 2267.270 ;
        RECT 459.130 2264.490 460.310 2265.670 ;
        RECT 460.730 2264.490 461.910 2265.670 ;
        RECT 459.130 2086.090 460.310 2087.270 ;
        RECT 460.730 2086.090 461.910 2087.270 ;
        RECT 459.130 2084.490 460.310 2085.670 ;
        RECT 460.730 2084.490 461.910 2085.670 ;
        RECT 459.130 1906.090 460.310 1907.270 ;
        RECT 460.730 1906.090 461.910 1907.270 ;
        RECT 459.130 1904.490 460.310 1905.670 ;
        RECT 460.730 1904.490 461.910 1905.670 ;
        RECT 459.130 1726.090 460.310 1727.270 ;
        RECT 460.730 1726.090 461.910 1727.270 ;
        RECT 459.130 1724.490 460.310 1725.670 ;
        RECT 460.730 1724.490 461.910 1725.670 ;
        RECT 459.130 1546.090 460.310 1547.270 ;
        RECT 460.730 1546.090 461.910 1547.270 ;
        RECT 459.130 1544.490 460.310 1545.670 ;
        RECT 460.730 1544.490 461.910 1545.670 ;
        RECT 459.130 1366.090 460.310 1367.270 ;
        RECT 460.730 1366.090 461.910 1367.270 ;
        RECT 459.130 1364.490 460.310 1365.670 ;
        RECT 460.730 1364.490 461.910 1365.670 ;
        RECT 459.130 1186.090 460.310 1187.270 ;
        RECT 460.730 1186.090 461.910 1187.270 ;
        RECT 459.130 1184.490 460.310 1185.670 ;
        RECT 460.730 1184.490 461.910 1185.670 ;
        RECT 639.130 3527.810 640.310 3528.990 ;
        RECT 640.730 3527.810 641.910 3528.990 ;
        RECT 639.130 3526.210 640.310 3527.390 ;
        RECT 640.730 3526.210 641.910 3527.390 ;
        RECT 639.130 3346.090 640.310 3347.270 ;
        RECT 640.730 3346.090 641.910 3347.270 ;
        RECT 639.130 3344.490 640.310 3345.670 ;
        RECT 640.730 3344.490 641.910 3345.670 ;
        RECT 639.130 3166.090 640.310 3167.270 ;
        RECT 640.730 3166.090 641.910 3167.270 ;
        RECT 639.130 3164.490 640.310 3165.670 ;
        RECT 640.730 3164.490 641.910 3165.670 ;
        RECT 639.130 2986.090 640.310 2987.270 ;
        RECT 640.730 2986.090 641.910 2987.270 ;
        RECT 639.130 2984.490 640.310 2985.670 ;
        RECT 640.730 2984.490 641.910 2985.670 ;
        RECT 639.130 2806.090 640.310 2807.270 ;
        RECT 640.730 2806.090 641.910 2807.270 ;
        RECT 639.130 2804.490 640.310 2805.670 ;
        RECT 640.730 2804.490 641.910 2805.670 ;
        RECT 639.130 2626.090 640.310 2627.270 ;
        RECT 640.730 2626.090 641.910 2627.270 ;
        RECT 639.130 2624.490 640.310 2625.670 ;
        RECT 640.730 2624.490 641.910 2625.670 ;
        RECT 639.130 2446.090 640.310 2447.270 ;
        RECT 640.730 2446.090 641.910 2447.270 ;
        RECT 639.130 2444.490 640.310 2445.670 ;
        RECT 640.730 2444.490 641.910 2445.670 ;
        RECT 639.130 2266.090 640.310 2267.270 ;
        RECT 640.730 2266.090 641.910 2267.270 ;
        RECT 639.130 2264.490 640.310 2265.670 ;
        RECT 640.730 2264.490 641.910 2265.670 ;
        RECT 639.130 2086.090 640.310 2087.270 ;
        RECT 640.730 2086.090 641.910 2087.270 ;
        RECT 639.130 2084.490 640.310 2085.670 ;
        RECT 640.730 2084.490 641.910 2085.670 ;
        RECT 639.130 1906.090 640.310 1907.270 ;
        RECT 640.730 1906.090 641.910 1907.270 ;
        RECT 639.130 1904.490 640.310 1905.670 ;
        RECT 640.730 1904.490 641.910 1905.670 ;
        RECT 639.130 1726.090 640.310 1727.270 ;
        RECT 640.730 1726.090 641.910 1727.270 ;
        RECT 639.130 1724.490 640.310 1725.670 ;
        RECT 640.730 1724.490 641.910 1725.670 ;
        RECT 639.130 1546.090 640.310 1547.270 ;
        RECT 640.730 1546.090 641.910 1547.270 ;
        RECT 639.130 1544.490 640.310 1545.670 ;
        RECT 640.730 1544.490 641.910 1545.670 ;
        RECT 639.130 1366.090 640.310 1367.270 ;
        RECT 640.730 1366.090 641.910 1367.270 ;
        RECT 639.130 1364.490 640.310 1365.670 ;
        RECT 640.730 1364.490 641.910 1365.670 ;
        RECT 639.130 1186.090 640.310 1187.270 ;
        RECT 640.730 1186.090 641.910 1187.270 ;
        RECT 639.130 1184.490 640.310 1185.670 ;
        RECT 640.730 1184.490 641.910 1185.670 ;
        RECT 819.130 3527.810 820.310 3528.990 ;
        RECT 820.730 3527.810 821.910 3528.990 ;
        RECT 819.130 3526.210 820.310 3527.390 ;
        RECT 820.730 3526.210 821.910 3527.390 ;
        RECT 819.130 3346.090 820.310 3347.270 ;
        RECT 820.730 3346.090 821.910 3347.270 ;
        RECT 819.130 3344.490 820.310 3345.670 ;
        RECT 820.730 3344.490 821.910 3345.670 ;
        RECT 819.130 3166.090 820.310 3167.270 ;
        RECT 820.730 3166.090 821.910 3167.270 ;
        RECT 819.130 3164.490 820.310 3165.670 ;
        RECT 820.730 3164.490 821.910 3165.670 ;
        RECT 819.130 2986.090 820.310 2987.270 ;
        RECT 820.730 2986.090 821.910 2987.270 ;
        RECT 819.130 2984.490 820.310 2985.670 ;
        RECT 820.730 2984.490 821.910 2985.670 ;
        RECT 819.130 2806.090 820.310 2807.270 ;
        RECT 820.730 2806.090 821.910 2807.270 ;
        RECT 819.130 2804.490 820.310 2805.670 ;
        RECT 820.730 2804.490 821.910 2805.670 ;
        RECT 819.130 2626.090 820.310 2627.270 ;
        RECT 820.730 2626.090 821.910 2627.270 ;
        RECT 819.130 2624.490 820.310 2625.670 ;
        RECT 820.730 2624.490 821.910 2625.670 ;
        RECT 819.130 2446.090 820.310 2447.270 ;
        RECT 820.730 2446.090 821.910 2447.270 ;
        RECT 819.130 2444.490 820.310 2445.670 ;
        RECT 820.730 2444.490 821.910 2445.670 ;
        RECT 819.130 2266.090 820.310 2267.270 ;
        RECT 820.730 2266.090 821.910 2267.270 ;
        RECT 819.130 2264.490 820.310 2265.670 ;
        RECT 820.730 2264.490 821.910 2265.670 ;
        RECT 819.130 2086.090 820.310 2087.270 ;
        RECT 820.730 2086.090 821.910 2087.270 ;
        RECT 819.130 2084.490 820.310 2085.670 ;
        RECT 820.730 2084.490 821.910 2085.670 ;
        RECT 819.130 1906.090 820.310 1907.270 ;
        RECT 820.730 1906.090 821.910 1907.270 ;
        RECT 819.130 1904.490 820.310 1905.670 ;
        RECT 820.730 1904.490 821.910 1905.670 ;
        RECT 819.130 1726.090 820.310 1727.270 ;
        RECT 820.730 1726.090 821.910 1727.270 ;
        RECT 819.130 1724.490 820.310 1725.670 ;
        RECT 820.730 1724.490 821.910 1725.670 ;
        RECT 819.130 1546.090 820.310 1547.270 ;
        RECT 820.730 1546.090 821.910 1547.270 ;
        RECT 819.130 1544.490 820.310 1545.670 ;
        RECT 820.730 1544.490 821.910 1545.670 ;
        RECT 819.130 1366.090 820.310 1367.270 ;
        RECT 820.730 1366.090 821.910 1367.270 ;
        RECT 819.130 1364.490 820.310 1365.670 ;
        RECT 820.730 1364.490 821.910 1365.670 ;
        RECT 819.130 1186.090 820.310 1187.270 ;
        RECT 820.730 1186.090 821.910 1187.270 ;
        RECT 819.130 1184.490 820.310 1185.670 ;
        RECT 820.730 1184.490 821.910 1185.670 ;
        RECT 999.130 3527.810 1000.310 3528.990 ;
        RECT 1000.730 3527.810 1001.910 3528.990 ;
        RECT 999.130 3526.210 1000.310 3527.390 ;
        RECT 1000.730 3526.210 1001.910 3527.390 ;
        RECT 999.130 3346.090 1000.310 3347.270 ;
        RECT 1000.730 3346.090 1001.910 3347.270 ;
        RECT 999.130 3344.490 1000.310 3345.670 ;
        RECT 1000.730 3344.490 1001.910 3345.670 ;
        RECT 999.130 3166.090 1000.310 3167.270 ;
        RECT 1000.730 3166.090 1001.910 3167.270 ;
        RECT 999.130 3164.490 1000.310 3165.670 ;
        RECT 1000.730 3164.490 1001.910 3165.670 ;
        RECT 999.130 2986.090 1000.310 2987.270 ;
        RECT 1000.730 2986.090 1001.910 2987.270 ;
        RECT 999.130 2984.490 1000.310 2985.670 ;
        RECT 1000.730 2984.490 1001.910 2985.670 ;
        RECT 999.130 2806.090 1000.310 2807.270 ;
        RECT 1000.730 2806.090 1001.910 2807.270 ;
        RECT 999.130 2804.490 1000.310 2805.670 ;
        RECT 1000.730 2804.490 1001.910 2805.670 ;
        RECT 999.130 2626.090 1000.310 2627.270 ;
        RECT 1000.730 2626.090 1001.910 2627.270 ;
        RECT 999.130 2624.490 1000.310 2625.670 ;
        RECT 1000.730 2624.490 1001.910 2625.670 ;
        RECT 999.130 2446.090 1000.310 2447.270 ;
        RECT 1000.730 2446.090 1001.910 2447.270 ;
        RECT 999.130 2444.490 1000.310 2445.670 ;
        RECT 1000.730 2444.490 1001.910 2445.670 ;
        RECT 999.130 2266.090 1000.310 2267.270 ;
        RECT 1000.730 2266.090 1001.910 2267.270 ;
        RECT 999.130 2264.490 1000.310 2265.670 ;
        RECT 1000.730 2264.490 1001.910 2265.670 ;
        RECT 999.130 2086.090 1000.310 2087.270 ;
        RECT 1000.730 2086.090 1001.910 2087.270 ;
        RECT 999.130 2084.490 1000.310 2085.670 ;
        RECT 1000.730 2084.490 1001.910 2085.670 ;
        RECT 999.130 1906.090 1000.310 1907.270 ;
        RECT 1000.730 1906.090 1001.910 1907.270 ;
        RECT 999.130 1904.490 1000.310 1905.670 ;
        RECT 1000.730 1904.490 1001.910 1905.670 ;
        RECT 999.130 1726.090 1000.310 1727.270 ;
        RECT 1000.730 1726.090 1001.910 1727.270 ;
        RECT 999.130 1724.490 1000.310 1725.670 ;
        RECT 1000.730 1724.490 1001.910 1725.670 ;
        RECT 999.130 1546.090 1000.310 1547.270 ;
        RECT 1000.730 1546.090 1001.910 1547.270 ;
        RECT 999.130 1544.490 1000.310 1545.670 ;
        RECT 1000.730 1544.490 1001.910 1545.670 ;
        RECT 999.130 1366.090 1000.310 1367.270 ;
        RECT 1000.730 1366.090 1001.910 1367.270 ;
        RECT 999.130 1364.490 1000.310 1365.670 ;
        RECT 1000.730 1364.490 1001.910 1365.670 ;
        RECT 999.130 1186.090 1000.310 1187.270 ;
        RECT 1000.730 1186.090 1001.910 1187.270 ;
        RECT 999.130 1184.490 1000.310 1185.670 ;
        RECT 1000.730 1184.490 1001.910 1185.670 ;
        RECT 1179.130 3527.810 1180.310 3528.990 ;
        RECT 1180.730 3527.810 1181.910 3528.990 ;
        RECT 1179.130 3526.210 1180.310 3527.390 ;
        RECT 1180.730 3526.210 1181.910 3527.390 ;
        RECT 1179.130 3346.090 1180.310 3347.270 ;
        RECT 1180.730 3346.090 1181.910 3347.270 ;
        RECT 1179.130 3344.490 1180.310 3345.670 ;
        RECT 1180.730 3344.490 1181.910 3345.670 ;
        RECT 1179.130 3166.090 1180.310 3167.270 ;
        RECT 1180.730 3166.090 1181.910 3167.270 ;
        RECT 1179.130 3164.490 1180.310 3165.670 ;
        RECT 1180.730 3164.490 1181.910 3165.670 ;
        RECT 1179.130 2986.090 1180.310 2987.270 ;
        RECT 1180.730 2986.090 1181.910 2987.270 ;
        RECT 1179.130 2984.490 1180.310 2985.670 ;
        RECT 1180.730 2984.490 1181.910 2985.670 ;
        RECT 1179.130 2806.090 1180.310 2807.270 ;
        RECT 1180.730 2806.090 1181.910 2807.270 ;
        RECT 1179.130 2804.490 1180.310 2805.670 ;
        RECT 1180.730 2804.490 1181.910 2805.670 ;
        RECT 1179.130 2626.090 1180.310 2627.270 ;
        RECT 1180.730 2626.090 1181.910 2627.270 ;
        RECT 1179.130 2624.490 1180.310 2625.670 ;
        RECT 1180.730 2624.490 1181.910 2625.670 ;
        RECT 1179.130 2446.090 1180.310 2447.270 ;
        RECT 1180.730 2446.090 1181.910 2447.270 ;
        RECT 1179.130 2444.490 1180.310 2445.670 ;
        RECT 1180.730 2444.490 1181.910 2445.670 ;
        RECT 1179.130 2266.090 1180.310 2267.270 ;
        RECT 1180.730 2266.090 1181.910 2267.270 ;
        RECT 1179.130 2264.490 1180.310 2265.670 ;
        RECT 1180.730 2264.490 1181.910 2265.670 ;
        RECT 1179.130 2086.090 1180.310 2087.270 ;
        RECT 1180.730 2086.090 1181.910 2087.270 ;
        RECT 1179.130 2084.490 1180.310 2085.670 ;
        RECT 1180.730 2084.490 1181.910 2085.670 ;
        RECT 1179.130 1906.090 1180.310 1907.270 ;
        RECT 1180.730 1906.090 1181.910 1907.270 ;
        RECT 1179.130 1904.490 1180.310 1905.670 ;
        RECT 1180.730 1904.490 1181.910 1905.670 ;
        RECT 1179.130 1726.090 1180.310 1727.270 ;
        RECT 1180.730 1726.090 1181.910 1727.270 ;
        RECT 1179.130 1724.490 1180.310 1725.670 ;
        RECT 1180.730 1724.490 1181.910 1725.670 ;
        RECT 1179.130 1546.090 1180.310 1547.270 ;
        RECT 1180.730 1546.090 1181.910 1547.270 ;
        RECT 1179.130 1544.490 1180.310 1545.670 ;
        RECT 1180.730 1544.490 1181.910 1545.670 ;
        RECT 1179.130 1366.090 1180.310 1367.270 ;
        RECT 1180.730 1366.090 1181.910 1367.270 ;
        RECT 1179.130 1364.490 1180.310 1365.670 ;
        RECT 1180.730 1364.490 1181.910 1365.670 ;
        RECT 1179.130 1186.090 1180.310 1187.270 ;
        RECT 1180.730 1186.090 1181.910 1187.270 ;
        RECT 1179.130 1184.490 1180.310 1185.670 ;
        RECT 1180.730 1184.490 1181.910 1185.670 ;
        RECT 99.130 1006.090 100.310 1007.270 ;
        RECT 100.730 1006.090 101.910 1007.270 ;
        RECT 99.130 1004.490 100.310 1005.670 ;
        RECT 100.730 1004.490 101.910 1005.670 ;
        RECT 1179.130 1006.090 1180.310 1007.270 ;
        RECT 1180.730 1006.090 1181.910 1007.270 ;
        RECT 1179.130 1004.490 1180.310 1005.670 ;
        RECT 1180.730 1004.490 1181.910 1005.670 ;
        RECT 99.130 826.090 100.310 827.270 ;
        RECT 100.730 826.090 101.910 827.270 ;
        RECT 99.130 824.490 100.310 825.670 ;
        RECT 100.730 824.490 101.910 825.670 ;
        RECT 99.130 646.090 100.310 647.270 ;
        RECT 100.730 646.090 101.910 647.270 ;
        RECT 99.130 644.490 100.310 645.670 ;
        RECT 100.730 644.490 101.910 645.670 ;
        RECT 99.130 466.090 100.310 467.270 ;
        RECT 100.730 466.090 101.910 467.270 ;
        RECT 99.130 464.490 100.310 465.670 ;
        RECT 100.730 464.490 101.910 465.670 ;
        RECT 298.050 826.090 299.230 827.270 ;
        RECT 298.050 824.490 299.230 825.670 ;
        RECT 298.050 646.090 299.230 647.270 ;
        RECT 298.050 644.490 299.230 645.670 ;
        RECT 298.050 466.090 299.230 467.270 ;
        RECT 298.050 464.490 299.230 465.670 ;
        RECT 451.650 826.090 452.830 827.270 ;
        RECT 451.650 824.490 452.830 825.670 ;
        RECT 451.650 646.090 452.830 647.270 ;
        RECT 451.650 644.490 452.830 645.670 ;
        RECT 451.650 466.090 452.830 467.270 ;
        RECT 451.650 464.490 452.830 465.670 ;
        RECT 605.250 826.090 606.430 827.270 ;
        RECT 605.250 824.490 606.430 825.670 ;
        RECT 605.250 646.090 606.430 647.270 ;
        RECT 605.250 644.490 606.430 645.670 ;
        RECT 605.250 466.090 606.430 467.270 ;
        RECT 605.250 464.490 606.430 465.670 ;
        RECT 758.850 826.090 760.030 827.270 ;
        RECT 758.850 824.490 760.030 825.670 ;
        RECT 758.850 646.090 760.030 647.270 ;
        RECT 758.850 644.490 760.030 645.670 ;
        RECT 758.850 466.090 760.030 467.270 ;
        RECT 758.850 464.490 760.030 465.670 ;
        RECT 912.450 826.090 913.630 827.270 ;
        RECT 912.450 824.490 913.630 825.670 ;
        RECT 912.450 646.090 913.630 647.270 ;
        RECT 912.450 644.490 913.630 645.670 ;
        RECT 912.450 466.090 913.630 467.270 ;
        RECT 912.450 464.490 913.630 465.670 ;
        RECT 1066.050 826.090 1067.230 827.270 ;
        RECT 1066.050 824.490 1067.230 825.670 ;
        RECT 1066.050 646.090 1067.230 647.270 ;
        RECT 1066.050 644.490 1067.230 645.670 ;
        RECT 1066.050 466.090 1067.230 467.270 ;
        RECT 1066.050 464.490 1067.230 465.670 ;
        RECT 1179.130 826.090 1180.310 827.270 ;
        RECT 1180.730 826.090 1181.910 827.270 ;
        RECT 1179.130 824.490 1180.310 825.670 ;
        RECT 1180.730 824.490 1181.910 825.670 ;
        RECT 1179.130 646.090 1180.310 647.270 ;
        RECT 1180.730 646.090 1181.910 647.270 ;
        RECT 1179.130 644.490 1180.310 645.670 ;
        RECT 1180.730 644.490 1181.910 645.670 ;
        RECT 1179.130 466.090 1180.310 467.270 ;
        RECT 1180.730 466.090 1181.910 467.270 ;
        RECT 1179.130 464.490 1180.310 465.670 ;
        RECT 1180.730 464.490 1181.910 465.670 ;
        RECT 99.130 286.090 100.310 287.270 ;
        RECT 100.730 286.090 101.910 287.270 ;
        RECT 99.130 284.490 100.310 285.670 ;
        RECT 100.730 284.490 101.910 285.670 ;
        RECT 99.130 106.090 100.310 107.270 ;
        RECT 100.730 106.090 101.910 107.270 ;
        RECT 99.130 104.490 100.310 105.670 ;
        RECT 100.730 104.490 101.910 105.670 ;
        RECT 99.130 -7.710 100.310 -6.530 ;
        RECT 100.730 -7.710 101.910 -6.530 ;
        RECT 99.130 -9.310 100.310 -8.130 ;
        RECT 100.730 -9.310 101.910 -8.130 ;
        RECT 279.130 286.090 280.310 287.270 ;
        RECT 280.730 286.090 281.910 287.270 ;
        RECT 279.130 284.490 280.310 285.670 ;
        RECT 280.730 284.490 281.910 285.670 ;
        RECT 279.130 106.090 280.310 107.270 ;
        RECT 280.730 106.090 281.910 107.270 ;
        RECT 279.130 104.490 280.310 105.670 ;
        RECT 280.730 104.490 281.910 105.670 ;
        RECT 279.130 -7.710 280.310 -6.530 ;
        RECT 280.730 -7.710 281.910 -6.530 ;
        RECT 279.130 -9.310 280.310 -8.130 ;
        RECT 280.730 -9.310 281.910 -8.130 ;
        RECT 459.130 286.090 460.310 287.270 ;
        RECT 460.730 286.090 461.910 287.270 ;
        RECT 459.130 284.490 460.310 285.670 ;
        RECT 460.730 284.490 461.910 285.670 ;
        RECT 459.130 106.090 460.310 107.270 ;
        RECT 460.730 106.090 461.910 107.270 ;
        RECT 459.130 104.490 460.310 105.670 ;
        RECT 460.730 104.490 461.910 105.670 ;
        RECT 459.130 -7.710 460.310 -6.530 ;
        RECT 460.730 -7.710 461.910 -6.530 ;
        RECT 459.130 -9.310 460.310 -8.130 ;
        RECT 460.730 -9.310 461.910 -8.130 ;
        RECT 639.130 286.090 640.310 287.270 ;
        RECT 640.730 286.090 641.910 287.270 ;
        RECT 639.130 284.490 640.310 285.670 ;
        RECT 640.730 284.490 641.910 285.670 ;
        RECT 639.130 106.090 640.310 107.270 ;
        RECT 640.730 106.090 641.910 107.270 ;
        RECT 639.130 104.490 640.310 105.670 ;
        RECT 640.730 104.490 641.910 105.670 ;
        RECT 639.130 -7.710 640.310 -6.530 ;
        RECT 640.730 -7.710 641.910 -6.530 ;
        RECT 639.130 -9.310 640.310 -8.130 ;
        RECT 640.730 -9.310 641.910 -8.130 ;
        RECT 819.130 286.090 820.310 287.270 ;
        RECT 820.730 286.090 821.910 287.270 ;
        RECT 819.130 284.490 820.310 285.670 ;
        RECT 820.730 284.490 821.910 285.670 ;
        RECT 819.130 106.090 820.310 107.270 ;
        RECT 820.730 106.090 821.910 107.270 ;
        RECT 819.130 104.490 820.310 105.670 ;
        RECT 820.730 104.490 821.910 105.670 ;
        RECT 819.130 -7.710 820.310 -6.530 ;
        RECT 820.730 -7.710 821.910 -6.530 ;
        RECT 819.130 -9.310 820.310 -8.130 ;
        RECT 820.730 -9.310 821.910 -8.130 ;
        RECT 999.130 286.090 1000.310 287.270 ;
        RECT 1000.730 286.090 1001.910 287.270 ;
        RECT 999.130 284.490 1000.310 285.670 ;
        RECT 1000.730 284.490 1001.910 285.670 ;
        RECT 999.130 106.090 1000.310 107.270 ;
        RECT 1000.730 106.090 1001.910 107.270 ;
        RECT 999.130 104.490 1000.310 105.670 ;
        RECT 1000.730 104.490 1001.910 105.670 ;
        RECT 999.130 -7.710 1000.310 -6.530 ;
        RECT 1000.730 -7.710 1001.910 -6.530 ;
        RECT 999.130 -9.310 1000.310 -8.130 ;
        RECT 1000.730 -9.310 1001.910 -8.130 ;
        RECT 1179.130 286.090 1180.310 287.270 ;
        RECT 1180.730 286.090 1181.910 287.270 ;
        RECT 1179.130 284.490 1180.310 285.670 ;
        RECT 1180.730 284.490 1181.910 285.670 ;
        RECT 1179.130 106.090 1180.310 107.270 ;
        RECT 1180.730 106.090 1181.910 107.270 ;
        RECT 1179.130 104.490 1180.310 105.670 ;
        RECT 1180.730 104.490 1181.910 105.670 ;
        RECT 1179.130 -7.710 1180.310 -6.530 ;
        RECT 1180.730 -7.710 1181.910 -6.530 ;
        RECT 1179.130 -9.310 1180.310 -8.130 ;
        RECT 1180.730 -9.310 1181.910 -8.130 ;
        RECT 1359.130 3527.810 1360.310 3528.990 ;
        RECT 1360.730 3527.810 1361.910 3528.990 ;
        RECT 1359.130 3526.210 1360.310 3527.390 ;
        RECT 1360.730 3526.210 1361.910 3527.390 ;
        RECT 1359.130 3346.090 1360.310 3347.270 ;
        RECT 1360.730 3346.090 1361.910 3347.270 ;
        RECT 1359.130 3344.490 1360.310 3345.670 ;
        RECT 1360.730 3344.490 1361.910 3345.670 ;
        RECT 1359.130 3166.090 1360.310 3167.270 ;
        RECT 1360.730 3166.090 1361.910 3167.270 ;
        RECT 1359.130 3164.490 1360.310 3165.670 ;
        RECT 1360.730 3164.490 1361.910 3165.670 ;
        RECT 1359.130 2986.090 1360.310 2987.270 ;
        RECT 1360.730 2986.090 1361.910 2987.270 ;
        RECT 1359.130 2984.490 1360.310 2985.670 ;
        RECT 1360.730 2984.490 1361.910 2985.670 ;
        RECT 1359.130 2806.090 1360.310 2807.270 ;
        RECT 1360.730 2806.090 1361.910 2807.270 ;
        RECT 1359.130 2804.490 1360.310 2805.670 ;
        RECT 1360.730 2804.490 1361.910 2805.670 ;
        RECT 1359.130 2626.090 1360.310 2627.270 ;
        RECT 1360.730 2626.090 1361.910 2627.270 ;
        RECT 1359.130 2624.490 1360.310 2625.670 ;
        RECT 1360.730 2624.490 1361.910 2625.670 ;
        RECT 1359.130 2446.090 1360.310 2447.270 ;
        RECT 1360.730 2446.090 1361.910 2447.270 ;
        RECT 1359.130 2444.490 1360.310 2445.670 ;
        RECT 1360.730 2444.490 1361.910 2445.670 ;
        RECT 1359.130 2266.090 1360.310 2267.270 ;
        RECT 1360.730 2266.090 1361.910 2267.270 ;
        RECT 1359.130 2264.490 1360.310 2265.670 ;
        RECT 1360.730 2264.490 1361.910 2265.670 ;
        RECT 1359.130 2086.090 1360.310 2087.270 ;
        RECT 1360.730 2086.090 1361.910 2087.270 ;
        RECT 1359.130 2084.490 1360.310 2085.670 ;
        RECT 1360.730 2084.490 1361.910 2085.670 ;
        RECT 1359.130 1906.090 1360.310 1907.270 ;
        RECT 1360.730 1906.090 1361.910 1907.270 ;
        RECT 1359.130 1904.490 1360.310 1905.670 ;
        RECT 1360.730 1904.490 1361.910 1905.670 ;
        RECT 1359.130 1726.090 1360.310 1727.270 ;
        RECT 1360.730 1726.090 1361.910 1727.270 ;
        RECT 1359.130 1724.490 1360.310 1725.670 ;
        RECT 1360.730 1724.490 1361.910 1725.670 ;
        RECT 1359.130 1546.090 1360.310 1547.270 ;
        RECT 1360.730 1546.090 1361.910 1547.270 ;
        RECT 1359.130 1544.490 1360.310 1545.670 ;
        RECT 1360.730 1544.490 1361.910 1545.670 ;
        RECT 1359.130 1366.090 1360.310 1367.270 ;
        RECT 1360.730 1366.090 1361.910 1367.270 ;
        RECT 1359.130 1364.490 1360.310 1365.670 ;
        RECT 1360.730 1364.490 1361.910 1365.670 ;
        RECT 1359.130 1186.090 1360.310 1187.270 ;
        RECT 1360.730 1186.090 1361.910 1187.270 ;
        RECT 1359.130 1184.490 1360.310 1185.670 ;
        RECT 1360.730 1184.490 1361.910 1185.670 ;
        RECT 1359.130 1006.090 1360.310 1007.270 ;
        RECT 1360.730 1006.090 1361.910 1007.270 ;
        RECT 1359.130 1004.490 1360.310 1005.670 ;
        RECT 1360.730 1004.490 1361.910 1005.670 ;
        RECT 1359.130 826.090 1360.310 827.270 ;
        RECT 1360.730 826.090 1361.910 827.270 ;
        RECT 1359.130 824.490 1360.310 825.670 ;
        RECT 1360.730 824.490 1361.910 825.670 ;
        RECT 1359.130 646.090 1360.310 647.270 ;
        RECT 1360.730 646.090 1361.910 647.270 ;
        RECT 1359.130 644.490 1360.310 645.670 ;
        RECT 1360.730 644.490 1361.910 645.670 ;
        RECT 1359.130 466.090 1360.310 467.270 ;
        RECT 1360.730 466.090 1361.910 467.270 ;
        RECT 1359.130 464.490 1360.310 465.670 ;
        RECT 1360.730 464.490 1361.910 465.670 ;
        RECT 1359.130 286.090 1360.310 287.270 ;
        RECT 1360.730 286.090 1361.910 287.270 ;
        RECT 1359.130 284.490 1360.310 285.670 ;
        RECT 1360.730 284.490 1361.910 285.670 ;
        RECT 1359.130 106.090 1360.310 107.270 ;
        RECT 1360.730 106.090 1361.910 107.270 ;
        RECT 1359.130 104.490 1360.310 105.670 ;
        RECT 1360.730 104.490 1361.910 105.670 ;
        RECT 1359.130 -7.710 1360.310 -6.530 ;
        RECT 1360.730 -7.710 1361.910 -6.530 ;
        RECT 1359.130 -9.310 1360.310 -8.130 ;
        RECT 1360.730 -9.310 1361.910 -8.130 ;
        RECT 1539.130 3527.810 1540.310 3528.990 ;
        RECT 1540.730 3527.810 1541.910 3528.990 ;
        RECT 1539.130 3526.210 1540.310 3527.390 ;
        RECT 1540.730 3526.210 1541.910 3527.390 ;
        RECT 1539.130 3346.090 1540.310 3347.270 ;
        RECT 1540.730 3346.090 1541.910 3347.270 ;
        RECT 1539.130 3344.490 1540.310 3345.670 ;
        RECT 1540.730 3344.490 1541.910 3345.670 ;
        RECT 1539.130 3166.090 1540.310 3167.270 ;
        RECT 1540.730 3166.090 1541.910 3167.270 ;
        RECT 1539.130 3164.490 1540.310 3165.670 ;
        RECT 1540.730 3164.490 1541.910 3165.670 ;
        RECT 1539.130 2986.090 1540.310 2987.270 ;
        RECT 1540.730 2986.090 1541.910 2987.270 ;
        RECT 1539.130 2984.490 1540.310 2985.670 ;
        RECT 1540.730 2984.490 1541.910 2985.670 ;
        RECT 1539.130 2806.090 1540.310 2807.270 ;
        RECT 1540.730 2806.090 1541.910 2807.270 ;
        RECT 1539.130 2804.490 1540.310 2805.670 ;
        RECT 1540.730 2804.490 1541.910 2805.670 ;
        RECT 1539.130 2626.090 1540.310 2627.270 ;
        RECT 1540.730 2626.090 1541.910 2627.270 ;
        RECT 1539.130 2624.490 1540.310 2625.670 ;
        RECT 1540.730 2624.490 1541.910 2625.670 ;
        RECT 1539.130 2446.090 1540.310 2447.270 ;
        RECT 1540.730 2446.090 1541.910 2447.270 ;
        RECT 1539.130 2444.490 1540.310 2445.670 ;
        RECT 1540.730 2444.490 1541.910 2445.670 ;
        RECT 1539.130 2266.090 1540.310 2267.270 ;
        RECT 1540.730 2266.090 1541.910 2267.270 ;
        RECT 1539.130 2264.490 1540.310 2265.670 ;
        RECT 1540.730 2264.490 1541.910 2265.670 ;
        RECT 1539.130 2086.090 1540.310 2087.270 ;
        RECT 1540.730 2086.090 1541.910 2087.270 ;
        RECT 1539.130 2084.490 1540.310 2085.670 ;
        RECT 1540.730 2084.490 1541.910 2085.670 ;
        RECT 1539.130 1906.090 1540.310 1907.270 ;
        RECT 1540.730 1906.090 1541.910 1907.270 ;
        RECT 1539.130 1904.490 1540.310 1905.670 ;
        RECT 1540.730 1904.490 1541.910 1905.670 ;
        RECT 1539.130 1726.090 1540.310 1727.270 ;
        RECT 1540.730 1726.090 1541.910 1727.270 ;
        RECT 1539.130 1724.490 1540.310 1725.670 ;
        RECT 1540.730 1724.490 1541.910 1725.670 ;
        RECT 1539.130 1546.090 1540.310 1547.270 ;
        RECT 1540.730 1546.090 1541.910 1547.270 ;
        RECT 1539.130 1544.490 1540.310 1545.670 ;
        RECT 1540.730 1544.490 1541.910 1545.670 ;
        RECT 1539.130 1366.090 1540.310 1367.270 ;
        RECT 1540.730 1366.090 1541.910 1367.270 ;
        RECT 1539.130 1364.490 1540.310 1365.670 ;
        RECT 1540.730 1364.490 1541.910 1365.670 ;
        RECT 1539.130 1186.090 1540.310 1187.270 ;
        RECT 1540.730 1186.090 1541.910 1187.270 ;
        RECT 1539.130 1184.490 1540.310 1185.670 ;
        RECT 1540.730 1184.490 1541.910 1185.670 ;
        RECT 1539.130 1006.090 1540.310 1007.270 ;
        RECT 1540.730 1006.090 1541.910 1007.270 ;
        RECT 1539.130 1004.490 1540.310 1005.670 ;
        RECT 1540.730 1004.490 1541.910 1005.670 ;
        RECT 1539.130 826.090 1540.310 827.270 ;
        RECT 1540.730 826.090 1541.910 827.270 ;
        RECT 1539.130 824.490 1540.310 825.670 ;
        RECT 1540.730 824.490 1541.910 825.670 ;
        RECT 1539.130 646.090 1540.310 647.270 ;
        RECT 1540.730 646.090 1541.910 647.270 ;
        RECT 1539.130 644.490 1540.310 645.670 ;
        RECT 1540.730 644.490 1541.910 645.670 ;
        RECT 1539.130 466.090 1540.310 467.270 ;
        RECT 1540.730 466.090 1541.910 467.270 ;
        RECT 1539.130 464.490 1540.310 465.670 ;
        RECT 1540.730 464.490 1541.910 465.670 ;
        RECT 1539.130 286.090 1540.310 287.270 ;
        RECT 1540.730 286.090 1541.910 287.270 ;
        RECT 1539.130 284.490 1540.310 285.670 ;
        RECT 1540.730 284.490 1541.910 285.670 ;
        RECT 1539.130 106.090 1540.310 107.270 ;
        RECT 1540.730 106.090 1541.910 107.270 ;
        RECT 1539.130 104.490 1540.310 105.670 ;
        RECT 1540.730 104.490 1541.910 105.670 ;
        RECT 1539.130 -7.710 1540.310 -6.530 ;
        RECT 1540.730 -7.710 1541.910 -6.530 ;
        RECT 1539.130 -9.310 1540.310 -8.130 ;
        RECT 1540.730 -9.310 1541.910 -8.130 ;
        RECT 1719.130 3527.810 1720.310 3528.990 ;
        RECT 1720.730 3527.810 1721.910 3528.990 ;
        RECT 1719.130 3526.210 1720.310 3527.390 ;
        RECT 1720.730 3526.210 1721.910 3527.390 ;
        RECT 1719.130 3346.090 1720.310 3347.270 ;
        RECT 1720.730 3346.090 1721.910 3347.270 ;
        RECT 1719.130 3344.490 1720.310 3345.670 ;
        RECT 1720.730 3344.490 1721.910 3345.670 ;
        RECT 1719.130 3166.090 1720.310 3167.270 ;
        RECT 1720.730 3166.090 1721.910 3167.270 ;
        RECT 1719.130 3164.490 1720.310 3165.670 ;
        RECT 1720.730 3164.490 1721.910 3165.670 ;
        RECT 1719.130 2986.090 1720.310 2987.270 ;
        RECT 1720.730 2986.090 1721.910 2987.270 ;
        RECT 1719.130 2984.490 1720.310 2985.670 ;
        RECT 1720.730 2984.490 1721.910 2985.670 ;
        RECT 1719.130 2806.090 1720.310 2807.270 ;
        RECT 1720.730 2806.090 1721.910 2807.270 ;
        RECT 1719.130 2804.490 1720.310 2805.670 ;
        RECT 1720.730 2804.490 1721.910 2805.670 ;
        RECT 1719.130 2626.090 1720.310 2627.270 ;
        RECT 1720.730 2626.090 1721.910 2627.270 ;
        RECT 1719.130 2624.490 1720.310 2625.670 ;
        RECT 1720.730 2624.490 1721.910 2625.670 ;
        RECT 1719.130 2446.090 1720.310 2447.270 ;
        RECT 1720.730 2446.090 1721.910 2447.270 ;
        RECT 1719.130 2444.490 1720.310 2445.670 ;
        RECT 1720.730 2444.490 1721.910 2445.670 ;
        RECT 1719.130 2266.090 1720.310 2267.270 ;
        RECT 1720.730 2266.090 1721.910 2267.270 ;
        RECT 1719.130 2264.490 1720.310 2265.670 ;
        RECT 1720.730 2264.490 1721.910 2265.670 ;
        RECT 1719.130 2086.090 1720.310 2087.270 ;
        RECT 1720.730 2086.090 1721.910 2087.270 ;
        RECT 1719.130 2084.490 1720.310 2085.670 ;
        RECT 1720.730 2084.490 1721.910 2085.670 ;
        RECT 1719.130 1906.090 1720.310 1907.270 ;
        RECT 1720.730 1906.090 1721.910 1907.270 ;
        RECT 1719.130 1904.490 1720.310 1905.670 ;
        RECT 1720.730 1904.490 1721.910 1905.670 ;
        RECT 1719.130 1726.090 1720.310 1727.270 ;
        RECT 1720.730 1726.090 1721.910 1727.270 ;
        RECT 1719.130 1724.490 1720.310 1725.670 ;
        RECT 1720.730 1724.490 1721.910 1725.670 ;
        RECT 1719.130 1546.090 1720.310 1547.270 ;
        RECT 1720.730 1546.090 1721.910 1547.270 ;
        RECT 1719.130 1544.490 1720.310 1545.670 ;
        RECT 1720.730 1544.490 1721.910 1545.670 ;
        RECT 1719.130 1366.090 1720.310 1367.270 ;
        RECT 1720.730 1366.090 1721.910 1367.270 ;
        RECT 1719.130 1364.490 1720.310 1365.670 ;
        RECT 1720.730 1364.490 1721.910 1365.670 ;
        RECT 1719.130 1186.090 1720.310 1187.270 ;
        RECT 1720.730 1186.090 1721.910 1187.270 ;
        RECT 1719.130 1184.490 1720.310 1185.670 ;
        RECT 1720.730 1184.490 1721.910 1185.670 ;
        RECT 1719.130 1006.090 1720.310 1007.270 ;
        RECT 1720.730 1006.090 1721.910 1007.270 ;
        RECT 1719.130 1004.490 1720.310 1005.670 ;
        RECT 1720.730 1004.490 1721.910 1005.670 ;
        RECT 1719.130 826.090 1720.310 827.270 ;
        RECT 1720.730 826.090 1721.910 827.270 ;
        RECT 1719.130 824.490 1720.310 825.670 ;
        RECT 1720.730 824.490 1721.910 825.670 ;
        RECT 1719.130 646.090 1720.310 647.270 ;
        RECT 1720.730 646.090 1721.910 647.270 ;
        RECT 1719.130 644.490 1720.310 645.670 ;
        RECT 1720.730 644.490 1721.910 645.670 ;
        RECT 1719.130 466.090 1720.310 467.270 ;
        RECT 1720.730 466.090 1721.910 467.270 ;
        RECT 1719.130 464.490 1720.310 465.670 ;
        RECT 1720.730 464.490 1721.910 465.670 ;
        RECT 1719.130 286.090 1720.310 287.270 ;
        RECT 1720.730 286.090 1721.910 287.270 ;
        RECT 1719.130 284.490 1720.310 285.670 ;
        RECT 1720.730 284.490 1721.910 285.670 ;
        RECT 1719.130 106.090 1720.310 107.270 ;
        RECT 1720.730 106.090 1721.910 107.270 ;
        RECT 1719.130 104.490 1720.310 105.670 ;
        RECT 1720.730 104.490 1721.910 105.670 ;
        RECT 1719.130 -7.710 1720.310 -6.530 ;
        RECT 1720.730 -7.710 1721.910 -6.530 ;
        RECT 1719.130 -9.310 1720.310 -8.130 ;
        RECT 1720.730 -9.310 1721.910 -8.130 ;
        RECT 1899.130 3527.810 1900.310 3528.990 ;
        RECT 1900.730 3527.810 1901.910 3528.990 ;
        RECT 1899.130 3526.210 1900.310 3527.390 ;
        RECT 1900.730 3526.210 1901.910 3527.390 ;
        RECT 1899.130 3346.090 1900.310 3347.270 ;
        RECT 1900.730 3346.090 1901.910 3347.270 ;
        RECT 1899.130 3344.490 1900.310 3345.670 ;
        RECT 1900.730 3344.490 1901.910 3345.670 ;
        RECT 1899.130 3166.090 1900.310 3167.270 ;
        RECT 1900.730 3166.090 1901.910 3167.270 ;
        RECT 1899.130 3164.490 1900.310 3165.670 ;
        RECT 1900.730 3164.490 1901.910 3165.670 ;
        RECT 1899.130 2986.090 1900.310 2987.270 ;
        RECT 1900.730 2986.090 1901.910 2987.270 ;
        RECT 1899.130 2984.490 1900.310 2985.670 ;
        RECT 1900.730 2984.490 1901.910 2985.670 ;
        RECT 1899.130 2806.090 1900.310 2807.270 ;
        RECT 1900.730 2806.090 1901.910 2807.270 ;
        RECT 1899.130 2804.490 1900.310 2805.670 ;
        RECT 1900.730 2804.490 1901.910 2805.670 ;
        RECT 1899.130 2626.090 1900.310 2627.270 ;
        RECT 1900.730 2626.090 1901.910 2627.270 ;
        RECT 1899.130 2624.490 1900.310 2625.670 ;
        RECT 1900.730 2624.490 1901.910 2625.670 ;
        RECT 1899.130 2446.090 1900.310 2447.270 ;
        RECT 1900.730 2446.090 1901.910 2447.270 ;
        RECT 1899.130 2444.490 1900.310 2445.670 ;
        RECT 1900.730 2444.490 1901.910 2445.670 ;
        RECT 1899.130 2266.090 1900.310 2267.270 ;
        RECT 1900.730 2266.090 1901.910 2267.270 ;
        RECT 1899.130 2264.490 1900.310 2265.670 ;
        RECT 1900.730 2264.490 1901.910 2265.670 ;
        RECT 1899.130 2086.090 1900.310 2087.270 ;
        RECT 1900.730 2086.090 1901.910 2087.270 ;
        RECT 1899.130 2084.490 1900.310 2085.670 ;
        RECT 1900.730 2084.490 1901.910 2085.670 ;
        RECT 1899.130 1906.090 1900.310 1907.270 ;
        RECT 1900.730 1906.090 1901.910 1907.270 ;
        RECT 1899.130 1904.490 1900.310 1905.670 ;
        RECT 1900.730 1904.490 1901.910 1905.670 ;
        RECT 1899.130 1726.090 1900.310 1727.270 ;
        RECT 1900.730 1726.090 1901.910 1727.270 ;
        RECT 1899.130 1724.490 1900.310 1725.670 ;
        RECT 1900.730 1724.490 1901.910 1725.670 ;
        RECT 1899.130 1546.090 1900.310 1547.270 ;
        RECT 1900.730 1546.090 1901.910 1547.270 ;
        RECT 1899.130 1544.490 1900.310 1545.670 ;
        RECT 1900.730 1544.490 1901.910 1545.670 ;
        RECT 1899.130 1366.090 1900.310 1367.270 ;
        RECT 1900.730 1366.090 1901.910 1367.270 ;
        RECT 1899.130 1364.490 1900.310 1365.670 ;
        RECT 1900.730 1364.490 1901.910 1365.670 ;
        RECT 1899.130 1186.090 1900.310 1187.270 ;
        RECT 1900.730 1186.090 1901.910 1187.270 ;
        RECT 1899.130 1184.490 1900.310 1185.670 ;
        RECT 1900.730 1184.490 1901.910 1185.670 ;
        RECT 1899.130 1006.090 1900.310 1007.270 ;
        RECT 1900.730 1006.090 1901.910 1007.270 ;
        RECT 1899.130 1004.490 1900.310 1005.670 ;
        RECT 1900.730 1004.490 1901.910 1005.670 ;
        RECT 1899.130 826.090 1900.310 827.270 ;
        RECT 1900.730 826.090 1901.910 827.270 ;
        RECT 1899.130 824.490 1900.310 825.670 ;
        RECT 1900.730 824.490 1901.910 825.670 ;
        RECT 1899.130 646.090 1900.310 647.270 ;
        RECT 1900.730 646.090 1901.910 647.270 ;
        RECT 1899.130 644.490 1900.310 645.670 ;
        RECT 1900.730 644.490 1901.910 645.670 ;
        RECT 1899.130 466.090 1900.310 467.270 ;
        RECT 1900.730 466.090 1901.910 467.270 ;
        RECT 1899.130 464.490 1900.310 465.670 ;
        RECT 1900.730 464.490 1901.910 465.670 ;
        RECT 1899.130 286.090 1900.310 287.270 ;
        RECT 1900.730 286.090 1901.910 287.270 ;
        RECT 1899.130 284.490 1900.310 285.670 ;
        RECT 1900.730 284.490 1901.910 285.670 ;
        RECT 1899.130 106.090 1900.310 107.270 ;
        RECT 1900.730 106.090 1901.910 107.270 ;
        RECT 1899.130 104.490 1900.310 105.670 ;
        RECT 1900.730 104.490 1901.910 105.670 ;
        RECT 1899.130 -7.710 1900.310 -6.530 ;
        RECT 1900.730 -7.710 1901.910 -6.530 ;
        RECT 1899.130 -9.310 1900.310 -8.130 ;
        RECT 1900.730 -9.310 1901.910 -8.130 ;
        RECT 2079.130 3527.810 2080.310 3528.990 ;
        RECT 2080.730 3527.810 2081.910 3528.990 ;
        RECT 2079.130 3526.210 2080.310 3527.390 ;
        RECT 2080.730 3526.210 2081.910 3527.390 ;
        RECT 2079.130 3346.090 2080.310 3347.270 ;
        RECT 2080.730 3346.090 2081.910 3347.270 ;
        RECT 2079.130 3344.490 2080.310 3345.670 ;
        RECT 2080.730 3344.490 2081.910 3345.670 ;
        RECT 2079.130 3166.090 2080.310 3167.270 ;
        RECT 2080.730 3166.090 2081.910 3167.270 ;
        RECT 2079.130 3164.490 2080.310 3165.670 ;
        RECT 2080.730 3164.490 2081.910 3165.670 ;
        RECT 2079.130 2986.090 2080.310 2987.270 ;
        RECT 2080.730 2986.090 2081.910 2987.270 ;
        RECT 2079.130 2984.490 2080.310 2985.670 ;
        RECT 2080.730 2984.490 2081.910 2985.670 ;
        RECT 2079.130 2806.090 2080.310 2807.270 ;
        RECT 2080.730 2806.090 2081.910 2807.270 ;
        RECT 2079.130 2804.490 2080.310 2805.670 ;
        RECT 2080.730 2804.490 2081.910 2805.670 ;
        RECT 2079.130 2626.090 2080.310 2627.270 ;
        RECT 2080.730 2626.090 2081.910 2627.270 ;
        RECT 2079.130 2624.490 2080.310 2625.670 ;
        RECT 2080.730 2624.490 2081.910 2625.670 ;
        RECT 2079.130 2446.090 2080.310 2447.270 ;
        RECT 2080.730 2446.090 2081.910 2447.270 ;
        RECT 2079.130 2444.490 2080.310 2445.670 ;
        RECT 2080.730 2444.490 2081.910 2445.670 ;
        RECT 2079.130 2266.090 2080.310 2267.270 ;
        RECT 2080.730 2266.090 2081.910 2267.270 ;
        RECT 2079.130 2264.490 2080.310 2265.670 ;
        RECT 2080.730 2264.490 2081.910 2265.670 ;
        RECT 2079.130 2086.090 2080.310 2087.270 ;
        RECT 2080.730 2086.090 2081.910 2087.270 ;
        RECT 2079.130 2084.490 2080.310 2085.670 ;
        RECT 2080.730 2084.490 2081.910 2085.670 ;
        RECT 2079.130 1906.090 2080.310 1907.270 ;
        RECT 2080.730 1906.090 2081.910 1907.270 ;
        RECT 2079.130 1904.490 2080.310 1905.670 ;
        RECT 2080.730 1904.490 2081.910 1905.670 ;
        RECT 2079.130 1726.090 2080.310 1727.270 ;
        RECT 2080.730 1726.090 2081.910 1727.270 ;
        RECT 2079.130 1724.490 2080.310 1725.670 ;
        RECT 2080.730 1724.490 2081.910 1725.670 ;
        RECT 2079.130 1546.090 2080.310 1547.270 ;
        RECT 2080.730 1546.090 2081.910 1547.270 ;
        RECT 2079.130 1544.490 2080.310 1545.670 ;
        RECT 2080.730 1544.490 2081.910 1545.670 ;
        RECT 2079.130 1366.090 2080.310 1367.270 ;
        RECT 2080.730 1366.090 2081.910 1367.270 ;
        RECT 2079.130 1364.490 2080.310 1365.670 ;
        RECT 2080.730 1364.490 2081.910 1365.670 ;
        RECT 2079.130 1186.090 2080.310 1187.270 ;
        RECT 2080.730 1186.090 2081.910 1187.270 ;
        RECT 2079.130 1184.490 2080.310 1185.670 ;
        RECT 2080.730 1184.490 2081.910 1185.670 ;
        RECT 2079.130 1006.090 2080.310 1007.270 ;
        RECT 2080.730 1006.090 2081.910 1007.270 ;
        RECT 2079.130 1004.490 2080.310 1005.670 ;
        RECT 2080.730 1004.490 2081.910 1005.670 ;
        RECT 2079.130 826.090 2080.310 827.270 ;
        RECT 2080.730 826.090 2081.910 827.270 ;
        RECT 2079.130 824.490 2080.310 825.670 ;
        RECT 2080.730 824.490 2081.910 825.670 ;
        RECT 2079.130 646.090 2080.310 647.270 ;
        RECT 2080.730 646.090 2081.910 647.270 ;
        RECT 2079.130 644.490 2080.310 645.670 ;
        RECT 2080.730 644.490 2081.910 645.670 ;
        RECT 2079.130 466.090 2080.310 467.270 ;
        RECT 2080.730 466.090 2081.910 467.270 ;
        RECT 2079.130 464.490 2080.310 465.670 ;
        RECT 2080.730 464.490 2081.910 465.670 ;
        RECT 2079.130 286.090 2080.310 287.270 ;
        RECT 2080.730 286.090 2081.910 287.270 ;
        RECT 2079.130 284.490 2080.310 285.670 ;
        RECT 2080.730 284.490 2081.910 285.670 ;
        RECT 2079.130 106.090 2080.310 107.270 ;
        RECT 2080.730 106.090 2081.910 107.270 ;
        RECT 2079.130 104.490 2080.310 105.670 ;
        RECT 2080.730 104.490 2081.910 105.670 ;
        RECT 2079.130 -7.710 2080.310 -6.530 ;
        RECT 2080.730 -7.710 2081.910 -6.530 ;
        RECT 2079.130 -9.310 2080.310 -8.130 ;
        RECT 2080.730 -9.310 2081.910 -8.130 ;
        RECT 2259.130 3527.810 2260.310 3528.990 ;
        RECT 2260.730 3527.810 2261.910 3528.990 ;
        RECT 2259.130 3526.210 2260.310 3527.390 ;
        RECT 2260.730 3526.210 2261.910 3527.390 ;
        RECT 2259.130 3346.090 2260.310 3347.270 ;
        RECT 2260.730 3346.090 2261.910 3347.270 ;
        RECT 2259.130 3344.490 2260.310 3345.670 ;
        RECT 2260.730 3344.490 2261.910 3345.670 ;
        RECT 2259.130 3166.090 2260.310 3167.270 ;
        RECT 2260.730 3166.090 2261.910 3167.270 ;
        RECT 2259.130 3164.490 2260.310 3165.670 ;
        RECT 2260.730 3164.490 2261.910 3165.670 ;
        RECT 2259.130 2986.090 2260.310 2987.270 ;
        RECT 2260.730 2986.090 2261.910 2987.270 ;
        RECT 2259.130 2984.490 2260.310 2985.670 ;
        RECT 2260.730 2984.490 2261.910 2985.670 ;
        RECT 2259.130 2806.090 2260.310 2807.270 ;
        RECT 2260.730 2806.090 2261.910 2807.270 ;
        RECT 2259.130 2804.490 2260.310 2805.670 ;
        RECT 2260.730 2804.490 2261.910 2805.670 ;
        RECT 2259.130 2626.090 2260.310 2627.270 ;
        RECT 2260.730 2626.090 2261.910 2627.270 ;
        RECT 2259.130 2624.490 2260.310 2625.670 ;
        RECT 2260.730 2624.490 2261.910 2625.670 ;
        RECT 2259.130 2446.090 2260.310 2447.270 ;
        RECT 2260.730 2446.090 2261.910 2447.270 ;
        RECT 2259.130 2444.490 2260.310 2445.670 ;
        RECT 2260.730 2444.490 2261.910 2445.670 ;
        RECT 2259.130 2266.090 2260.310 2267.270 ;
        RECT 2260.730 2266.090 2261.910 2267.270 ;
        RECT 2259.130 2264.490 2260.310 2265.670 ;
        RECT 2260.730 2264.490 2261.910 2265.670 ;
        RECT 2259.130 2086.090 2260.310 2087.270 ;
        RECT 2260.730 2086.090 2261.910 2087.270 ;
        RECT 2259.130 2084.490 2260.310 2085.670 ;
        RECT 2260.730 2084.490 2261.910 2085.670 ;
        RECT 2259.130 1906.090 2260.310 1907.270 ;
        RECT 2260.730 1906.090 2261.910 1907.270 ;
        RECT 2259.130 1904.490 2260.310 1905.670 ;
        RECT 2260.730 1904.490 2261.910 1905.670 ;
        RECT 2259.130 1726.090 2260.310 1727.270 ;
        RECT 2260.730 1726.090 2261.910 1727.270 ;
        RECT 2259.130 1724.490 2260.310 1725.670 ;
        RECT 2260.730 1724.490 2261.910 1725.670 ;
        RECT 2259.130 1546.090 2260.310 1547.270 ;
        RECT 2260.730 1546.090 2261.910 1547.270 ;
        RECT 2259.130 1544.490 2260.310 1545.670 ;
        RECT 2260.730 1544.490 2261.910 1545.670 ;
        RECT 2259.130 1366.090 2260.310 1367.270 ;
        RECT 2260.730 1366.090 2261.910 1367.270 ;
        RECT 2259.130 1364.490 2260.310 1365.670 ;
        RECT 2260.730 1364.490 2261.910 1365.670 ;
        RECT 2259.130 1186.090 2260.310 1187.270 ;
        RECT 2260.730 1186.090 2261.910 1187.270 ;
        RECT 2259.130 1184.490 2260.310 1185.670 ;
        RECT 2260.730 1184.490 2261.910 1185.670 ;
        RECT 2259.130 1006.090 2260.310 1007.270 ;
        RECT 2260.730 1006.090 2261.910 1007.270 ;
        RECT 2259.130 1004.490 2260.310 1005.670 ;
        RECT 2260.730 1004.490 2261.910 1005.670 ;
        RECT 2259.130 826.090 2260.310 827.270 ;
        RECT 2260.730 826.090 2261.910 827.270 ;
        RECT 2259.130 824.490 2260.310 825.670 ;
        RECT 2260.730 824.490 2261.910 825.670 ;
        RECT 2259.130 646.090 2260.310 647.270 ;
        RECT 2260.730 646.090 2261.910 647.270 ;
        RECT 2259.130 644.490 2260.310 645.670 ;
        RECT 2260.730 644.490 2261.910 645.670 ;
        RECT 2259.130 466.090 2260.310 467.270 ;
        RECT 2260.730 466.090 2261.910 467.270 ;
        RECT 2259.130 464.490 2260.310 465.670 ;
        RECT 2260.730 464.490 2261.910 465.670 ;
        RECT 2259.130 286.090 2260.310 287.270 ;
        RECT 2260.730 286.090 2261.910 287.270 ;
        RECT 2259.130 284.490 2260.310 285.670 ;
        RECT 2260.730 284.490 2261.910 285.670 ;
        RECT 2259.130 106.090 2260.310 107.270 ;
        RECT 2260.730 106.090 2261.910 107.270 ;
        RECT 2259.130 104.490 2260.310 105.670 ;
        RECT 2260.730 104.490 2261.910 105.670 ;
        RECT 2259.130 -7.710 2260.310 -6.530 ;
        RECT 2260.730 -7.710 2261.910 -6.530 ;
        RECT 2259.130 -9.310 2260.310 -8.130 ;
        RECT 2260.730 -9.310 2261.910 -8.130 ;
        RECT 2439.130 3527.810 2440.310 3528.990 ;
        RECT 2440.730 3527.810 2441.910 3528.990 ;
        RECT 2439.130 3526.210 2440.310 3527.390 ;
        RECT 2440.730 3526.210 2441.910 3527.390 ;
        RECT 2439.130 3346.090 2440.310 3347.270 ;
        RECT 2440.730 3346.090 2441.910 3347.270 ;
        RECT 2439.130 3344.490 2440.310 3345.670 ;
        RECT 2440.730 3344.490 2441.910 3345.670 ;
        RECT 2439.130 3166.090 2440.310 3167.270 ;
        RECT 2440.730 3166.090 2441.910 3167.270 ;
        RECT 2439.130 3164.490 2440.310 3165.670 ;
        RECT 2440.730 3164.490 2441.910 3165.670 ;
        RECT 2439.130 2986.090 2440.310 2987.270 ;
        RECT 2440.730 2986.090 2441.910 2987.270 ;
        RECT 2439.130 2984.490 2440.310 2985.670 ;
        RECT 2440.730 2984.490 2441.910 2985.670 ;
        RECT 2439.130 2806.090 2440.310 2807.270 ;
        RECT 2440.730 2806.090 2441.910 2807.270 ;
        RECT 2439.130 2804.490 2440.310 2805.670 ;
        RECT 2440.730 2804.490 2441.910 2805.670 ;
        RECT 2439.130 2626.090 2440.310 2627.270 ;
        RECT 2440.730 2626.090 2441.910 2627.270 ;
        RECT 2439.130 2624.490 2440.310 2625.670 ;
        RECT 2440.730 2624.490 2441.910 2625.670 ;
        RECT 2439.130 2446.090 2440.310 2447.270 ;
        RECT 2440.730 2446.090 2441.910 2447.270 ;
        RECT 2439.130 2444.490 2440.310 2445.670 ;
        RECT 2440.730 2444.490 2441.910 2445.670 ;
        RECT 2439.130 2266.090 2440.310 2267.270 ;
        RECT 2440.730 2266.090 2441.910 2267.270 ;
        RECT 2439.130 2264.490 2440.310 2265.670 ;
        RECT 2440.730 2264.490 2441.910 2265.670 ;
        RECT 2439.130 2086.090 2440.310 2087.270 ;
        RECT 2440.730 2086.090 2441.910 2087.270 ;
        RECT 2439.130 2084.490 2440.310 2085.670 ;
        RECT 2440.730 2084.490 2441.910 2085.670 ;
        RECT 2439.130 1906.090 2440.310 1907.270 ;
        RECT 2440.730 1906.090 2441.910 1907.270 ;
        RECT 2439.130 1904.490 2440.310 1905.670 ;
        RECT 2440.730 1904.490 2441.910 1905.670 ;
        RECT 2439.130 1726.090 2440.310 1727.270 ;
        RECT 2440.730 1726.090 2441.910 1727.270 ;
        RECT 2439.130 1724.490 2440.310 1725.670 ;
        RECT 2440.730 1724.490 2441.910 1725.670 ;
        RECT 2439.130 1546.090 2440.310 1547.270 ;
        RECT 2440.730 1546.090 2441.910 1547.270 ;
        RECT 2439.130 1544.490 2440.310 1545.670 ;
        RECT 2440.730 1544.490 2441.910 1545.670 ;
        RECT 2439.130 1366.090 2440.310 1367.270 ;
        RECT 2440.730 1366.090 2441.910 1367.270 ;
        RECT 2439.130 1364.490 2440.310 1365.670 ;
        RECT 2440.730 1364.490 2441.910 1365.670 ;
        RECT 2439.130 1186.090 2440.310 1187.270 ;
        RECT 2440.730 1186.090 2441.910 1187.270 ;
        RECT 2439.130 1184.490 2440.310 1185.670 ;
        RECT 2440.730 1184.490 2441.910 1185.670 ;
        RECT 2439.130 1006.090 2440.310 1007.270 ;
        RECT 2440.730 1006.090 2441.910 1007.270 ;
        RECT 2439.130 1004.490 2440.310 1005.670 ;
        RECT 2440.730 1004.490 2441.910 1005.670 ;
        RECT 2439.130 826.090 2440.310 827.270 ;
        RECT 2440.730 826.090 2441.910 827.270 ;
        RECT 2439.130 824.490 2440.310 825.670 ;
        RECT 2440.730 824.490 2441.910 825.670 ;
        RECT 2439.130 646.090 2440.310 647.270 ;
        RECT 2440.730 646.090 2441.910 647.270 ;
        RECT 2439.130 644.490 2440.310 645.670 ;
        RECT 2440.730 644.490 2441.910 645.670 ;
        RECT 2439.130 466.090 2440.310 467.270 ;
        RECT 2440.730 466.090 2441.910 467.270 ;
        RECT 2439.130 464.490 2440.310 465.670 ;
        RECT 2440.730 464.490 2441.910 465.670 ;
        RECT 2439.130 286.090 2440.310 287.270 ;
        RECT 2440.730 286.090 2441.910 287.270 ;
        RECT 2439.130 284.490 2440.310 285.670 ;
        RECT 2440.730 284.490 2441.910 285.670 ;
        RECT 2439.130 106.090 2440.310 107.270 ;
        RECT 2440.730 106.090 2441.910 107.270 ;
        RECT 2439.130 104.490 2440.310 105.670 ;
        RECT 2440.730 104.490 2441.910 105.670 ;
        RECT 2439.130 -7.710 2440.310 -6.530 ;
        RECT 2440.730 -7.710 2441.910 -6.530 ;
        RECT 2439.130 -9.310 2440.310 -8.130 ;
        RECT 2440.730 -9.310 2441.910 -8.130 ;
        RECT 2619.130 3527.810 2620.310 3528.990 ;
        RECT 2620.730 3527.810 2621.910 3528.990 ;
        RECT 2619.130 3526.210 2620.310 3527.390 ;
        RECT 2620.730 3526.210 2621.910 3527.390 ;
        RECT 2619.130 3346.090 2620.310 3347.270 ;
        RECT 2620.730 3346.090 2621.910 3347.270 ;
        RECT 2619.130 3344.490 2620.310 3345.670 ;
        RECT 2620.730 3344.490 2621.910 3345.670 ;
        RECT 2619.130 3166.090 2620.310 3167.270 ;
        RECT 2620.730 3166.090 2621.910 3167.270 ;
        RECT 2619.130 3164.490 2620.310 3165.670 ;
        RECT 2620.730 3164.490 2621.910 3165.670 ;
        RECT 2619.130 2986.090 2620.310 2987.270 ;
        RECT 2620.730 2986.090 2621.910 2987.270 ;
        RECT 2619.130 2984.490 2620.310 2985.670 ;
        RECT 2620.730 2984.490 2621.910 2985.670 ;
        RECT 2619.130 2806.090 2620.310 2807.270 ;
        RECT 2620.730 2806.090 2621.910 2807.270 ;
        RECT 2619.130 2804.490 2620.310 2805.670 ;
        RECT 2620.730 2804.490 2621.910 2805.670 ;
        RECT 2619.130 2626.090 2620.310 2627.270 ;
        RECT 2620.730 2626.090 2621.910 2627.270 ;
        RECT 2619.130 2624.490 2620.310 2625.670 ;
        RECT 2620.730 2624.490 2621.910 2625.670 ;
        RECT 2619.130 2446.090 2620.310 2447.270 ;
        RECT 2620.730 2446.090 2621.910 2447.270 ;
        RECT 2619.130 2444.490 2620.310 2445.670 ;
        RECT 2620.730 2444.490 2621.910 2445.670 ;
        RECT 2619.130 2266.090 2620.310 2267.270 ;
        RECT 2620.730 2266.090 2621.910 2267.270 ;
        RECT 2619.130 2264.490 2620.310 2265.670 ;
        RECT 2620.730 2264.490 2621.910 2265.670 ;
        RECT 2619.130 2086.090 2620.310 2087.270 ;
        RECT 2620.730 2086.090 2621.910 2087.270 ;
        RECT 2619.130 2084.490 2620.310 2085.670 ;
        RECT 2620.730 2084.490 2621.910 2085.670 ;
        RECT 2619.130 1906.090 2620.310 1907.270 ;
        RECT 2620.730 1906.090 2621.910 1907.270 ;
        RECT 2619.130 1904.490 2620.310 1905.670 ;
        RECT 2620.730 1904.490 2621.910 1905.670 ;
        RECT 2619.130 1726.090 2620.310 1727.270 ;
        RECT 2620.730 1726.090 2621.910 1727.270 ;
        RECT 2619.130 1724.490 2620.310 1725.670 ;
        RECT 2620.730 1724.490 2621.910 1725.670 ;
        RECT 2619.130 1546.090 2620.310 1547.270 ;
        RECT 2620.730 1546.090 2621.910 1547.270 ;
        RECT 2619.130 1544.490 2620.310 1545.670 ;
        RECT 2620.730 1544.490 2621.910 1545.670 ;
        RECT 2619.130 1366.090 2620.310 1367.270 ;
        RECT 2620.730 1366.090 2621.910 1367.270 ;
        RECT 2619.130 1364.490 2620.310 1365.670 ;
        RECT 2620.730 1364.490 2621.910 1365.670 ;
        RECT 2619.130 1186.090 2620.310 1187.270 ;
        RECT 2620.730 1186.090 2621.910 1187.270 ;
        RECT 2619.130 1184.490 2620.310 1185.670 ;
        RECT 2620.730 1184.490 2621.910 1185.670 ;
        RECT 2619.130 1006.090 2620.310 1007.270 ;
        RECT 2620.730 1006.090 2621.910 1007.270 ;
        RECT 2619.130 1004.490 2620.310 1005.670 ;
        RECT 2620.730 1004.490 2621.910 1005.670 ;
        RECT 2619.130 826.090 2620.310 827.270 ;
        RECT 2620.730 826.090 2621.910 827.270 ;
        RECT 2619.130 824.490 2620.310 825.670 ;
        RECT 2620.730 824.490 2621.910 825.670 ;
        RECT 2619.130 646.090 2620.310 647.270 ;
        RECT 2620.730 646.090 2621.910 647.270 ;
        RECT 2619.130 644.490 2620.310 645.670 ;
        RECT 2620.730 644.490 2621.910 645.670 ;
        RECT 2619.130 466.090 2620.310 467.270 ;
        RECT 2620.730 466.090 2621.910 467.270 ;
        RECT 2619.130 464.490 2620.310 465.670 ;
        RECT 2620.730 464.490 2621.910 465.670 ;
        RECT 2619.130 286.090 2620.310 287.270 ;
        RECT 2620.730 286.090 2621.910 287.270 ;
        RECT 2619.130 284.490 2620.310 285.670 ;
        RECT 2620.730 284.490 2621.910 285.670 ;
        RECT 2619.130 106.090 2620.310 107.270 ;
        RECT 2620.730 106.090 2621.910 107.270 ;
        RECT 2619.130 104.490 2620.310 105.670 ;
        RECT 2620.730 104.490 2621.910 105.670 ;
        RECT 2619.130 -7.710 2620.310 -6.530 ;
        RECT 2620.730 -7.710 2621.910 -6.530 ;
        RECT 2619.130 -9.310 2620.310 -8.130 ;
        RECT 2620.730 -9.310 2621.910 -8.130 ;
        RECT 2799.130 3527.810 2800.310 3528.990 ;
        RECT 2800.730 3527.810 2801.910 3528.990 ;
        RECT 2799.130 3526.210 2800.310 3527.390 ;
        RECT 2800.730 3526.210 2801.910 3527.390 ;
        RECT 2799.130 3346.090 2800.310 3347.270 ;
        RECT 2800.730 3346.090 2801.910 3347.270 ;
        RECT 2799.130 3344.490 2800.310 3345.670 ;
        RECT 2800.730 3344.490 2801.910 3345.670 ;
        RECT 2799.130 3166.090 2800.310 3167.270 ;
        RECT 2800.730 3166.090 2801.910 3167.270 ;
        RECT 2799.130 3164.490 2800.310 3165.670 ;
        RECT 2800.730 3164.490 2801.910 3165.670 ;
        RECT 2799.130 2986.090 2800.310 2987.270 ;
        RECT 2800.730 2986.090 2801.910 2987.270 ;
        RECT 2799.130 2984.490 2800.310 2985.670 ;
        RECT 2800.730 2984.490 2801.910 2985.670 ;
        RECT 2799.130 2806.090 2800.310 2807.270 ;
        RECT 2800.730 2806.090 2801.910 2807.270 ;
        RECT 2799.130 2804.490 2800.310 2805.670 ;
        RECT 2800.730 2804.490 2801.910 2805.670 ;
        RECT 2799.130 2626.090 2800.310 2627.270 ;
        RECT 2800.730 2626.090 2801.910 2627.270 ;
        RECT 2799.130 2624.490 2800.310 2625.670 ;
        RECT 2800.730 2624.490 2801.910 2625.670 ;
        RECT 2799.130 2446.090 2800.310 2447.270 ;
        RECT 2800.730 2446.090 2801.910 2447.270 ;
        RECT 2799.130 2444.490 2800.310 2445.670 ;
        RECT 2800.730 2444.490 2801.910 2445.670 ;
        RECT 2799.130 2266.090 2800.310 2267.270 ;
        RECT 2800.730 2266.090 2801.910 2267.270 ;
        RECT 2799.130 2264.490 2800.310 2265.670 ;
        RECT 2800.730 2264.490 2801.910 2265.670 ;
        RECT 2799.130 2086.090 2800.310 2087.270 ;
        RECT 2800.730 2086.090 2801.910 2087.270 ;
        RECT 2799.130 2084.490 2800.310 2085.670 ;
        RECT 2800.730 2084.490 2801.910 2085.670 ;
        RECT 2799.130 1906.090 2800.310 1907.270 ;
        RECT 2800.730 1906.090 2801.910 1907.270 ;
        RECT 2799.130 1904.490 2800.310 1905.670 ;
        RECT 2800.730 1904.490 2801.910 1905.670 ;
        RECT 2799.130 1726.090 2800.310 1727.270 ;
        RECT 2800.730 1726.090 2801.910 1727.270 ;
        RECT 2799.130 1724.490 2800.310 1725.670 ;
        RECT 2800.730 1724.490 2801.910 1725.670 ;
        RECT 2799.130 1546.090 2800.310 1547.270 ;
        RECT 2800.730 1546.090 2801.910 1547.270 ;
        RECT 2799.130 1544.490 2800.310 1545.670 ;
        RECT 2800.730 1544.490 2801.910 1545.670 ;
        RECT 2799.130 1366.090 2800.310 1367.270 ;
        RECT 2800.730 1366.090 2801.910 1367.270 ;
        RECT 2799.130 1364.490 2800.310 1365.670 ;
        RECT 2800.730 1364.490 2801.910 1365.670 ;
        RECT 2799.130 1186.090 2800.310 1187.270 ;
        RECT 2800.730 1186.090 2801.910 1187.270 ;
        RECT 2799.130 1184.490 2800.310 1185.670 ;
        RECT 2800.730 1184.490 2801.910 1185.670 ;
        RECT 2799.130 1006.090 2800.310 1007.270 ;
        RECT 2800.730 1006.090 2801.910 1007.270 ;
        RECT 2799.130 1004.490 2800.310 1005.670 ;
        RECT 2800.730 1004.490 2801.910 1005.670 ;
        RECT 2799.130 826.090 2800.310 827.270 ;
        RECT 2800.730 826.090 2801.910 827.270 ;
        RECT 2799.130 824.490 2800.310 825.670 ;
        RECT 2800.730 824.490 2801.910 825.670 ;
        RECT 2799.130 646.090 2800.310 647.270 ;
        RECT 2800.730 646.090 2801.910 647.270 ;
        RECT 2799.130 644.490 2800.310 645.670 ;
        RECT 2800.730 644.490 2801.910 645.670 ;
        RECT 2799.130 466.090 2800.310 467.270 ;
        RECT 2800.730 466.090 2801.910 467.270 ;
        RECT 2799.130 464.490 2800.310 465.670 ;
        RECT 2800.730 464.490 2801.910 465.670 ;
        RECT 2799.130 286.090 2800.310 287.270 ;
        RECT 2800.730 286.090 2801.910 287.270 ;
        RECT 2799.130 284.490 2800.310 285.670 ;
        RECT 2800.730 284.490 2801.910 285.670 ;
        RECT 2799.130 106.090 2800.310 107.270 ;
        RECT 2800.730 106.090 2801.910 107.270 ;
        RECT 2799.130 104.490 2800.310 105.670 ;
        RECT 2800.730 104.490 2801.910 105.670 ;
        RECT 2799.130 -7.710 2800.310 -6.530 ;
        RECT 2800.730 -7.710 2801.910 -6.530 ;
        RECT 2799.130 -9.310 2800.310 -8.130 ;
        RECT 2800.730 -9.310 2801.910 -8.130 ;
        RECT 2931.510 3527.810 2932.690 3528.990 ;
        RECT 2933.110 3527.810 2934.290 3528.990 ;
        RECT 2931.510 3526.210 2932.690 3527.390 ;
        RECT 2933.110 3526.210 2934.290 3527.390 ;
        RECT 2931.510 3346.090 2932.690 3347.270 ;
        RECT 2933.110 3346.090 2934.290 3347.270 ;
        RECT 2931.510 3344.490 2932.690 3345.670 ;
        RECT 2933.110 3344.490 2934.290 3345.670 ;
        RECT 2931.510 3166.090 2932.690 3167.270 ;
        RECT 2933.110 3166.090 2934.290 3167.270 ;
        RECT 2931.510 3164.490 2932.690 3165.670 ;
        RECT 2933.110 3164.490 2934.290 3165.670 ;
        RECT 2931.510 2986.090 2932.690 2987.270 ;
        RECT 2933.110 2986.090 2934.290 2987.270 ;
        RECT 2931.510 2984.490 2932.690 2985.670 ;
        RECT 2933.110 2984.490 2934.290 2985.670 ;
        RECT 2931.510 2806.090 2932.690 2807.270 ;
        RECT 2933.110 2806.090 2934.290 2807.270 ;
        RECT 2931.510 2804.490 2932.690 2805.670 ;
        RECT 2933.110 2804.490 2934.290 2805.670 ;
        RECT 2931.510 2626.090 2932.690 2627.270 ;
        RECT 2933.110 2626.090 2934.290 2627.270 ;
        RECT 2931.510 2624.490 2932.690 2625.670 ;
        RECT 2933.110 2624.490 2934.290 2625.670 ;
        RECT 2931.510 2446.090 2932.690 2447.270 ;
        RECT 2933.110 2446.090 2934.290 2447.270 ;
        RECT 2931.510 2444.490 2932.690 2445.670 ;
        RECT 2933.110 2444.490 2934.290 2445.670 ;
        RECT 2931.510 2266.090 2932.690 2267.270 ;
        RECT 2933.110 2266.090 2934.290 2267.270 ;
        RECT 2931.510 2264.490 2932.690 2265.670 ;
        RECT 2933.110 2264.490 2934.290 2265.670 ;
        RECT 2931.510 2086.090 2932.690 2087.270 ;
        RECT 2933.110 2086.090 2934.290 2087.270 ;
        RECT 2931.510 2084.490 2932.690 2085.670 ;
        RECT 2933.110 2084.490 2934.290 2085.670 ;
        RECT 2931.510 1906.090 2932.690 1907.270 ;
        RECT 2933.110 1906.090 2934.290 1907.270 ;
        RECT 2931.510 1904.490 2932.690 1905.670 ;
        RECT 2933.110 1904.490 2934.290 1905.670 ;
        RECT 2931.510 1726.090 2932.690 1727.270 ;
        RECT 2933.110 1726.090 2934.290 1727.270 ;
        RECT 2931.510 1724.490 2932.690 1725.670 ;
        RECT 2933.110 1724.490 2934.290 1725.670 ;
        RECT 2931.510 1546.090 2932.690 1547.270 ;
        RECT 2933.110 1546.090 2934.290 1547.270 ;
        RECT 2931.510 1544.490 2932.690 1545.670 ;
        RECT 2933.110 1544.490 2934.290 1545.670 ;
        RECT 2931.510 1366.090 2932.690 1367.270 ;
        RECT 2933.110 1366.090 2934.290 1367.270 ;
        RECT 2931.510 1364.490 2932.690 1365.670 ;
        RECT 2933.110 1364.490 2934.290 1365.670 ;
        RECT 2931.510 1186.090 2932.690 1187.270 ;
        RECT 2933.110 1186.090 2934.290 1187.270 ;
        RECT 2931.510 1184.490 2932.690 1185.670 ;
        RECT 2933.110 1184.490 2934.290 1185.670 ;
        RECT 2931.510 1006.090 2932.690 1007.270 ;
        RECT 2933.110 1006.090 2934.290 1007.270 ;
        RECT 2931.510 1004.490 2932.690 1005.670 ;
        RECT 2933.110 1004.490 2934.290 1005.670 ;
        RECT 2931.510 826.090 2932.690 827.270 ;
        RECT 2933.110 826.090 2934.290 827.270 ;
        RECT 2931.510 824.490 2932.690 825.670 ;
        RECT 2933.110 824.490 2934.290 825.670 ;
        RECT 2931.510 646.090 2932.690 647.270 ;
        RECT 2933.110 646.090 2934.290 647.270 ;
        RECT 2931.510 644.490 2932.690 645.670 ;
        RECT 2933.110 644.490 2934.290 645.670 ;
        RECT 2931.510 466.090 2932.690 467.270 ;
        RECT 2933.110 466.090 2934.290 467.270 ;
        RECT 2931.510 464.490 2932.690 465.670 ;
        RECT 2933.110 464.490 2934.290 465.670 ;
        RECT 2931.510 286.090 2932.690 287.270 ;
        RECT 2933.110 286.090 2934.290 287.270 ;
        RECT 2931.510 284.490 2932.690 285.670 ;
        RECT 2933.110 284.490 2934.290 285.670 ;
        RECT 2931.510 106.090 2932.690 107.270 ;
        RECT 2933.110 106.090 2934.290 107.270 ;
        RECT 2931.510 104.490 2932.690 105.670 ;
        RECT 2933.110 104.490 2934.290 105.670 ;
        RECT 2931.510 -7.710 2932.690 -6.530 ;
        RECT 2933.110 -7.710 2934.290 -6.530 ;
        RECT 2931.510 -9.310 2932.690 -8.130 ;
        RECT 2933.110 -9.310 2934.290 -8.130 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
        RECT -14.830 824.330 2934.450 827.430 ;
        RECT -14.830 644.330 2934.450 647.430 ;
        RECT -14.830 464.330 2934.450 467.430 ;
        RECT -14.830 284.330 2934.450 287.430 ;
        RECT -14.830 104.330 2934.450 107.430 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
        RECT 297.570 1010.000 300.670 3538.750 ;
        RECT 477.570 1010.000 480.670 3538.750 ;
        RECT 657.570 1010.000 660.670 3538.750 ;
        RECT 837.570 1010.000 840.670 3538.750 ;
        RECT 1017.570 1010.000 1020.670 3538.750 ;
        RECT 297.570 -19.070 300.670 390.000 ;
        RECT 477.570 -19.070 480.670 390.000 ;
        RECT 657.570 -19.070 660.670 390.000 ;
        RECT 837.570 -19.070 840.670 390.000 ;
        RECT 1017.570 -19.070 1020.670 390.000 ;
        RECT 1197.570 -19.070 1200.670 3538.750 ;
        RECT 1377.570 -19.070 1380.670 3538.750 ;
        RECT 1557.570 -19.070 1560.670 3538.750 ;
        RECT 1737.570 -19.070 1740.670 3538.750 ;
        RECT 1917.570 -19.070 1920.670 3538.750 ;
        RECT 2097.570 -19.070 2100.670 3538.750 ;
        RECT 2277.570 -19.070 2280.670 3538.750 ;
        RECT 2457.570 -19.070 2460.670 3538.750 ;
        RECT 2637.570 -19.070 2640.670 3538.750 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER via4 ;
        RECT -24.270 3537.410 -23.090 3538.590 ;
        RECT -22.670 3537.410 -21.490 3538.590 ;
        RECT -24.270 3535.810 -23.090 3536.990 ;
        RECT -22.670 3535.810 -21.490 3536.990 ;
        RECT -24.270 3364.690 -23.090 3365.870 ;
        RECT -22.670 3364.690 -21.490 3365.870 ;
        RECT -24.270 3363.090 -23.090 3364.270 ;
        RECT -22.670 3363.090 -21.490 3364.270 ;
        RECT -24.270 3184.690 -23.090 3185.870 ;
        RECT -22.670 3184.690 -21.490 3185.870 ;
        RECT -24.270 3183.090 -23.090 3184.270 ;
        RECT -22.670 3183.090 -21.490 3184.270 ;
        RECT -24.270 3004.690 -23.090 3005.870 ;
        RECT -22.670 3004.690 -21.490 3005.870 ;
        RECT -24.270 3003.090 -23.090 3004.270 ;
        RECT -22.670 3003.090 -21.490 3004.270 ;
        RECT -24.270 2824.690 -23.090 2825.870 ;
        RECT -22.670 2824.690 -21.490 2825.870 ;
        RECT -24.270 2823.090 -23.090 2824.270 ;
        RECT -22.670 2823.090 -21.490 2824.270 ;
        RECT -24.270 2644.690 -23.090 2645.870 ;
        RECT -22.670 2644.690 -21.490 2645.870 ;
        RECT -24.270 2643.090 -23.090 2644.270 ;
        RECT -22.670 2643.090 -21.490 2644.270 ;
        RECT -24.270 2464.690 -23.090 2465.870 ;
        RECT -22.670 2464.690 -21.490 2465.870 ;
        RECT -24.270 2463.090 -23.090 2464.270 ;
        RECT -22.670 2463.090 -21.490 2464.270 ;
        RECT -24.270 2284.690 -23.090 2285.870 ;
        RECT -22.670 2284.690 -21.490 2285.870 ;
        RECT -24.270 2283.090 -23.090 2284.270 ;
        RECT -22.670 2283.090 -21.490 2284.270 ;
        RECT -24.270 2104.690 -23.090 2105.870 ;
        RECT -22.670 2104.690 -21.490 2105.870 ;
        RECT -24.270 2103.090 -23.090 2104.270 ;
        RECT -22.670 2103.090 -21.490 2104.270 ;
        RECT -24.270 1924.690 -23.090 1925.870 ;
        RECT -22.670 1924.690 -21.490 1925.870 ;
        RECT -24.270 1923.090 -23.090 1924.270 ;
        RECT -22.670 1923.090 -21.490 1924.270 ;
        RECT -24.270 1744.690 -23.090 1745.870 ;
        RECT -22.670 1744.690 -21.490 1745.870 ;
        RECT -24.270 1743.090 -23.090 1744.270 ;
        RECT -22.670 1743.090 -21.490 1744.270 ;
        RECT -24.270 1564.690 -23.090 1565.870 ;
        RECT -22.670 1564.690 -21.490 1565.870 ;
        RECT -24.270 1563.090 -23.090 1564.270 ;
        RECT -22.670 1563.090 -21.490 1564.270 ;
        RECT -24.270 1384.690 -23.090 1385.870 ;
        RECT -22.670 1384.690 -21.490 1385.870 ;
        RECT -24.270 1383.090 -23.090 1384.270 ;
        RECT -22.670 1383.090 -21.490 1384.270 ;
        RECT -24.270 1204.690 -23.090 1205.870 ;
        RECT -22.670 1204.690 -21.490 1205.870 ;
        RECT -24.270 1203.090 -23.090 1204.270 ;
        RECT -22.670 1203.090 -21.490 1204.270 ;
        RECT -24.270 1024.690 -23.090 1025.870 ;
        RECT -22.670 1024.690 -21.490 1025.870 ;
        RECT -24.270 1023.090 -23.090 1024.270 ;
        RECT -22.670 1023.090 -21.490 1024.270 ;
        RECT -24.270 844.690 -23.090 845.870 ;
        RECT -22.670 844.690 -21.490 845.870 ;
        RECT -24.270 843.090 -23.090 844.270 ;
        RECT -22.670 843.090 -21.490 844.270 ;
        RECT -24.270 664.690 -23.090 665.870 ;
        RECT -22.670 664.690 -21.490 665.870 ;
        RECT -24.270 663.090 -23.090 664.270 ;
        RECT -22.670 663.090 -21.490 664.270 ;
        RECT -24.270 484.690 -23.090 485.870 ;
        RECT -22.670 484.690 -21.490 485.870 ;
        RECT -24.270 483.090 -23.090 484.270 ;
        RECT -22.670 483.090 -21.490 484.270 ;
        RECT -24.270 304.690 -23.090 305.870 ;
        RECT -22.670 304.690 -21.490 305.870 ;
        RECT -24.270 303.090 -23.090 304.270 ;
        RECT -22.670 303.090 -21.490 304.270 ;
        RECT -24.270 124.690 -23.090 125.870 ;
        RECT -22.670 124.690 -21.490 125.870 ;
        RECT -24.270 123.090 -23.090 124.270 ;
        RECT -22.670 123.090 -21.490 124.270 ;
        RECT -24.270 -17.310 -23.090 -16.130 ;
        RECT -22.670 -17.310 -21.490 -16.130 ;
        RECT -24.270 -18.910 -23.090 -17.730 ;
        RECT -22.670 -18.910 -21.490 -17.730 ;
        RECT 117.730 3537.410 118.910 3538.590 ;
        RECT 119.330 3537.410 120.510 3538.590 ;
        RECT 117.730 3535.810 118.910 3536.990 ;
        RECT 119.330 3535.810 120.510 3536.990 ;
        RECT 117.730 3364.690 118.910 3365.870 ;
        RECT 119.330 3364.690 120.510 3365.870 ;
        RECT 117.730 3363.090 118.910 3364.270 ;
        RECT 119.330 3363.090 120.510 3364.270 ;
        RECT 117.730 3184.690 118.910 3185.870 ;
        RECT 119.330 3184.690 120.510 3185.870 ;
        RECT 117.730 3183.090 118.910 3184.270 ;
        RECT 119.330 3183.090 120.510 3184.270 ;
        RECT 117.730 3004.690 118.910 3005.870 ;
        RECT 119.330 3004.690 120.510 3005.870 ;
        RECT 117.730 3003.090 118.910 3004.270 ;
        RECT 119.330 3003.090 120.510 3004.270 ;
        RECT 117.730 2824.690 118.910 2825.870 ;
        RECT 119.330 2824.690 120.510 2825.870 ;
        RECT 117.730 2823.090 118.910 2824.270 ;
        RECT 119.330 2823.090 120.510 2824.270 ;
        RECT 117.730 2644.690 118.910 2645.870 ;
        RECT 119.330 2644.690 120.510 2645.870 ;
        RECT 117.730 2643.090 118.910 2644.270 ;
        RECT 119.330 2643.090 120.510 2644.270 ;
        RECT 117.730 2464.690 118.910 2465.870 ;
        RECT 119.330 2464.690 120.510 2465.870 ;
        RECT 117.730 2463.090 118.910 2464.270 ;
        RECT 119.330 2463.090 120.510 2464.270 ;
        RECT 117.730 2284.690 118.910 2285.870 ;
        RECT 119.330 2284.690 120.510 2285.870 ;
        RECT 117.730 2283.090 118.910 2284.270 ;
        RECT 119.330 2283.090 120.510 2284.270 ;
        RECT 117.730 2104.690 118.910 2105.870 ;
        RECT 119.330 2104.690 120.510 2105.870 ;
        RECT 117.730 2103.090 118.910 2104.270 ;
        RECT 119.330 2103.090 120.510 2104.270 ;
        RECT 117.730 1924.690 118.910 1925.870 ;
        RECT 119.330 1924.690 120.510 1925.870 ;
        RECT 117.730 1923.090 118.910 1924.270 ;
        RECT 119.330 1923.090 120.510 1924.270 ;
        RECT 117.730 1744.690 118.910 1745.870 ;
        RECT 119.330 1744.690 120.510 1745.870 ;
        RECT 117.730 1743.090 118.910 1744.270 ;
        RECT 119.330 1743.090 120.510 1744.270 ;
        RECT 117.730 1564.690 118.910 1565.870 ;
        RECT 119.330 1564.690 120.510 1565.870 ;
        RECT 117.730 1563.090 118.910 1564.270 ;
        RECT 119.330 1563.090 120.510 1564.270 ;
        RECT 117.730 1384.690 118.910 1385.870 ;
        RECT 119.330 1384.690 120.510 1385.870 ;
        RECT 117.730 1383.090 118.910 1384.270 ;
        RECT 119.330 1383.090 120.510 1384.270 ;
        RECT 117.730 1204.690 118.910 1205.870 ;
        RECT 119.330 1204.690 120.510 1205.870 ;
        RECT 117.730 1203.090 118.910 1204.270 ;
        RECT 119.330 1203.090 120.510 1204.270 ;
        RECT 117.730 1024.690 118.910 1025.870 ;
        RECT 119.330 1024.690 120.510 1025.870 ;
        RECT 117.730 1023.090 118.910 1024.270 ;
        RECT 119.330 1023.090 120.510 1024.270 ;
        RECT 297.730 3537.410 298.910 3538.590 ;
        RECT 299.330 3537.410 300.510 3538.590 ;
        RECT 297.730 3535.810 298.910 3536.990 ;
        RECT 299.330 3535.810 300.510 3536.990 ;
        RECT 297.730 3364.690 298.910 3365.870 ;
        RECT 299.330 3364.690 300.510 3365.870 ;
        RECT 297.730 3363.090 298.910 3364.270 ;
        RECT 299.330 3363.090 300.510 3364.270 ;
        RECT 297.730 3184.690 298.910 3185.870 ;
        RECT 299.330 3184.690 300.510 3185.870 ;
        RECT 297.730 3183.090 298.910 3184.270 ;
        RECT 299.330 3183.090 300.510 3184.270 ;
        RECT 297.730 3004.690 298.910 3005.870 ;
        RECT 299.330 3004.690 300.510 3005.870 ;
        RECT 297.730 3003.090 298.910 3004.270 ;
        RECT 299.330 3003.090 300.510 3004.270 ;
        RECT 297.730 2824.690 298.910 2825.870 ;
        RECT 299.330 2824.690 300.510 2825.870 ;
        RECT 297.730 2823.090 298.910 2824.270 ;
        RECT 299.330 2823.090 300.510 2824.270 ;
        RECT 297.730 2644.690 298.910 2645.870 ;
        RECT 299.330 2644.690 300.510 2645.870 ;
        RECT 297.730 2643.090 298.910 2644.270 ;
        RECT 299.330 2643.090 300.510 2644.270 ;
        RECT 297.730 2464.690 298.910 2465.870 ;
        RECT 299.330 2464.690 300.510 2465.870 ;
        RECT 297.730 2463.090 298.910 2464.270 ;
        RECT 299.330 2463.090 300.510 2464.270 ;
        RECT 297.730 2284.690 298.910 2285.870 ;
        RECT 299.330 2284.690 300.510 2285.870 ;
        RECT 297.730 2283.090 298.910 2284.270 ;
        RECT 299.330 2283.090 300.510 2284.270 ;
        RECT 297.730 2104.690 298.910 2105.870 ;
        RECT 299.330 2104.690 300.510 2105.870 ;
        RECT 297.730 2103.090 298.910 2104.270 ;
        RECT 299.330 2103.090 300.510 2104.270 ;
        RECT 297.730 1924.690 298.910 1925.870 ;
        RECT 299.330 1924.690 300.510 1925.870 ;
        RECT 297.730 1923.090 298.910 1924.270 ;
        RECT 299.330 1923.090 300.510 1924.270 ;
        RECT 297.730 1744.690 298.910 1745.870 ;
        RECT 299.330 1744.690 300.510 1745.870 ;
        RECT 297.730 1743.090 298.910 1744.270 ;
        RECT 299.330 1743.090 300.510 1744.270 ;
        RECT 297.730 1564.690 298.910 1565.870 ;
        RECT 299.330 1564.690 300.510 1565.870 ;
        RECT 297.730 1563.090 298.910 1564.270 ;
        RECT 299.330 1563.090 300.510 1564.270 ;
        RECT 297.730 1384.690 298.910 1385.870 ;
        RECT 299.330 1384.690 300.510 1385.870 ;
        RECT 297.730 1383.090 298.910 1384.270 ;
        RECT 299.330 1383.090 300.510 1384.270 ;
        RECT 297.730 1204.690 298.910 1205.870 ;
        RECT 299.330 1204.690 300.510 1205.870 ;
        RECT 297.730 1203.090 298.910 1204.270 ;
        RECT 299.330 1203.090 300.510 1204.270 ;
        RECT 297.730 1024.690 298.910 1025.870 ;
        RECT 299.330 1024.690 300.510 1025.870 ;
        RECT 297.730 1023.090 298.910 1024.270 ;
        RECT 299.330 1023.090 300.510 1024.270 ;
        RECT 477.730 3537.410 478.910 3538.590 ;
        RECT 479.330 3537.410 480.510 3538.590 ;
        RECT 477.730 3535.810 478.910 3536.990 ;
        RECT 479.330 3535.810 480.510 3536.990 ;
        RECT 477.730 3364.690 478.910 3365.870 ;
        RECT 479.330 3364.690 480.510 3365.870 ;
        RECT 477.730 3363.090 478.910 3364.270 ;
        RECT 479.330 3363.090 480.510 3364.270 ;
        RECT 477.730 3184.690 478.910 3185.870 ;
        RECT 479.330 3184.690 480.510 3185.870 ;
        RECT 477.730 3183.090 478.910 3184.270 ;
        RECT 479.330 3183.090 480.510 3184.270 ;
        RECT 477.730 3004.690 478.910 3005.870 ;
        RECT 479.330 3004.690 480.510 3005.870 ;
        RECT 477.730 3003.090 478.910 3004.270 ;
        RECT 479.330 3003.090 480.510 3004.270 ;
        RECT 477.730 2824.690 478.910 2825.870 ;
        RECT 479.330 2824.690 480.510 2825.870 ;
        RECT 477.730 2823.090 478.910 2824.270 ;
        RECT 479.330 2823.090 480.510 2824.270 ;
        RECT 477.730 2644.690 478.910 2645.870 ;
        RECT 479.330 2644.690 480.510 2645.870 ;
        RECT 477.730 2643.090 478.910 2644.270 ;
        RECT 479.330 2643.090 480.510 2644.270 ;
        RECT 477.730 2464.690 478.910 2465.870 ;
        RECT 479.330 2464.690 480.510 2465.870 ;
        RECT 477.730 2463.090 478.910 2464.270 ;
        RECT 479.330 2463.090 480.510 2464.270 ;
        RECT 477.730 2284.690 478.910 2285.870 ;
        RECT 479.330 2284.690 480.510 2285.870 ;
        RECT 477.730 2283.090 478.910 2284.270 ;
        RECT 479.330 2283.090 480.510 2284.270 ;
        RECT 477.730 2104.690 478.910 2105.870 ;
        RECT 479.330 2104.690 480.510 2105.870 ;
        RECT 477.730 2103.090 478.910 2104.270 ;
        RECT 479.330 2103.090 480.510 2104.270 ;
        RECT 477.730 1924.690 478.910 1925.870 ;
        RECT 479.330 1924.690 480.510 1925.870 ;
        RECT 477.730 1923.090 478.910 1924.270 ;
        RECT 479.330 1923.090 480.510 1924.270 ;
        RECT 477.730 1744.690 478.910 1745.870 ;
        RECT 479.330 1744.690 480.510 1745.870 ;
        RECT 477.730 1743.090 478.910 1744.270 ;
        RECT 479.330 1743.090 480.510 1744.270 ;
        RECT 477.730 1564.690 478.910 1565.870 ;
        RECT 479.330 1564.690 480.510 1565.870 ;
        RECT 477.730 1563.090 478.910 1564.270 ;
        RECT 479.330 1563.090 480.510 1564.270 ;
        RECT 477.730 1384.690 478.910 1385.870 ;
        RECT 479.330 1384.690 480.510 1385.870 ;
        RECT 477.730 1383.090 478.910 1384.270 ;
        RECT 479.330 1383.090 480.510 1384.270 ;
        RECT 477.730 1204.690 478.910 1205.870 ;
        RECT 479.330 1204.690 480.510 1205.870 ;
        RECT 477.730 1203.090 478.910 1204.270 ;
        RECT 479.330 1203.090 480.510 1204.270 ;
        RECT 477.730 1024.690 478.910 1025.870 ;
        RECT 479.330 1024.690 480.510 1025.870 ;
        RECT 477.730 1023.090 478.910 1024.270 ;
        RECT 479.330 1023.090 480.510 1024.270 ;
        RECT 657.730 3537.410 658.910 3538.590 ;
        RECT 659.330 3537.410 660.510 3538.590 ;
        RECT 657.730 3535.810 658.910 3536.990 ;
        RECT 659.330 3535.810 660.510 3536.990 ;
        RECT 657.730 3364.690 658.910 3365.870 ;
        RECT 659.330 3364.690 660.510 3365.870 ;
        RECT 657.730 3363.090 658.910 3364.270 ;
        RECT 659.330 3363.090 660.510 3364.270 ;
        RECT 657.730 3184.690 658.910 3185.870 ;
        RECT 659.330 3184.690 660.510 3185.870 ;
        RECT 657.730 3183.090 658.910 3184.270 ;
        RECT 659.330 3183.090 660.510 3184.270 ;
        RECT 657.730 3004.690 658.910 3005.870 ;
        RECT 659.330 3004.690 660.510 3005.870 ;
        RECT 657.730 3003.090 658.910 3004.270 ;
        RECT 659.330 3003.090 660.510 3004.270 ;
        RECT 657.730 2824.690 658.910 2825.870 ;
        RECT 659.330 2824.690 660.510 2825.870 ;
        RECT 657.730 2823.090 658.910 2824.270 ;
        RECT 659.330 2823.090 660.510 2824.270 ;
        RECT 657.730 2644.690 658.910 2645.870 ;
        RECT 659.330 2644.690 660.510 2645.870 ;
        RECT 657.730 2643.090 658.910 2644.270 ;
        RECT 659.330 2643.090 660.510 2644.270 ;
        RECT 657.730 2464.690 658.910 2465.870 ;
        RECT 659.330 2464.690 660.510 2465.870 ;
        RECT 657.730 2463.090 658.910 2464.270 ;
        RECT 659.330 2463.090 660.510 2464.270 ;
        RECT 657.730 2284.690 658.910 2285.870 ;
        RECT 659.330 2284.690 660.510 2285.870 ;
        RECT 657.730 2283.090 658.910 2284.270 ;
        RECT 659.330 2283.090 660.510 2284.270 ;
        RECT 657.730 2104.690 658.910 2105.870 ;
        RECT 659.330 2104.690 660.510 2105.870 ;
        RECT 657.730 2103.090 658.910 2104.270 ;
        RECT 659.330 2103.090 660.510 2104.270 ;
        RECT 657.730 1924.690 658.910 1925.870 ;
        RECT 659.330 1924.690 660.510 1925.870 ;
        RECT 657.730 1923.090 658.910 1924.270 ;
        RECT 659.330 1923.090 660.510 1924.270 ;
        RECT 657.730 1744.690 658.910 1745.870 ;
        RECT 659.330 1744.690 660.510 1745.870 ;
        RECT 657.730 1743.090 658.910 1744.270 ;
        RECT 659.330 1743.090 660.510 1744.270 ;
        RECT 657.730 1564.690 658.910 1565.870 ;
        RECT 659.330 1564.690 660.510 1565.870 ;
        RECT 657.730 1563.090 658.910 1564.270 ;
        RECT 659.330 1563.090 660.510 1564.270 ;
        RECT 657.730 1384.690 658.910 1385.870 ;
        RECT 659.330 1384.690 660.510 1385.870 ;
        RECT 657.730 1383.090 658.910 1384.270 ;
        RECT 659.330 1383.090 660.510 1384.270 ;
        RECT 657.730 1204.690 658.910 1205.870 ;
        RECT 659.330 1204.690 660.510 1205.870 ;
        RECT 657.730 1203.090 658.910 1204.270 ;
        RECT 659.330 1203.090 660.510 1204.270 ;
        RECT 657.730 1024.690 658.910 1025.870 ;
        RECT 659.330 1024.690 660.510 1025.870 ;
        RECT 657.730 1023.090 658.910 1024.270 ;
        RECT 659.330 1023.090 660.510 1024.270 ;
        RECT 837.730 3537.410 838.910 3538.590 ;
        RECT 839.330 3537.410 840.510 3538.590 ;
        RECT 837.730 3535.810 838.910 3536.990 ;
        RECT 839.330 3535.810 840.510 3536.990 ;
        RECT 837.730 3364.690 838.910 3365.870 ;
        RECT 839.330 3364.690 840.510 3365.870 ;
        RECT 837.730 3363.090 838.910 3364.270 ;
        RECT 839.330 3363.090 840.510 3364.270 ;
        RECT 837.730 3184.690 838.910 3185.870 ;
        RECT 839.330 3184.690 840.510 3185.870 ;
        RECT 837.730 3183.090 838.910 3184.270 ;
        RECT 839.330 3183.090 840.510 3184.270 ;
        RECT 837.730 3004.690 838.910 3005.870 ;
        RECT 839.330 3004.690 840.510 3005.870 ;
        RECT 837.730 3003.090 838.910 3004.270 ;
        RECT 839.330 3003.090 840.510 3004.270 ;
        RECT 837.730 2824.690 838.910 2825.870 ;
        RECT 839.330 2824.690 840.510 2825.870 ;
        RECT 837.730 2823.090 838.910 2824.270 ;
        RECT 839.330 2823.090 840.510 2824.270 ;
        RECT 837.730 2644.690 838.910 2645.870 ;
        RECT 839.330 2644.690 840.510 2645.870 ;
        RECT 837.730 2643.090 838.910 2644.270 ;
        RECT 839.330 2643.090 840.510 2644.270 ;
        RECT 837.730 2464.690 838.910 2465.870 ;
        RECT 839.330 2464.690 840.510 2465.870 ;
        RECT 837.730 2463.090 838.910 2464.270 ;
        RECT 839.330 2463.090 840.510 2464.270 ;
        RECT 837.730 2284.690 838.910 2285.870 ;
        RECT 839.330 2284.690 840.510 2285.870 ;
        RECT 837.730 2283.090 838.910 2284.270 ;
        RECT 839.330 2283.090 840.510 2284.270 ;
        RECT 837.730 2104.690 838.910 2105.870 ;
        RECT 839.330 2104.690 840.510 2105.870 ;
        RECT 837.730 2103.090 838.910 2104.270 ;
        RECT 839.330 2103.090 840.510 2104.270 ;
        RECT 837.730 1924.690 838.910 1925.870 ;
        RECT 839.330 1924.690 840.510 1925.870 ;
        RECT 837.730 1923.090 838.910 1924.270 ;
        RECT 839.330 1923.090 840.510 1924.270 ;
        RECT 837.730 1744.690 838.910 1745.870 ;
        RECT 839.330 1744.690 840.510 1745.870 ;
        RECT 837.730 1743.090 838.910 1744.270 ;
        RECT 839.330 1743.090 840.510 1744.270 ;
        RECT 837.730 1564.690 838.910 1565.870 ;
        RECT 839.330 1564.690 840.510 1565.870 ;
        RECT 837.730 1563.090 838.910 1564.270 ;
        RECT 839.330 1563.090 840.510 1564.270 ;
        RECT 837.730 1384.690 838.910 1385.870 ;
        RECT 839.330 1384.690 840.510 1385.870 ;
        RECT 837.730 1383.090 838.910 1384.270 ;
        RECT 839.330 1383.090 840.510 1384.270 ;
        RECT 837.730 1204.690 838.910 1205.870 ;
        RECT 839.330 1204.690 840.510 1205.870 ;
        RECT 837.730 1203.090 838.910 1204.270 ;
        RECT 839.330 1203.090 840.510 1204.270 ;
        RECT 837.730 1024.690 838.910 1025.870 ;
        RECT 839.330 1024.690 840.510 1025.870 ;
        RECT 837.730 1023.090 838.910 1024.270 ;
        RECT 839.330 1023.090 840.510 1024.270 ;
        RECT 1017.730 3537.410 1018.910 3538.590 ;
        RECT 1019.330 3537.410 1020.510 3538.590 ;
        RECT 1017.730 3535.810 1018.910 3536.990 ;
        RECT 1019.330 3535.810 1020.510 3536.990 ;
        RECT 1017.730 3364.690 1018.910 3365.870 ;
        RECT 1019.330 3364.690 1020.510 3365.870 ;
        RECT 1017.730 3363.090 1018.910 3364.270 ;
        RECT 1019.330 3363.090 1020.510 3364.270 ;
        RECT 1017.730 3184.690 1018.910 3185.870 ;
        RECT 1019.330 3184.690 1020.510 3185.870 ;
        RECT 1017.730 3183.090 1018.910 3184.270 ;
        RECT 1019.330 3183.090 1020.510 3184.270 ;
        RECT 1017.730 3004.690 1018.910 3005.870 ;
        RECT 1019.330 3004.690 1020.510 3005.870 ;
        RECT 1017.730 3003.090 1018.910 3004.270 ;
        RECT 1019.330 3003.090 1020.510 3004.270 ;
        RECT 1017.730 2824.690 1018.910 2825.870 ;
        RECT 1019.330 2824.690 1020.510 2825.870 ;
        RECT 1017.730 2823.090 1018.910 2824.270 ;
        RECT 1019.330 2823.090 1020.510 2824.270 ;
        RECT 1017.730 2644.690 1018.910 2645.870 ;
        RECT 1019.330 2644.690 1020.510 2645.870 ;
        RECT 1017.730 2643.090 1018.910 2644.270 ;
        RECT 1019.330 2643.090 1020.510 2644.270 ;
        RECT 1017.730 2464.690 1018.910 2465.870 ;
        RECT 1019.330 2464.690 1020.510 2465.870 ;
        RECT 1017.730 2463.090 1018.910 2464.270 ;
        RECT 1019.330 2463.090 1020.510 2464.270 ;
        RECT 1017.730 2284.690 1018.910 2285.870 ;
        RECT 1019.330 2284.690 1020.510 2285.870 ;
        RECT 1017.730 2283.090 1018.910 2284.270 ;
        RECT 1019.330 2283.090 1020.510 2284.270 ;
        RECT 1017.730 2104.690 1018.910 2105.870 ;
        RECT 1019.330 2104.690 1020.510 2105.870 ;
        RECT 1017.730 2103.090 1018.910 2104.270 ;
        RECT 1019.330 2103.090 1020.510 2104.270 ;
        RECT 1017.730 1924.690 1018.910 1925.870 ;
        RECT 1019.330 1924.690 1020.510 1925.870 ;
        RECT 1017.730 1923.090 1018.910 1924.270 ;
        RECT 1019.330 1923.090 1020.510 1924.270 ;
        RECT 1017.730 1744.690 1018.910 1745.870 ;
        RECT 1019.330 1744.690 1020.510 1745.870 ;
        RECT 1017.730 1743.090 1018.910 1744.270 ;
        RECT 1019.330 1743.090 1020.510 1744.270 ;
        RECT 1017.730 1564.690 1018.910 1565.870 ;
        RECT 1019.330 1564.690 1020.510 1565.870 ;
        RECT 1017.730 1563.090 1018.910 1564.270 ;
        RECT 1019.330 1563.090 1020.510 1564.270 ;
        RECT 1017.730 1384.690 1018.910 1385.870 ;
        RECT 1019.330 1384.690 1020.510 1385.870 ;
        RECT 1017.730 1383.090 1018.910 1384.270 ;
        RECT 1019.330 1383.090 1020.510 1384.270 ;
        RECT 1017.730 1204.690 1018.910 1205.870 ;
        RECT 1019.330 1204.690 1020.510 1205.870 ;
        RECT 1017.730 1203.090 1018.910 1204.270 ;
        RECT 1019.330 1203.090 1020.510 1204.270 ;
        RECT 1017.730 1024.690 1018.910 1025.870 ;
        RECT 1019.330 1024.690 1020.510 1025.870 ;
        RECT 1017.730 1023.090 1018.910 1024.270 ;
        RECT 1019.330 1023.090 1020.510 1024.270 ;
        RECT 1197.730 3537.410 1198.910 3538.590 ;
        RECT 1199.330 3537.410 1200.510 3538.590 ;
        RECT 1197.730 3535.810 1198.910 3536.990 ;
        RECT 1199.330 3535.810 1200.510 3536.990 ;
        RECT 1197.730 3364.690 1198.910 3365.870 ;
        RECT 1199.330 3364.690 1200.510 3365.870 ;
        RECT 1197.730 3363.090 1198.910 3364.270 ;
        RECT 1199.330 3363.090 1200.510 3364.270 ;
        RECT 1197.730 3184.690 1198.910 3185.870 ;
        RECT 1199.330 3184.690 1200.510 3185.870 ;
        RECT 1197.730 3183.090 1198.910 3184.270 ;
        RECT 1199.330 3183.090 1200.510 3184.270 ;
        RECT 1197.730 3004.690 1198.910 3005.870 ;
        RECT 1199.330 3004.690 1200.510 3005.870 ;
        RECT 1197.730 3003.090 1198.910 3004.270 ;
        RECT 1199.330 3003.090 1200.510 3004.270 ;
        RECT 1197.730 2824.690 1198.910 2825.870 ;
        RECT 1199.330 2824.690 1200.510 2825.870 ;
        RECT 1197.730 2823.090 1198.910 2824.270 ;
        RECT 1199.330 2823.090 1200.510 2824.270 ;
        RECT 1197.730 2644.690 1198.910 2645.870 ;
        RECT 1199.330 2644.690 1200.510 2645.870 ;
        RECT 1197.730 2643.090 1198.910 2644.270 ;
        RECT 1199.330 2643.090 1200.510 2644.270 ;
        RECT 1197.730 2464.690 1198.910 2465.870 ;
        RECT 1199.330 2464.690 1200.510 2465.870 ;
        RECT 1197.730 2463.090 1198.910 2464.270 ;
        RECT 1199.330 2463.090 1200.510 2464.270 ;
        RECT 1197.730 2284.690 1198.910 2285.870 ;
        RECT 1199.330 2284.690 1200.510 2285.870 ;
        RECT 1197.730 2283.090 1198.910 2284.270 ;
        RECT 1199.330 2283.090 1200.510 2284.270 ;
        RECT 1197.730 2104.690 1198.910 2105.870 ;
        RECT 1199.330 2104.690 1200.510 2105.870 ;
        RECT 1197.730 2103.090 1198.910 2104.270 ;
        RECT 1199.330 2103.090 1200.510 2104.270 ;
        RECT 1197.730 1924.690 1198.910 1925.870 ;
        RECT 1199.330 1924.690 1200.510 1925.870 ;
        RECT 1197.730 1923.090 1198.910 1924.270 ;
        RECT 1199.330 1923.090 1200.510 1924.270 ;
        RECT 1197.730 1744.690 1198.910 1745.870 ;
        RECT 1199.330 1744.690 1200.510 1745.870 ;
        RECT 1197.730 1743.090 1198.910 1744.270 ;
        RECT 1199.330 1743.090 1200.510 1744.270 ;
        RECT 1197.730 1564.690 1198.910 1565.870 ;
        RECT 1199.330 1564.690 1200.510 1565.870 ;
        RECT 1197.730 1563.090 1198.910 1564.270 ;
        RECT 1199.330 1563.090 1200.510 1564.270 ;
        RECT 1197.730 1384.690 1198.910 1385.870 ;
        RECT 1199.330 1384.690 1200.510 1385.870 ;
        RECT 1197.730 1383.090 1198.910 1384.270 ;
        RECT 1199.330 1383.090 1200.510 1384.270 ;
        RECT 1197.730 1204.690 1198.910 1205.870 ;
        RECT 1199.330 1204.690 1200.510 1205.870 ;
        RECT 1197.730 1203.090 1198.910 1204.270 ;
        RECT 1199.330 1203.090 1200.510 1204.270 ;
        RECT 1197.730 1024.690 1198.910 1025.870 ;
        RECT 1199.330 1024.690 1200.510 1025.870 ;
        RECT 1197.730 1023.090 1198.910 1024.270 ;
        RECT 1199.330 1023.090 1200.510 1024.270 ;
        RECT 117.730 844.690 118.910 845.870 ;
        RECT 119.330 844.690 120.510 845.870 ;
        RECT 117.730 843.090 118.910 844.270 ;
        RECT 119.330 843.090 120.510 844.270 ;
        RECT 117.730 664.690 118.910 665.870 ;
        RECT 119.330 664.690 120.510 665.870 ;
        RECT 117.730 663.090 118.910 664.270 ;
        RECT 119.330 663.090 120.510 664.270 ;
        RECT 117.730 484.690 118.910 485.870 ;
        RECT 119.330 484.690 120.510 485.870 ;
        RECT 117.730 483.090 118.910 484.270 ;
        RECT 119.330 483.090 120.510 484.270 ;
        RECT 1197.730 844.690 1198.910 845.870 ;
        RECT 1199.330 844.690 1200.510 845.870 ;
        RECT 1197.730 843.090 1198.910 844.270 ;
        RECT 1199.330 843.090 1200.510 844.270 ;
        RECT 1197.730 664.690 1198.910 665.870 ;
        RECT 1199.330 664.690 1200.510 665.870 ;
        RECT 1197.730 663.090 1198.910 664.270 ;
        RECT 1199.330 663.090 1200.510 664.270 ;
        RECT 1197.730 484.690 1198.910 485.870 ;
        RECT 1199.330 484.690 1200.510 485.870 ;
        RECT 1197.730 483.090 1198.910 484.270 ;
        RECT 1199.330 483.090 1200.510 484.270 ;
        RECT 117.730 304.690 118.910 305.870 ;
        RECT 119.330 304.690 120.510 305.870 ;
        RECT 117.730 303.090 118.910 304.270 ;
        RECT 119.330 303.090 120.510 304.270 ;
        RECT 117.730 124.690 118.910 125.870 ;
        RECT 119.330 124.690 120.510 125.870 ;
        RECT 117.730 123.090 118.910 124.270 ;
        RECT 119.330 123.090 120.510 124.270 ;
        RECT 117.730 -17.310 118.910 -16.130 ;
        RECT 119.330 -17.310 120.510 -16.130 ;
        RECT 117.730 -18.910 118.910 -17.730 ;
        RECT 119.330 -18.910 120.510 -17.730 ;
        RECT 297.730 304.690 298.910 305.870 ;
        RECT 299.330 304.690 300.510 305.870 ;
        RECT 297.730 303.090 298.910 304.270 ;
        RECT 299.330 303.090 300.510 304.270 ;
        RECT 297.730 124.690 298.910 125.870 ;
        RECT 299.330 124.690 300.510 125.870 ;
        RECT 297.730 123.090 298.910 124.270 ;
        RECT 299.330 123.090 300.510 124.270 ;
        RECT 297.730 -17.310 298.910 -16.130 ;
        RECT 299.330 -17.310 300.510 -16.130 ;
        RECT 297.730 -18.910 298.910 -17.730 ;
        RECT 299.330 -18.910 300.510 -17.730 ;
        RECT 477.730 304.690 478.910 305.870 ;
        RECT 479.330 304.690 480.510 305.870 ;
        RECT 477.730 303.090 478.910 304.270 ;
        RECT 479.330 303.090 480.510 304.270 ;
        RECT 477.730 124.690 478.910 125.870 ;
        RECT 479.330 124.690 480.510 125.870 ;
        RECT 477.730 123.090 478.910 124.270 ;
        RECT 479.330 123.090 480.510 124.270 ;
        RECT 477.730 -17.310 478.910 -16.130 ;
        RECT 479.330 -17.310 480.510 -16.130 ;
        RECT 477.730 -18.910 478.910 -17.730 ;
        RECT 479.330 -18.910 480.510 -17.730 ;
        RECT 657.730 304.690 658.910 305.870 ;
        RECT 659.330 304.690 660.510 305.870 ;
        RECT 657.730 303.090 658.910 304.270 ;
        RECT 659.330 303.090 660.510 304.270 ;
        RECT 657.730 124.690 658.910 125.870 ;
        RECT 659.330 124.690 660.510 125.870 ;
        RECT 657.730 123.090 658.910 124.270 ;
        RECT 659.330 123.090 660.510 124.270 ;
        RECT 657.730 -17.310 658.910 -16.130 ;
        RECT 659.330 -17.310 660.510 -16.130 ;
        RECT 657.730 -18.910 658.910 -17.730 ;
        RECT 659.330 -18.910 660.510 -17.730 ;
        RECT 837.730 304.690 838.910 305.870 ;
        RECT 839.330 304.690 840.510 305.870 ;
        RECT 837.730 303.090 838.910 304.270 ;
        RECT 839.330 303.090 840.510 304.270 ;
        RECT 837.730 124.690 838.910 125.870 ;
        RECT 839.330 124.690 840.510 125.870 ;
        RECT 837.730 123.090 838.910 124.270 ;
        RECT 839.330 123.090 840.510 124.270 ;
        RECT 837.730 -17.310 838.910 -16.130 ;
        RECT 839.330 -17.310 840.510 -16.130 ;
        RECT 837.730 -18.910 838.910 -17.730 ;
        RECT 839.330 -18.910 840.510 -17.730 ;
        RECT 1017.730 304.690 1018.910 305.870 ;
        RECT 1019.330 304.690 1020.510 305.870 ;
        RECT 1017.730 303.090 1018.910 304.270 ;
        RECT 1019.330 303.090 1020.510 304.270 ;
        RECT 1017.730 124.690 1018.910 125.870 ;
        RECT 1019.330 124.690 1020.510 125.870 ;
        RECT 1017.730 123.090 1018.910 124.270 ;
        RECT 1019.330 123.090 1020.510 124.270 ;
        RECT 1017.730 -17.310 1018.910 -16.130 ;
        RECT 1019.330 -17.310 1020.510 -16.130 ;
        RECT 1017.730 -18.910 1018.910 -17.730 ;
        RECT 1019.330 -18.910 1020.510 -17.730 ;
        RECT 1197.730 304.690 1198.910 305.870 ;
        RECT 1199.330 304.690 1200.510 305.870 ;
        RECT 1197.730 303.090 1198.910 304.270 ;
        RECT 1199.330 303.090 1200.510 304.270 ;
        RECT 1197.730 124.690 1198.910 125.870 ;
        RECT 1199.330 124.690 1200.510 125.870 ;
        RECT 1197.730 123.090 1198.910 124.270 ;
        RECT 1199.330 123.090 1200.510 124.270 ;
        RECT 1197.730 -17.310 1198.910 -16.130 ;
        RECT 1199.330 -17.310 1200.510 -16.130 ;
        RECT 1197.730 -18.910 1198.910 -17.730 ;
        RECT 1199.330 -18.910 1200.510 -17.730 ;
        RECT 1377.730 3537.410 1378.910 3538.590 ;
        RECT 1379.330 3537.410 1380.510 3538.590 ;
        RECT 1377.730 3535.810 1378.910 3536.990 ;
        RECT 1379.330 3535.810 1380.510 3536.990 ;
        RECT 1377.730 3364.690 1378.910 3365.870 ;
        RECT 1379.330 3364.690 1380.510 3365.870 ;
        RECT 1377.730 3363.090 1378.910 3364.270 ;
        RECT 1379.330 3363.090 1380.510 3364.270 ;
        RECT 1377.730 3184.690 1378.910 3185.870 ;
        RECT 1379.330 3184.690 1380.510 3185.870 ;
        RECT 1377.730 3183.090 1378.910 3184.270 ;
        RECT 1379.330 3183.090 1380.510 3184.270 ;
        RECT 1377.730 3004.690 1378.910 3005.870 ;
        RECT 1379.330 3004.690 1380.510 3005.870 ;
        RECT 1377.730 3003.090 1378.910 3004.270 ;
        RECT 1379.330 3003.090 1380.510 3004.270 ;
        RECT 1377.730 2824.690 1378.910 2825.870 ;
        RECT 1379.330 2824.690 1380.510 2825.870 ;
        RECT 1377.730 2823.090 1378.910 2824.270 ;
        RECT 1379.330 2823.090 1380.510 2824.270 ;
        RECT 1377.730 2644.690 1378.910 2645.870 ;
        RECT 1379.330 2644.690 1380.510 2645.870 ;
        RECT 1377.730 2643.090 1378.910 2644.270 ;
        RECT 1379.330 2643.090 1380.510 2644.270 ;
        RECT 1377.730 2464.690 1378.910 2465.870 ;
        RECT 1379.330 2464.690 1380.510 2465.870 ;
        RECT 1377.730 2463.090 1378.910 2464.270 ;
        RECT 1379.330 2463.090 1380.510 2464.270 ;
        RECT 1377.730 2284.690 1378.910 2285.870 ;
        RECT 1379.330 2284.690 1380.510 2285.870 ;
        RECT 1377.730 2283.090 1378.910 2284.270 ;
        RECT 1379.330 2283.090 1380.510 2284.270 ;
        RECT 1377.730 2104.690 1378.910 2105.870 ;
        RECT 1379.330 2104.690 1380.510 2105.870 ;
        RECT 1377.730 2103.090 1378.910 2104.270 ;
        RECT 1379.330 2103.090 1380.510 2104.270 ;
        RECT 1377.730 1924.690 1378.910 1925.870 ;
        RECT 1379.330 1924.690 1380.510 1925.870 ;
        RECT 1377.730 1923.090 1378.910 1924.270 ;
        RECT 1379.330 1923.090 1380.510 1924.270 ;
        RECT 1377.730 1744.690 1378.910 1745.870 ;
        RECT 1379.330 1744.690 1380.510 1745.870 ;
        RECT 1377.730 1743.090 1378.910 1744.270 ;
        RECT 1379.330 1743.090 1380.510 1744.270 ;
        RECT 1377.730 1564.690 1378.910 1565.870 ;
        RECT 1379.330 1564.690 1380.510 1565.870 ;
        RECT 1377.730 1563.090 1378.910 1564.270 ;
        RECT 1379.330 1563.090 1380.510 1564.270 ;
        RECT 1377.730 1384.690 1378.910 1385.870 ;
        RECT 1379.330 1384.690 1380.510 1385.870 ;
        RECT 1377.730 1383.090 1378.910 1384.270 ;
        RECT 1379.330 1383.090 1380.510 1384.270 ;
        RECT 1377.730 1204.690 1378.910 1205.870 ;
        RECT 1379.330 1204.690 1380.510 1205.870 ;
        RECT 1377.730 1203.090 1378.910 1204.270 ;
        RECT 1379.330 1203.090 1380.510 1204.270 ;
        RECT 1377.730 1024.690 1378.910 1025.870 ;
        RECT 1379.330 1024.690 1380.510 1025.870 ;
        RECT 1377.730 1023.090 1378.910 1024.270 ;
        RECT 1379.330 1023.090 1380.510 1024.270 ;
        RECT 1377.730 844.690 1378.910 845.870 ;
        RECT 1379.330 844.690 1380.510 845.870 ;
        RECT 1377.730 843.090 1378.910 844.270 ;
        RECT 1379.330 843.090 1380.510 844.270 ;
        RECT 1377.730 664.690 1378.910 665.870 ;
        RECT 1379.330 664.690 1380.510 665.870 ;
        RECT 1377.730 663.090 1378.910 664.270 ;
        RECT 1379.330 663.090 1380.510 664.270 ;
        RECT 1377.730 484.690 1378.910 485.870 ;
        RECT 1379.330 484.690 1380.510 485.870 ;
        RECT 1377.730 483.090 1378.910 484.270 ;
        RECT 1379.330 483.090 1380.510 484.270 ;
        RECT 1377.730 304.690 1378.910 305.870 ;
        RECT 1379.330 304.690 1380.510 305.870 ;
        RECT 1377.730 303.090 1378.910 304.270 ;
        RECT 1379.330 303.090 1380.510 304.270 ;
        RECT 1377.730 124.690 1378.910 125.870 ;
        RECT 1379.330 124.690 1380.510 125.870 ;
        RECT 1377.730 123.090 1378.910 124.270 ;
        RECT 1379.330 123.090 1380.510 124.270 ;
        RECT 1377.730 -17.310 1378.910 -16.130 ;
        RECT 1379.330 -17.310 1380.510 -16.130 ;
        RECT 1377.730 -18.910 1378.910 -17.730 ;
        RECT 1379.330 -18.910 1380.510 -17.730 ;
        RECT 1557.730 3537.410 1558.910 3538.590 ;
        RECT 1559.330 3537.410 1560.510 3538.590 ;
        RECT 1557.730 3535.810 1558.910 3536.990 ;
        RECT 1559.330 3535.810 1560.510 3536.990 ;
        RECT 1557.730 3364.690 1558.910 3365.870 ;
        RECT 1559.330 3364.690 1560.510 3365.870 ;
        RECT 1557.730 3363.090 1558.910 3364.270 ;
        RECT 1559.330 3363.090 1560.510 3364.270 ;
        RECT 1557.730 3184.690 1558.910 3185.870 ;
        RECT 1559.330 3184.690 1560.510 3185.870 ;
        RECT 1557.730 3183.090 1558.910 3184.270 ;
        RECT 1559.330 3183.090 1560.510 3184.270 ;
        RECT 1557.730 3004.690 1558.910 3005.870 ;
        RECT 1559.330 3004.690 1560.510 3005.870 ;
        RECT 1557.730 3003.090 1558.910 3004.270 ;
        RECT 1559.330 3003.090 1560.510 3004.270 ;
        RECT 1557.730 2824.690 1558.910 2825.870 ;
        RECT 1559.330 2824.690 1560.510 2825.870 ;
        RECT 1557.730 2823.090 1558.910 2824.270 ;
        RECT 1559.330 2823.090 1560.510 2824.270 ;
        RECT 1557.730 2644.690 1558.910 2645.870 ;
        RECT 1559.330 2644.690 1560.510 2645.870 ;
        RECT 1557.730 2643.090 1558.910 2644.270 ;
        RECT 1559.330 2643.090 1560.510 2644.270 ;
        RECT 1557.730 2464.690 1558.910 2465.870 ;
        RECT 1559.330 2464.690 1560.510 2465.870 ;
        RECT 1557.730 2463.090 1558.910 2464.270 ;
        RECT 1559.330 2463.090 1560.510 2464.270 ;
        RECT 1557.730 2284.690 1558.910 2285.870 ;
        RECT 1559.330 2284.690 1560.510 2285.870 ;
        RECT 1557.730 2283.090 1558.910 2284.270 ;
        RECT 1559.330 2283.090 1560.510 2284.270 ;
        RECT 1557.730 2104.690 1558.910 2105.870 ;
        RECT 1559.330 2104.690 1560.510 2105.870 ;
        RECT 1557.730 2103.090 1558.910 2104.270 ;
        RECT 1559.330 2103.090 1560.510 2104.270 ;
        RECT 1557.730 1924.690 1558.910 1925.870 ;
        RECT 1559.330 1924.690 1560.510 1925.870 ;
        RECT 1557.730 1923.090 1558.910 1924.270 ;
        RECT 1559.330 1923.090 1560.510 1924.270 ;
        RECT 1557.730 1744.690 1558.910 1745.870 ;
        RECT 1559.330 1744.690 1560.510 1745.870 ;
        RECT 1557.730 1743.090 1558.910 1744.270 ;
        RECT 1559.330 1743.090 1560.510 1744.270 ;
        RECT 1557.730 1564.690 1558.910 1565.870 ;
        RECT 1559.330 1564.690 1560.510 1565.870 ;
        RECT 1557.730 1563.090 1558.910 1564.270 ;
        RECT 1559.330 1563.090 1560.510 1564.270 ;
        RECT 1557.730 1384.690 1558.910 1385.870 ;
        RECT 1559.330 1384.690 1560.510 1385.870 ;
        RECT 1557.730 1383.090 1558.910 1384.270 ;
        RECT 1559.330 1383.090 1560.510 1384.270 ;
        RECT 1557.730 1204.690 1558.910 1205.870 ;
        RECT 1559.330 1204.690 1560.510 1205.870 ;
        RECT 1557.730 1203.090 1558.910 1204.270 ;
        RECT 1559.330 1203.090 1560.510 1204.270 ;
        RECT 1557.730 1024.690 1558.910 1025.870 ;
        RECT 1559.330 1024.690 1560.510 1025.870 ;
        RECT 1557.730 1023.090 1558.910 1024.270 ;
        RECT 1559.330 1023.090 1560.510 1024.270 ;
        RECT 1557.730 844.690 1558.910 845.870 ;
        RECT 1559.330 844.690 1560.510 845.870 ;
        RECT 1557.730 843.090 1558.910 844.270 ;
        RECT 1559.330 843.090 1560.510 844.270 ;
        RECT 1557.730 664.690 1558.910 665.870 ;
        RECT 1559.330 664.690 1560.510 665.870 ;
        RECT 1557.730 663.090 1558.910 664.270 ;
        RECT 1559.330 663.090 1560.510 664.270 ;
        RECT 1557.730 484.690 1558.910 485.870 ;
        RECT 1559.330 484.690 1560.510 485.870 ;
        RECT 1557.730 483.090 1558.910 484.270 ;
        RECT 1559.330 483.090 1560.510 484.270 ;
        RECT 1557.730 304.690 1558.910 305.870 ;
        RECT 1559.330 304.690 1560.510 305.870 ;
        RECT 1557.730 303.090 1558.910 304.270 ;
        RECT 1559.330 303.090 1560.510 304.270 ;
        RECT 1557.730 124.690 1558.910 125.870 ;
        RECT 1559.330 124.690 1560.510 125.870 ;
        RECT 1557.730 123.090 1558.910 124.270 ;
        RECT 1559.330 123.090 1560.510 124.270 ;
        RECT 1557.730 -17.310 1558.910 -16.130 ;
        RECT 1559.330 -17.310 1560.510 -16.130 ;
        RECT 1557.730 -18.910 1558.910 -17.730 ;
        RECT 1559.330 -18.910 1560.510 -17.730 ;
        RECT 1737.730 3537.410 1738.910 3538.590 ;
        RECT 1739.330 3537.410 1740.510 3538.590 ;
        RECT 1737.730 3535.810 1738.910 3536.990 ;
        RECT 1739.330 3535.810 1740.510 3536.990 ;
        RECT 1737.730 3364.690 1738.910 3365.870 ;
        RECT 1739.330 3364.690 1740.510 3365.870 ;
        RECT 1737.730 3363.090 1738.910 3364.270 ;
        RECT 1739.330 3363.090 1740.510 3364.270 ;
        RECT 1737.730 3184.690 1738.910 3185.870 ;
        RECT 1739.330 3184.690 1740.510 3185.870 ;
        RECT 1737.730 3183.090 1738.910 3184.270 ;
        RECT 1739.330 3183.090 1740.510 3184.270 ;
        RECT 1737.730 3004.690 1738.910 3005.870 ;
        RECT 1739.330 3004.690 1740.510 3005.870 ;
        RECT 1737.730 3003.090 1738.910 3004.270 ;
        RECT 1739.330 3003.090 1740.510 3004.270 ;
        RECT 1737.730 2824.690 1738.910 2825.870 ;
        RECT 1739.330 2824.690 1740.510 2825.870 ;
        RECT 1737.730 2823.090 1738.910 2824.270 ;
        RECT 1739.330 2823.090 1740.510 2824.270 ;
        RECT 1737.730 2644.690 1738.910 2645.870 ;
        RECT 1739.330 2644.690 1740.510 2645.870 ;
        RECT 1737.730 2643.090 1738.910 2644.270 ;
        RECT 1739.330 2643.090 1740.510 2644.270 ;
        RECT 1737.730 2464.690 1738.910 2465.870 ;
        RECT 1739.330 2464.690 1740.510 2465.870 ;
        RECT 1737.730 2463.090 1738.910 2464.270 ;
        RECT 1739.330 2463.090 1740.510 2464.270 ;
        RECT 1737.730 2284.690 1738.910 2285.870 ;
        RECT 1739.330 2284.690 1740.510 2285.870 ;
        RECT 1737.730 2283.090 1738.910 2284.270 ;
        RECT 1739.330 2283.090 1740.510 2284.270 ;
        RECT 1737.730 2104.690 1738.910 2105.870 ;
        RECT 1739.330 2104.690 1740.510 2105.870 ;
        RECT 1737.730 2103.090 1738.910 2104.270 ;
        RECT 1739.330 2103.090 1740.510 2104.270 ;
        RECT 1737.730 1924.690 1738.910 1925.870 ;
        RECT 1739.330 1924.690 1740.510 1925.870 ;
        RECT 1737.730 1923.090 1738.910 1924.270 ;
        RECT 1739.330 1923.090 1740.510 1924.270 ;
        RECT 1737.730 1744.690 1738.910 1745.870 ;
        RECT 1739.330 1744.690 1740.510 1745.870 ;
        RECT 1737.730 1743.090 1738.910 1744.270 ;
        RECT 1739.330 1743.090 1740.510 1744.270 ;
        RECT 1737.730 1564.690 1738.910 1565.870 ;
        RECT 1739.330 1564.690 1740.510 1565.870 ;
        RECT 1737.730 1563.090 1738.910 1564.270 ;
        RECT 1739.330 1563.090 1740.510 1564.270 ;
        RECT 1737.730 1384.690 1738.910 1385.870 ;
        RECT 1739.330 1384.690 1740.510 1385.870 ;
        RECT 1737.730 1383.090 1738.910 1384.270 ;
        RECT 1739.330 1383.090 1740.510 1384.270 ;
        RECT 1737.730 1204.690 1738.910 1205.870 ;
        RECT 1739.330 1204.690 1740.510 1205.870 ;
        RECT 1737.730 1203.090 1738.910 1204.270 ;
        RECT 1739.330 1203.090 1740.510 1204.270 ;
        RECT 1737.730 1024.690 1738.910 1025.870 ;
        RECT 1739.330 1024.690 1740.510 1025.870 ;
        RECT 1737.730 1023.090 1738.910 1024.270 ;
        RECT 1739.330 1023.090 1740.510 1024.270 ;
        RECT 1737.730 844.690 1738.910 845.870 ;
        RECT 1739.330 844.690 1740.510 845.870 ;
        RECT 1737.730 843.090 1738.910 844.270 ;
        RECT 1739.330 843.090 1740.510 844.270 ;
        RECT 1737.730 664.690 1738.910 665.870 ;
        RECT 1739.330 664.690 1740.510 665.870 ;
        RECT 1737.730 663.090 1738.910 664.270 ;
        RECT 1739.330 663.090 1740.510 664.270 ;
        RECT 1737.730 484.690 1738.910 485.870 ;
        RECT 1739.330 484.690 1740.510 485.870 ;
        RECT 1737.730 483.090 1738.910 484.270 ;
        RECT 1739.330 483.090 1740.510 484.270 ;
        RECT 1737.730 304.690 1738.910 305.870 ;
        RECT 1739.330 304.690 1740.510 305.870 ;
        RECT 1737.730 303.090 1738.910 304.270 ;
        RECT 1739.330 303.090 1740.510 304.270 ;
        RECT 1737.730 124.690 1738.910 125.870 ;
        RECT 1739.330 124.690 1740.510 125.870 ;
        RECT 1737.730 123.090 1738.910 124.270 ;
        RECT 1739.330 123.090 1740.510 124.270 ;
        RECT 1737.730 -17.310 1738.910 -16.130 ;
        RECT 1739.330 -17.310 1740.510 -16.130 ;
        RECT 1737.730 -18.910 1738.910 -17.730 ;
        RECT 1739.330 -18.910 1740.510 -17.730 ;
        RECT 1917.730 3537.410 1918.910 3538.590 ;
        RECT 1919.330 3537.410 1920.510 3538.590 ;
        RECT 1917.730 3535.810 1918.910 3536.990 ;
        RECT 1919.330 3535.810 1920.510 3536.990 ;
        RECT 1917.730 3364.690 1918.910 3365.870 ;
        RECT 1919.330 3364.690 1920.510 3365.870 ;
        RECT 1917.730 3363.090 1918.910 3364.270 ;
        RECT 1919.330 3363.090 1920.510 3364.270 ;
        RECT 1917.730 3184.690 1918.910 3185.870 ;
        RECT 1919.330 3184.690 1920.510 3185.870 ;
        RECT 1917.730 3183.090 1918.910 3184.270 ;
        RECT 1919.330 3183.090 1920.510 3184.270 ;
        RECT 1917.730 3004.690 1918.910 3005.870 ;
        RECT 1919.330 3004.690 1920.510 3005.870 ;
        RECT 1917.730 3003.090 1918.910 3004.270 ;
        RECT 1919.330 3003.090 1920.510 3004.270 ;
        RECT 1917.730 2824.690 1918.910 2825.870 ;
        RECT 1919.330 2824.690 1920.510 2825.870 ;
        RECT 1917.730 2823.090 1918.910 2824.270 ;
        RECT 1919.330 2823.090 1920.510 2824.270 ;
        RECT 1917.730 2644.690 1918.910 2645.870 ;
        RECT 1919.330 2644.690 1920.510 2645.870 ;
        RECT 1917.730 2643.090 1918.910 2644.270 ;
        RECT 1919.330 2643.090 1920.510 2644.270 ;
        RECT 1917.730 2464.690 1918.910 2465.870 ;
        RECT 1919.330 2464.690 1920.510 2465.870 ;
        RECT 1917.730 2463.090 1918.910 2464.270 ;
        RECT 1919.330 2463.090 1920.510 2464.270 ;
        RECT 1917.730 2284.690 1918.910 2285.870 ;
        RECT 1919.330 2284.690 1920.510 2285.870 ;
        RECT 1917.730 2283.090 1918.910 2284.270 ;
        RECT 1919.330 2283.090 1920.510 2284.270 ;
        RECT 1917.730 2104.690 1918.910 2105.870 ;
        RECT 1919.330 2104.690 1920.510 2105.870 ;
        RECT 1917.730 2103.090 1918.910 2104.270 ;
        RECT 1919.330 2103.090 1920.510 2104.270 ;
        RECT 1917.730 1924.690 1918.910 1925.870 ;
        RECT 1919.330 1924.690 1920.510 1925.870 ;
        RECT 1917.730 1923.090 1918.910 1924.270 ;
        RECT 1919.330 1923.090 1920.510 1924.270 ;
        RECT 1917.730 1744.690 1918.910 1745.870 ;
        RECT 1919.330 1744.690 1920.510 1745.870 ;
        RECT 1917.730 1743.090 1918.910 1744.270 ;
        RECT 1919.330 1743.090 1920.510 1744.270 ;
        RECT 1917.730 1564.690 1918.910 1565.870 ;
        RECT 1919.330 1564.690 1920.510 1565.870 ;
        RECT 1917.730 1563.090 1918.910 1564.270 ;
        RECT 1919.330 1563.090 1920.510 1564.270 ;
        RECT 1917.730 1384.690 1918.910 1385.870 ;
        RECT 1919.330 1384.690 1920.510 1385.870 ;
        RECT 1917.730 1383.090 1918.910 1384.270 ;
        RECT 1919.330 1383.090 1920.510 1384.270 ;
        RECT 1917.730 1204.690 1918.910 1205.870 ;
        RECT 1919.330 1204.690 1920.510 1205.870 ;
        RECT 1917.730 1203.090 1918.910 1204.270 ;
        RECT 1919.330 1203.090 1920.510 1204.270 ;
        RECT 1917.730 1024.690 1918.910 1025.870 ;
        RECT 1919.330 1024.690 1920.510 1025.870 ;
        RECT 1917.730 1023.090 1918.910 1024.270 ;
        RECT 1919.330 1023.090 1920.510 1024.270 ;
        RECT 1917.730 844.690 1918.910 845.870 ;
        RECT 1919.330 844.690 1920.510 845.870 ;
        RECT 1917.730 843.090 1918.910 844.270 ;
        RECT 1919.330 843.090 1920.510 844.270 ;
        RECT 1917.730 664.690 1918.910 665.870 ;
        RECT 1919.330 664.690 1920.510 665.870 ;
        RECT 1917.730 663.090 1918.910 664.270 ;
        RECT 1919.330 663.090 1920.510 664.270 ;
        RECT 1917.730 484.690 1918.910 485.870 ;
        RECT 1919.330 484.690 1920.510 485.870 ;
        RECT 1917.730 483.090 1918.910 484.270 ;
        RECT 1919.330 483.090 1920.510 484.270 ;
        RECT 1917.730 304.690 1918.910 305.870 ;
        RECT 1919.330 304.690 1920.510 305.870 ;
        RECT 1917.730 303.090 1918.910 304.270 ;
        RECT 1919.330 303.090 1920.510 304.270 ;
        RECT 1917.730 124.690 1918.910 125.870 ;
        RECT 1919.330 124.690 1920.510 125.870 ;
        RECT 1917.730 123.090 1918.910 124.270 ;
        RECT 1919.330 123.090 1920.510 124.270 ;
        RECT 1917.730 -17.310 1918.910 -16.130 ;
        RECT 1919.330 -17.310 1920.510 -16.130 ;
        RECT 1917.730 -18.910 1918.910 -17.730 ;
        RECT 1919.330 -18.910 1920.510 -17.730 ;
        RECT 2097.730 3537.410 2098.910 3538.590 ;
        RECT 2099.330 3537.410 2100.510 3538.590 ;
        RECT 2097.730 3535.810 2098.910 3536.990 ;
        RECT 2099.330 3535.810 2100.510 3536.990 ;
        RECT 2097.730 3364.690 2098.910 3365.870 ;
        RECT 2099.330 3364.690 2100.510 3365.870 ;
        RECT 2097.730 3363.090 2098.910 3364.270 ;
        RECT 2099.330 3363.090 2100.510 3364.270 ;
        RECT 2097.730 3184.690 2098.910 3185.870 ;
        RECT 2099.330 3184.690 2100.510 3185.870 ;
        RECT 2097.730 3183.090 2098.910 3184.270 ;
        RECT 2099.330 3183.090 2100.510 3184.270 ;
        RECT 2097.730 3004.690 2098.910 3005.870 ;
        RECT 2099.330 3004.690 2100.510 3005.870 ;
        RECT 2097.730 3003.090 2098.910 3004.270 ;
        RECT 2099.330 3003.090 2100.510 3004.270 ;
        RECT 2097.730 2824.690 2098.910 2825.870 ;
        RECT 2099.330 2824.690 2100.510 2825.870 ;
        RECT 2097.730 2823.090 2098.910 2824.270 ;
        RECT 2099.330 2823.090 2100.510 2824.270 ;
        RECT 2097.730 2644.690 2098.910 2645.870 ;
        RECT 2099.330 2644.690 2100.510 2645.870 ;
        RECT 2097.730 2643.090 2098.910 2644.270 ;
        RECT 2099.330 2643.090 2100.510 2644.270 ;
        RECT 2097.730 2464.690 2098.910 2465.870 ;
        RECT 2099.330 2464.690 2100.510 2465.870 ;
        RECT 2097.730 2463.090 2098.910 2464.270 ;
        RECT 2099.330 2463.090 2100.510 2464.270 ;
        RECT 2097.730 2284.690 2098.910 2285.870 ;
        RECT 2099.330 2284.690 2100.510 2285.870 ;
        RECT 2097.730 2283.090 2098.910 2284.270 ;
        RECT 2099.330 2283.090 2100.510 2284.270 ;
        RECT 2097.730 2104.690 2098.910 2105.870 ;
        RECT 2099.330 2104.690 2100.510 2105.870 ;
        RECT 2097.730 2103.090 2098.910 2104.270 ;
        RECT 2099.330 2103.090 2100.510 2104.270 ;
        RECT 2097.730 1924.690 2098.910 1925.870 ;
        RECT 2099.330 1924.690 2100.510 1925.870 ;
        RECT 2097.730 1923.090 2098.910 1924.270 ;
        RECT 2099.330 1923.090 2100.510 1924.270 ;
        RECT 2097.730 1744.690 2098.910 1745.870 ;
        RECT 2099.330 1744.690 2100.510 1745.870 ;
        RECT 2097.730 1743.090 2098.910 1744.270 ;
        RECT 2099.330 1743.090 2100.510 1744.270 ;
        RECT 2097.730 1564.690 2098.910 1565.870 ;
        RECT 2099.330 1564.690 2100.510 1565.870 ;
        RECT 2097.730 1563.090 2098.910 1564.270 ;
        RECT 2099.330 1563.090 2100.510 1564.270 ;
        RECT 2097.730 1384.690 2098.910 1385.870 ;
        RECT 2099.330 1384.690 2100.510 1385.870 ;
        RECT 2097.730 1383.090 2098.910 1384.270 ;
        RECT 2099.330 1383.090 2100.510 1384.270 ;
        RECT 2097.730 1204.690 2098.910 1205.870 ;
        RECT 2099.330 1204.690 2100.510 1205.870 ;
        RECT 2097.730 1203.090 2098.910 1204.270 ;
        RECT 2099.330 1203.090 2100.510 1204.270 ;
        RECT 2097.730 1024.690 2098.910 1025.870 ;
        RECT 2099.330 1024.690 2100.510 1025.870 ;
        RECT 2097.730 1023.090 2098.910 1024.270 ;
        RECT 2099.330 1023.090 2100.510 1024.270 ;
        RECT 2097.730 844.690 2098.910 845.870 ;
        RECT 2099.330 844.690 2100.510 845.870 ;
        RECT 2097.730 843.090 2098.910 844.270 ;
        RECT 2099.330 843.090 2100.510 844.270 ;
        RECT 2097.730 664.690 2098.910 665.870 ;
        RECT 2099.330 664.690 2100.510 665.870 ;
        RECT 2097.730 663.090 2098.910 664.270 ;
        RECT 2099.330 663.090 2100.510 664.270 ;
        RECT 2097.730 484.690 2098.910 485.870 ;
        RECT 2099.330 484.690 2100.510 485.870 ;
        RECT 2097.730 483.090 2098.910 484.270 ;
        RECT 2099.330 483.090 2100.510 484.270 ;
        RECT 2097.730 304.690 2098.910 305.870 ;
        RECT 2099.330 304.690 2100.510 305.870 ;
        RECT 2097.730 303.090 2098.910 304.270 ;
        RECT 2099.330 303.090 2100.510 304.270 ;
        RECT 2097.730 124.690 2098.910 125.870 ;
        RECT 2099.330 124.690 2100.510 125.870 ;
        RECT 2097.730 123.090 2098.910 124.270 ;
        RECT 2099.330 123.090 2100.510 124.270 ;
        RECT 2097.730 -17.310 2098.910 -16.130 ;
        RECT 2099.330 -17.310 2100.510 -16.130 ;
        RECT 2097.730 -18.910 2098.910 -17.730 ;
        RECT 2099.330 -18.910 2100.510 -17.730 ;
        RECT 2277.730 3537.410 2278.910 3538.590 ;
        RECT 2279.330 3537.410 2280.510 3538.590 ;
        RECT 2277.730 3535.810 2278.910 3536.990 ;
        RECT 2279.330 3535.810 2280.510 3536.990 ;
        RECT 2277.730 3364.690 2278.910 3365.870 ;
        RECT 2279.330 3364.690 2280.510 3365.870 ;
        RECT 2277.730 3363.090 2278.910 3364.270 ;
        RECT 2279.330 3363.090 2280.510 3364.270 ;
        RECT 2277.730 3184.690 2278.910 3185.870 ;
        RECT 2279.330 3184.690 2280.510 3185.870 ;
        RECT 2277.730 3183.090 2278.910 3184.270 ;
        RECT 2279.330 3183.090 2280.510 3184.270 ;
        RECT 2277.730 3004.690 2278.910 3005.870 ;
        RECT 2279.330 3004.690 2280.510 3005.870 ;
        RECT 2277.730 3003.090 2278.910 3004.270 ;
        RECT 2279.330 3003.090 2280.510 3004.270 ;
        RECT 2277.730 2824.690 2278.910 2825.870 ;
        RECT 2279.330 2824.690 2280.510 2825.870 ;
        RECT 2277.730 2823.090 2278.910 2824.270 ;
        RECT 2279.330 2823.090 2280.510 2824.270 ;
        RECT 2277.730 2644.690 2278.910 2645.870 ;
        RECT 2279.330 2644.690 2280.510 2645.870 ;
        RECT 2277.730 2643.090 2278.910 2644.270 ;
        RECT 2279.330 2643.090 2280.510 2644.270 ;
        RECT 2277.730 2464.690 2278.910 2465.870 ;
        RECT 2279.330 2464.690 2280.510 2465.870 ;
        RECT 2277.730 2463.090 2278.910 2464.270 ;
        RECT 2279.330 2463.090 2280.510 2464.270 ;
        RECT 2277.730 2284.690 2278.910 2285.870 ;
        RECT 2279.330 2284.690 2280.510 2285.870 ;
        RECT 2277.730 2283.090 2278.910 2284.270 ;
        RECT 2279.330 2283.090 2280.510 2284.270 ;
        RECT 2277.730 2104.690 2278.910 2105.870 ;
        RECT 2279.330 2104.690 2280.510 2105.870 ;
        RECT 2277.730 2103.090 2278.910 2104.270 ;
        RECT 2279.330 2103.090 2280.510 2104.270 ;
        RECT 2277.730 1924.690 2278.910 1925.870 ;
        RECT 2279.330 1924.690 2280.510 1925.870 ;
        RECT 2277.730 1923.090 2278.910 1924.270 ;
        RECT 2279.330 1923.090 2280.510 1924.270 ;
        RECT 2277.730 1744.690 2278.910 1745.870 ;
        RECT 2279.330 1744.690 2280.510 1745.870 ;
        RECT 2277.730 1743.090 2278.910 1744.270 ;
        RECT 2279.330 1743.090 2280.510 1744.270 ;
        RECT 2277.730 1564.690 2278.910 1565.870 ;
        RECT 2279.330 1564.690 2280.510 1565.870 ;
        RECT 2277.730 1563.090 2278.910 1564.270 ;
        RECT 2279.330 1563.090 2280.510 1564.270 ;
        RECT 2277.730 1384.690 2278.910 1385.870 ;
        RECT 2279.330 1384.690 2280.510 1385.870 ;
        RECT 2277.730 1383.090 2278.910 1384.270 ;
        RECT 2279.330 1383.090 2280.510 1384.270 ;
        RECT 2277.730 1204.690 2278.910 1205.870 ;
        RECT 2279.330 1204.690 2280.510 1205.870 ;
        RECT 2277.730 1203.090 2278.910 1204.270 ;
        RECT 2279.330 1203.090 2280.510 1204.270 ;
        RECT 2277.730 1024.690 2278.910 1025.870 ;
        RECT 2279.330 1024.690 2280.510 1025.870 ;
        RECT 2277.730 1023.090 2278.910 1024.270 ;
        RECT 2279.330 1023.090 2280.510 1024.270 ;
        RECT 2277.730 844.690 2278.910 845.870 ;
        RECT 2279.330 844.690 2280.510 845.870 ;
        RECT 2277.730 843.090 2278.910 844.270 ;
        RECT 2279.330 843.090 2280.510 844.270 ;
        RECT 2277.730 664.690 2278.910 665.870 ;
        RECT 2279.330 664.690 2280.510 665.870 ;
        RECT 2277.730 663.090 2278.910 664.270 ;
        RECT 2279.330 663.090 2280.510 664.270 ;
        RECT 2277.730 484.690 2278.910 485.870 ;
        RECT 2279.330 484.690 2280.510 485.870 ;
        RECT 2277.730 483.090 2278.910 484.270 ;
        RECT 2279.330 483.090 2280.510 484.270 ;
        RECT 2277.730 304.690 2278.910 305.870 ;
        RECT 2279.330 304.690 2280.510 305.870 ;
        RECT 2277.730 303.090 2278.910 304.270 ;
        RECT 2279.330 303.090 2280.510 304.270 ;
        RECT 2277.730 124.690 2278.910 125.870 ;
        RECT 2279.330 124.690 2280.510 125.870 ;
        RECT 2277.730 123.090 2278.910 124.270 ;
        RECT 2279.330 123.090 2280.510 124.270 ;
        RECT 2277.730 -17.310 2278.910 -16.130 ;
        RECT 2279.330 -17.310 2280.510 -16.130 ;
        RECT 2277.730 -18.910 2278.910 -17.730 ;
        RECT 2279.330 -18.910 2280.510 -17.730 ;
        RECT 2457.730 3537.410 2458.910 3538.590 ;
        RECT 2459.330 3537.410 2460.510 3538.590 ;
        RECT 2457.730 3535.810 2458.910 3536.990 ;
        RECT 2459.330 3535.810 2460.510 3536.990 ;
        RECT 2457.730 3364.690 2458.910 3365.870 ;
        RECT 2459.330 3364.690 2460.510 3365.870 ;
        RECT 2457.730 3363.090 2458.910 3364.270 ;
        RECT 2459.330 3363.090 2460.510 3364.270 ;
        RECT 2457.730 3184.690 2458.910 3185.870 ;
        RECT 2459.330 3184.690 2460.510 3185.870 ;
        RECT 2457.730 3183.090 2458.910 3184.270 ;
        RECT 2459.330 3183.090 2460.510 3184.270 ;
        RECT 2457.730 3004.690 2458.910 3005.870 ;
        RECT 2459.330 3004.690 2460.510 3005.870 ;
        RECT 2457.730 3003.090 2458.910 3004.270 ;
        RECT 2459.330 3003.090 2460.510 3004.270 ;
        RECT 2457.730 2824.690 2458.910 2825.870 ;
        RECT 2459.330 2824.690 2460.510 2825.870 ;
        RECT 2457.730 2823.090 2458.910 2824.270 ;
        RECT 2459.330 2823.090 2460.510 2824.270 ;
        RECT 2457.730 2644.690 2458.910 2645.870 ;
        RECT 2459.330 2644.690 2460.510 2645.870 ;
        RECT 2457.730 2643.090 2458.910 2644.270 ;
        RECT 2459.330 2643.090 2460.510 2644.270 ;
        RECT 2457.730 2464.690 2458.910 2465.870 ;
        RECT 2459.330 2464.690 2460.510 2465.870 ;
        RECT 2457.730 2463.090 2458.910 2464.270 ;
        RECT 2459.330 2463.090 2460.510 2464.270 ;
        RECT 2457.730 2284.690 2458.910 2285.870 ;
        RECT 2459.330 2284.690 2460.510 2285.870 ;
        RECT 2457.730 2283.090 2458.910 2284.270 ;
        RECT 2459.330 2283.090 2460.510 2284.270 ;
        RECT 2457.730 2104.690 2458.910 2105.870 ;
        RECT 2459.330 2104.690 2460.510 2105.870 ;
        RECT 2457.730 2103.090 2458.910 2104.270 ;
        RECT 2459.330 2103.090 2460.510 2104.270 ;
        RECT 2457.730 1924.690 2458.910 1925.870 ;
        RECT 2459.330 1924.690 2460.510 1925.870 ;
        RECT 2457.730 1923.090 2458.910 1924.270 ;
        RECT 2459.330 1923.090 2460.510 1924.270 ;
        RECT 2457.730 1744.690 2458.910 1745.870 ;
        RECT 2459.330 1744.690 2460.510 1745.870 ;
        RECT 2457.730 1743.090 2458.910 1744.270 ;
        RECT 2459.330 1743.090 2460.510 1744.270 ;
        RECT 2457.730 1564.690 2458.910 1565.870 ;
        RECT 2459.330 1564.690 2460.510 1565.870 ;
        RECT 2457.730 1563.090 2458.910 1564.270 ;
        RECT 2459.330 1563.090 2460.510 1564.270 ;
        RECT 2457.730 1384.690 2458.910 1385.870 ;
        RECT 2459.330 1384.690 2460.510 1385.870 ;
        RECT 2457.730 1383.090 2458.910 1384.270 ;
        RECT 2459.330 1383.090 2460.510 1384.270 ;
        RECT 2457.730 1204.690 2458.910 1205.870 ;
        RECT 2459.330 1204.690 2460.510 1205.870 ;
        RECT 2457.730 1203.090 2458.910 1204.270 ;
        RECT 2459.330 1203.090 2460.510 1204.270 ;
        RECT 2457.730 1024.690 2458.910 1025.870 ;
        RECT 2459.330 1024.690 2460.510 1025.870 ;
        RECT 2457.730 1023.090 2458.910 1024.270 ;
        RECT 2459.330 1023.090 2460.510 1024.270 ;
        RECT 2457.730 844.690 2458.910 845.870 ;
        RECT 2459.330 844.690 2460.510 845.870 ;
        RECT 2457.730 843.090 2458.910 844.270 ;
        RECT 2459.330 843.090 2460.510 844.270 ;
        RECT 2457.730 664.690 2458.910 665.870 ;
        RECT 2459.330 664.690 2460.510 665.870 ;
        RECT 2457.730 663.090 2458.910 664.270 ;
        RECT 2459.330 663.090 2460.510 664.270 ;
        RECT 2457.730 484.690 2458.910 485.870 ;
        RECT 2459.330 484.690 2460.510 485.870 ;
        RECT 2457.730 483.090 2458.910 484.270 ;
        RECT 2459.330 483.090 2460.510 484.270 ;
        RECT 2457.730 304.690 2458.910 305.870 ;
        RECT 2459.330 304.690 2460.510 305.870 ;
        RECT 2457.730 303.090 2458.910 304.270 ;
        RECT 2459.330 303.090 2460.510 304.270 ;
        RECT 2457.730 124.690 2458.910 125.870 ;
        RECT 2459.330 124.690 2460.510 125.870 ;
        RECT 2457.730 123.090 2458.910 124.270 ;
        RECT 2459.330 123.090 2460.510 124.270 ;
        RECT 2457.730 -17.310 2458.910 -16.130 ;
        RECT 2459.330 -17.310 2460.510 -16.130 ;
        RECT 2457.730 -18.910 2458.910 -17.730 ;
        RECT 2459.330 -18.910 2460.510 -17.730 ;
        RECT 2637.730 3537.410 2638.910 3538.590 ;
        RECT 2639.330 3537.410 2640.510 3538.590 ;
        RECT 2637.730 3535.810 2638.910 3536.990 ;
        RECT 2639.330 3535.810 2640.510 3536.990 ;
        RECT 2637.730 3364.690 2638.910 3365.870 ;
        RECT 2639.330 3364.690 2640.510 3365.870 ;
        RECT 2637.730 3363.090 2638.910 3364.270 ;
        RECT 2639.330 3363.090 2640.510 3364.270 ;
        RECT 2637.730 3184.690 2638.910 3185.870 ;
        RECT 2639.330 3184.690 2640.510 3185.870 ;
        RECT 2637.730 3183.090 2638.910 3184.270 ;
        RECT 2639.330 3183.090 2640.510 3184.270 ;
        RECT 2637.730 3004.690 2638.910 3005.870 ;
        RECT 2639.330 3004.690 2640.510 3005.870 ;
        RECT 2637.730 3003.090 2638.910 3004.270 ;
        RECT 2639.330 3003.090 2640.510 3004.270 ;
        RECT 2637.730 2824.690 2638.910 2825.870 ;
        RECT 2639.330 2824.690 2640.510 2825.870 ;
        RECT 2637.730 2823.090 2638.910 2824.270 ;
        RECT 2639.330 2823.090 2640.510 2824.270 ;
        RECT 2637.730 2644.690 2638.910 2645.870 ;
        RECT 2639.330 2644.690 2640.510 2645.870 ;
        RECT 2637.730 2643.090 2638.910 2644.270 ;
        RECT 2639.330 2643.090 2640.510 2644.270 ;
        RECT 2637.730 2464.690 2638.910 2465.870 ;
        RECT 2639.330 2464.690 2640.510 2465.870 ;
        RECT 2637.730 2463.090 2638.910 2464.270 ;
        RECT 2639.330 2463.090 2640.510 2464.270 ;
        RECT 2637.730 2284.690 2638.910 2285.870 ;
        RECT 2639.330 2284.690 2640.510 2285.870 ;
        RECT 2637.730 2283.090 2638.910 2284.270 ;
        RECT 2639.330 2283.090 2640.510 2284.270 ;
        RECT 2637.730 2104.690 2638.910 2105.870 ;
        RECT 2639.330 2104.690 2640.510 2105.870 ;
        RECT 2637.730 2103.090 2638.910 2104.270 ;
        RECT 2639.330 2103.090 2640.510 2104.270 ;
        RECT 2637.730 1924.690 2638.910 1925.870 ;
        RECT 2639.330 1924.690 2640.510 1925.870 ;
        RECT 2637.730 1923.090 2638.910 1924.270 ;
        RECT 2639.330 1923.090 2640.510 1924.270 ;
        RECT 2637.730 1744.690 2638.910 1745.870 ;
        RECT 2639.330 1744.690 2640.510 1745.870 ;
        RECT 2637.730 1743.090 2638.910 1744.270 ;
        RECT 2639.330 1743.090 2640.510 1744.270 ;
        RECT 2637.730 1564.690 2638.910 1565.870 ;
        RECT 2639.330 1564.690 2640.510 1565.870 ;
        RECT 2637.730 1563.090 2638.910 1564.270 ;
        RECT 2639.330 1563.090 2640.510 1564.270 ;
        RECT 2637.730 1384.690 2638.910 1385.870 ;
        RECT 2639.330 1384.690 2640.510 1385.870 ;
        RECT 2637.730 1383.090 2638.910 1384.270 ;
        RECT 2639.330 1383.090 2640.510 1384.270 ;
        RECT 2637.730 1204.690 2638.910 1205.870 ;
        RECT 2639.330 1204.690 2640.510 1205.870 ;
        RECT 2637.730 1203.090 2638.910 1204.270 ;
        RECT 2639.330 1203.090 2640.510 1204.270 ;
        RECT 2637.730 1024.690 2638.910 1025.870 ;
        RECT 2639.330 1024.690 2640.510 1025.870 ;
        RECT 2637.730 1023.090 2638.910 1024.270 ;
        RECT 2639.330 1023.090 2640.510 1024.270 ;
        RECT 2637.730 844.690 2638.910 845.870 ;
        RECT 2639.330 844.690 2640.510 845.870 ;
        RECT 2637.730 843.090 2638.910 844.270 ;
        RECT 2639.330 843.090 2640.510 844.270 ;
        RECT 2637.730 664.690 2638.910 665.870 ;
        RECT 2639.330 664.690 2640.510 665.870 ;
        RECT 2637.730 663.090 2638.910 664.270 ;
        RECT 2639.330 663.090 2640.510 664.270 ;
        RECT 2637.730 484.690 2638.910 485.870 ;
        RECT 2639.330 484.690 2640.510 485.870 ;
        RECT 2637.730 483.090 2638.910 484.270 ;
        RECT 2639.330 483.090 2640.510 484.270 ;
        RECT 2637.730 304.690 2638.910 305.870 ;
        RECT 2639.330 304.690 2640.510 305.870 ;
        RECT 2637.730 303.090 2638.910 304.270 ;
        RECT 2639.330 303.090 2640.510 304.270 ;
        RECT 2637.730 124.690 2638.910 125.870 ;
        RECT 2639.330 124.690 2640.510 125.870 ;
        RECT 2637.730 123.090 2638.910 124.270 ;
        RECT 2639.330 123.090 2640.510 124.270 ;
        RECT 2637.730 -17.310 2638.910 -16.130 ;
        RECT 2639.330 -17.310 2640.510 -16.130 ;
        RECT 2637.730 -18.910 2638.910 -17.730 ;
        RECT 2639.330 -18.910 2640.510 -17.730 ;
        RECT 2817.730 3537.410 2818.910 3538.590 ;
        RECT 2819.330 3537.410 2820.510 3538.590 ;
        RECT 2817.730 3535.810 2818.910 3536.990 ;
        RECT 2819.330 3535.810 2820.510 3536.990 ;
        RECT 2817.730 3364.690 2818.910 3365.870 ;
        RECT 2819.330 3364.690 2820.510 3365.870 ;
        RECT 2817.730 3363.090 2818.910 3364.270 ;
        RECT 2819.330 3363.090 2820.510 3364.270 ;
        RECT 2817.730 3184.690 2818.910 3185.870 ;
        RECT 2819.330 3184.690 2820.510 3185.870 ;
        RECT 2817.730 3183.090 2818.910 3184.270 ;
        RECT 2819.330 3183.090 2820.510 3184.270 ;
        RECT 2817.730 3004.690 2818.910 3005.870 ;
        RECT 2819.330 3004.690 2820.510 3005.870 ;
        RECT 2817.730 3003.090 2818.910 3004.270 ;
        RECT 2819.330 3003.090 2820.510 3004.270 ;
        RECT 2817.730 2824.690 2818.910 2825.870 ;
        RECT 2819.330 2824.690 2820.510 2825.870 ;
        RECT 2817.730 2823.090 2818.910 2824.270 ;
        RECT 2819.330 2823.090 2820.510 2824.270 ;
        RECT 2817.730 2644.690 2818.910 2645.870 ;
        RECT 2819.330 2644.690 2820.510 2645.870 ;
        RECT 2817.730 2643.090 2818.910 2644.270 ;
        RECT 2819.330 2643.090 2820.510 2644.270 ;
        RECT 2817.730 2464.690 2818.910 2465.870 ;
        RECT 2819.330 2464.690 2820.510 2465.870 ;
        RECT 2817.730 2463.090 2818.910 2464.270 ;
        RECT 2819.330 2463.090 2820.510 2464.270 ;
        RECT 2817.730 2284.690 2818.910 2285.870 ;
        RECT 2819.330 2284.690 2820.510 2285.870 ;
        RECT 2817.730 2283.090 2818.910 2284.270 ;
        RECT 2819.330 2283.090 2820.510 2284.270 ;
        RECT 2817.730 2104.690 2818.910 2105.870 ;
        RECT 2819.330 2104.690 2820.510 2105.870 ;
        RECT 2817.730 2103.090 2818.910 2104.270 ;
        RECT 2819.330 2103.090 2820.510 2104.270 ;
        RECT 2817.730 1924.690 2818.910 1925.870 ;
        RECT 2819.330 1924.690 2820.510 1925.870 ;
        RECT 2817.730 1923.090 2818.910 1924.270 ;
        RECT 2819.330 1923.090 2820.510 1924.270 ;
        RECT 2817.730 1744.690 2818.910 1745.870 ;
        RECT 2819.330 1744.690 2820.510 1745.870 ;
        RECT 2817.730 1743.090 2818.910 1744.270 ;
        RECT 2819.330 1743.090 2820.510 1744.270 ;
        RECT 2817.730 1564.690 2818.910 1565.870 ;
        RECT 2819.330 1564.690 2820.510 1565.870 ;
        RECT 2817.730 1563.090 2818.910 1564.270 ;
        RECT 2819.330 1563.090 2820.510 1564.270 ;
        RECT 2817.730 1384.690 2818.910 1385.870 ;
        RECT 2819.330 1384.690 2820.510 1385.870 ;
        RECT 2817.730 1383.090 2818.910 1384.270 ;
        RECT 2819.330 1383.090 2820.510 1384.270 ;
        RECT 2817.730 1204.690 2818.910 1205.870 ;
        RECT 2819.330 1204.690 2820.510 1205.870 ;
        RECT 2817.730 1203.090 2818.910 1204.270 ;
        RECT 2819.330 1203.090 2820.510 1204.270 ;
        RECT 2817.730 1024.690 2818.910 1025.870 ;
        RECT 2819.330 1024.690 2820.510 1025.870 ;
        RECT 2817.730 1023.090 2818.910 1024.270 ;
        RECT 2819.330 1023.090 2820.510 1024.270 ;
        RECT 2817.730 844.690 2818.910 845.870 ;
        RECT 2819.330 844.690 2820.510 845.870 ;
        RECT 2817.730 843.090 2818.910 844.270 ;
        RECT 2819.330 843.090 2820.510 844.270 ;
        RECT 2817.730 664.690 2818.910 665.870 ;
        RECT 2819.330 664.690 2820.510 665.870 ;
        RECT 2817.730 663.090 2818.910 664.270 ;
        RECT 2819.330 663.090 2820.510 664.270 ;
        RECT 2817.730 484.690 2818.910 485.870 ;
        RECT 2819.330 484.690 2820.510 485.870 ;
        RECT 2817.730 483.090 2818.910 484.270 ;
        RECT 2819.330 483.090 2820.510 484.270 ;
        RECT 2817.730 304.690 2818.910 305.870 ;
        RECT 2819.330 304.690 2820.510 305.870 ;
        RECT 2817.730 303.090 2818.910 304.270 ;
        RECT 2819.330 303.090 2820.510 304.270 ;
        RECT 2817.730 124.690 2818.910 125.870 ;
        RECT 2819.330 124.690 2820.510 125.870 ;
        RECT 2817.730 123.090 2818.910 124.270 ;
        RECT 2819.330 123.090 2820.510 124.270 ;
        RECT 2817.730 -17.310 2818.910 -16.130 ;
        RECT 2819.330 -17.310 2820.510 -16.130 ;
        RECT 2817.730 -18.910 2818.910 -17.730 ;
        RECT 2819.330 -18.910 2820.510 -17.730 ;
        RECT 2941.110 3537.410 2942.290 3538.590 ;
        RECT 2942.710 3537.410 2943.890 3538.590 ;
        RECT 2941.110 3535.810 2942.290 3536.990 ;
        RECT 2942.710 3535.810 2943.890 3536.990 ;
        RECT 2941.110 3364.690 2942.290 3365.870 ;
        RECT 2942.710 3364.690 2943.890 3365.870 ;
        RECT 2941.110 3363.090 2942.290 3364.270 ;
        RECT 2942.710 3363.090 2943.890 3364.270 ;
        RECT 2941.110 3184.690 2942.290 3185.870 ;
        RECT 2942.710 3184.690 2943.890 3185.870 ;
        RECT 2941.110 3183.090 2942.290 3184.270 ;
        RECT 2942.710 3183.090 2943.890 3184.270 ;
        RECT 2941.110 3004.690 2942.290 3005.870 ;
        RECT 2942.710 3004.690 2943.890 3005.870 ;
        RECT 2941.110 3003.090 2942.290 3004.270 ;
        RECT 2942.710 3003.090 2943.890 3004.270 ;
        RECT 2941.110 2824.690 2942.290 2825.870 ;
        RECT 2942.710 2824.690 2943.890 2825.870 ;
        RECT 2941.110 2823.090 2942.290 2824.270 ;
        RECT 2942.710 2823.090 2943.890 2824.270 ;
        RECT 2941.110 2644.690 2942.290 2645.870 ;
        RECT 2942.710 2644.690 2943.890 2645.870 ;
        RECT 2941.110 2643.090 2942.290 2644.270 ;
        RECT 2942.710 2643.090 2943.890 2644.270 ;
        RECT 2941.110 2464.690 2942.290 2465.870 ;
        RECT 2942.710 2464.690 2943.890 2465.870 ;
        RECT 2941.110 2463.090 2942.290 2464.270 ;
        RECT 2942.710 2463.090 2943.890 2464.270 ;
        RECT 2941.110 2284.690 2942.290 2285.870 ;
        RECT 2942.710 2284.690 2943.890 2285.870 ;
        RECT 2941.110 2283.090 2942.290 2284.270 ;
        RECT 2942.710 2283.090 2943.890 2284.270 ;
        RECT 2941.110 2104.690 2942.290 2105.870 ;
        RECT 2942.710 2104.690 2943.890 2105.870 ;
        RECT 2941.110 2103.090 2942.290 2104.270 ;
        RECT 2942.710 2103.090 2943.890 2104.270 ;
        RECT 2941.110 1924.690 2942.290 1925.870 ;
        RECT 2942.710 1924.690 2943.890 1925.870 ;
        RECT 2941.110 1923.090 2942.290 1924.270 ;
        RECT 2942.710 1923.090 2943.890 1924.270 ;
        RECT 2941.110 1744.690 2942.290 1745.870 ;
        RECT 2942.710 1744.690 2943.890 1745.870 ;
        RECT 2941.110 1743.090 2942.290 1744.270 ;
        RECT 2942.710 1743.090 2943.890 1744.270 ;
        RECT 2941.110 1564.690 2942.290 1565.870 ;
        RECT 2942.710 1564.690 2943.890 1565.870 ;
        RECT 2941.110 1563.090 2942.290 1564.270 ;
        RECT 2942.710 1563.090 2943.890 1564.270 ;
        RECT 2941.110 1384.690 2942.290 1385.870 ;
        RECT 2942.710 1384.690 2943.890 1385.870 ;
        RECT 2941.110 1383.090 2942.290 1384.270 ;
        RECT 2942.710 1383.090 2943.890 1384.270 ;
        RECT 2941.110 1204.690 2942.290 1205.870 ;
        RECT 2942.710 1204.690 2943.890 1205.870 ;
        RECT 2941.110 1203.090 2942.290 1204.270 ;
        RECT 2942.710 1203.090 2943.890 1204.270 ;
        RECT 2941.110 1024.690 2942.290 1025.870 ;
        RECT 2942.710 1024.690 2943.890 1025.870 ;
        RECT 2941.110 1023.090 2942.290 1024.270 ;
        RECT 2942.710 1023.090 2943.890 1024.270 ;
        RECT 2941.110 844.690 2942.290 845.870 ;
        RECT 2942.710 844.690 2943.890 845.870 ;
        RECT 2941.110 843.090 2942.290 844.270 ;
        RECT 2942.710 843.090 2943.890 844.270 ;
        RECT 2941.110 664.690 2942.290 665.870 ;
        RECT 2942.710 664.690 2943.890 665.870 ;
        RECT 2941.110 663.090 2942.290 664.270 ;
        RECT 2942.710 663.090 2943.890 664.270 ;
        RECT 2941.110 484.690 2942.290 485.870 ;
        RECT 2942.710 484.690 2943.890 485.870 ;
        RECT 2941.110 483.090 2942.290 484.270 ;
        RECT 2942.710 483.090 2943.890 484.270 ;
        RECT 2941.110 304.690 2942.290 305.870 ;
        RECT 2942.710 304.690 2943.890 305.870 ;
        RECT 2941.110 303.090 2942.290 304.270 ;
        RECT 2942.710 303.090 2943.890 304.270 ;
        RECT 2941.110 124.690 2942.290 125.870 ;
        RECT 2942.710 124.690 2943.890 125.870 ;
        RECT 2941.110 123.090 2942.290 124.270 ;
        RECT 2942.710 123.090 2943.890 124.270 ;
        RECT 2941.110 -17.310 2942.290 -16.130 ;
        RECT 2942.710 -17.310 2943.890 -16.130 ;
        RECT 2941.110 -18.910 2942.290 -17.730 ;
        RECT 2942.710 -18.910 2943.890 -17.730 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
        RECT -24.430 842.930 2944.050 846.030 ;
        RECT -24.430 662.930 2944.050 666.030 ;
        RECT -24.430 482.930 2944.050 486.030 ;
        RECT -24.430 302.930 2944.050 306.030 ;
        RECT -24.430 122.930 2944.050 126.030 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.930 401.610 202.210 404.000 ;
        RECT 201.180 401.470 202.210 401.610 ;
        RECT 201.180 386.650 201.320 401.470 ;
        RECT 201.930 400.000 202.210 401.470 ;
        RECT 200.720 386.510 201.320 386.650 ;
        RECT 200.720 16.845 200.860 386.510 ;
        RECT 8.370 16.475 8.650 16.845 ;
        RECT 200.650 16.475 200.930 16.845 ;
        RECT 8.440 2.400 8.580 16.475 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 8.370 16.520 8.650 16.800 ;
        RECT 200.650 16.520 200.930 16.800 ;
      LAYER met3 ;
        RECT 8.345 16.810 8.675 16.825 ;
        RECT 200.625 16.810 200.955 16.825 ;
        RECT 8.345 16.510 200.955 16.810 ;
        RECT 8.345 16.495 8.675 16.510 ;
        RECT 200.625 16.495 200.955 16.510 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 201.090 17.580 201.410 17.640 ;
        RECT 14.330 17.440 201.410 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 201.090 17.380 201.410 17.440 ;
      LAYER via ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 201.120 17.380 201.380 17.640 ;
      LAYER met2 ;
        RECT 203.770 400.250 204.050 404.000 ;
        RECT 202.560 400.110 204.050 400.250 ;
        RECT 202.560 385.290 202.700 400.110 ;
        RECT 203.770 400.000 204.050 400.110 ;
        RECT 201.180 385.150 202.700 385.290 ;
        RECT 201.180 17.670 201.320 385.150 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 201.120 17.350 201.380 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 207.530 376.280 207.850 376.340 ;
        RECT 209.830 376.280 210.150 376.340 ;
        RECT 207.530 376.140 210.150 376.280 ;
        RECT 207.530 376.080 207.850 376.140 ;
        RECT 209.830 376.080 210.150 376.140 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 207.530 17.920 207.850 17.980 ;
        RECT 38.250 17.780 207.850 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 207.530 17.720 207.850 17.780 ;
      LAYER via ;
        RECT 207.560 376.080 207.820 376.340 ;
        RECT 209.860 376.080 210.120 376.340 ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 207.560 17.720 207.820 17.980 ;
      LAYER met2 ;
        RECT 211.130 400.250 211.410 404.000 ;
        RECT 209.920 400.110 211.410 400.250 ;
        RECT 209.920 376.370 210.060 400.110 ;
        RECT 211.130 400.000 211.410 400.110 ;
        RECT 207.560 376.050 207.820 376.370 ;
        RECT 209.860 376.050 210.120 376.370 ;
        RECT 207.620 18.010 207.760 376.050 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 207.560 17.690 207.820 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 239.270 17.920 239.590 17.980 ;
        RECT 269.630 17.920 269.950 17.980 ;
        RECT 239.270 17.780 269.950 17.920 ;
        RECT 239.270 17.720 239.590 17.780 ;
        RECT 269.630 17.720 269.950 17.780 ;
      LAYER via ;
        RECT 239.300 17.720 239.560 17.980 ;
        RECT 269.660 17.720 269.920 17.980 ;
      LAYER met2 ;
        RECT 271.850 400.250 272.130 404.000 ;
        RECT 270.640 400.110 272.130 400.250 ;
        RECT 270.640 324.370 270.780 400.110 ;
        RECT 271.850 400.000 272.130 400.110 ;
        RECT 269.720 324.230 270.780 324.370 ;
        RECT 269.720 18.010 269.860 324.230 ;
        RECT 239.300 17.690 239.560 18.010 ;
        RECT 269.660 17.690 269.920 18.010 ;
        RECT 239.360 2.400 239.500 17.690 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 255.370 391.920 255.690 391.980 ;
        RECT 276.990 391.920 277.310 391.980 ;
        RECT 255.370 391.780 277.310 391.920 ;
        RECT 255.370 391.720 255.690 391.780 ;
        RECT 276.990 391.720 277.310 391.780 ;
      LAYER via ;
        RECT 255.400 391.720 255.660 391.980 ;
        RECT 277.020 391.720 277.280 391.980 ;
      LAYER met2 ;
        RECT 276.910 400.180 277.190 404.000 ;
        RECT 276.910 400.000 277.220 400.180 ;
        RECT 277.080 392.010 277.220 400.000 ;
        RECT 255.400 391.690 255.660 392.010 ;
        RECT 277.020 391.690 277.280 392.010 ;
        RECT 255.460 1.770 255.600 391.690 ;
        RECT 256.630 1.770 257.190 2.400 ;
        RECT 255.460 1.630 257.190 1.770 ;
        RECT 256.630 -4.800 257.190 1.630 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 271.010 393.280 271.330 393.340 ;
        RECT 282.510 393.280 282.830 393.340 ;
        RECT 271.010 393.140 282.830 393.280 ;
        RECT 271.010 393.080 271.330 393.140 ;
        RECT 282.510 393.080 282.830 393.140 ;
      LAYER via ;
        RECT 271.040 393.080 271.300 393.340 ;
        RECT 282.540 393.080 282.800 393.340 ;
      LAYER met2 ;
        RECT 282.430 400.180 282.710 404.000 ;
        RECT 282.430 400.000 282.740 400.180 ;
        RECT 282.600 393.370 282.740 400.000 ;
        RECT 271.040 393.050 271.300 393.370 ;
        RECT 282.540 393.050 282.800 393.370 ;
        RECT 271.100 82.870 271.240 393.050 ;
        RECT 271.100 82.730 274.920 82.870 ;
        RECT 274.780 2.400 274.920 82.730 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.950 400.250 288.230 404.000 ;
        RECT 287.950 400.110 289.640 400.250 ;
        RECT 287.950 400.000 288.230 400.110 ;
        RECT 289.500 386.470 289.640 400.110 ;
        RECT 289.500 386.330 290.100 386.470 ;
        RECT 289.960 16.730 290.100 386.330 ;
        RECT 289.960 16.590 292.400 16.730 ;
        RECT 292.260 2.400 292.400 16.590 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.790 386.140 291.110 386.200 ;
        RECT 292.170 386.140 292.490 386.200 ;
        RECT 290.790 386.000 292.490 386.140 ;
        RECT 290.790 385.940 291.110 386.000 ;
        RECT 292.170 385.940 292.490 386.000 ;
        RECT 290.790 17.240 291.110 17.300 ;
        RECT 310.110 17.240 310.430 17.300 ;
        RECT 290.790 17.100 310.430 17.240 ;
        RECT 290.790 17.040 291.110 17.100 ;
        RECT 310.110 17.040 310.430 17.100 ;
      LAYER via ;
        RECT 290.820 385.940 291.080 386.200 ;
        RECT 292.200 385.940 292.460 386.200 ;
        RECT 290.820 17.040 291.080 17.300 ;
        RECT 310.140 17.040 310.400 17.300 ;
      LAYER met2 ;
        RECT 293.010 400.250 293.290 404.000 ;
        RECT 292.260 400.110 293.290 400.250 ;
        RECT 292.260 386.230 292.400 400.110 ;
        RECT 293.010 400.000 293.290 400.110 ;
        RECT 290.820 385.910 291.080 386.230 ;
        RECT 292.200 385.910 292.460 386.230 ;
        RECT 290.880 17.330 291.020 385.910 ;
        RECT 290.820 17.010 291.080 17.330 ;
        RECT 310.140 17.010 310.400 17.330 ;
        RECT 310.200 2.400 310.340 17.010 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 298.610 387.500 298.930 387.560 ;
        RECT 306.890 387.500 307.210 387.560 ;
        RECT 298.610 387.360 307.210 387.500 ;
        RECT 298.610 387.300 298.930 387.360 ;
        RECT 306.890 387.300 307.210 387.360 ;
        RECT 306.890 19.960 307.210 20.020 ;
        RECT 327.590 19.960 327.910 20.020 ;
        RECT 306.890 19.820 327.910 19.960 ;
        RECT 306.890 19.760 307.210 19.820 ;
        RECT 327.590 19.760 327.910 19.820 ;
      LAYER via ;
        RECT 298.640 387.300 298.900 387.560 ;
        RECT 306.920 387.300 307.180 387.560 ;
        RECT 306.920 19.760 307.180 20.020 ;
        RECT 327.620 19.760 327.880 20.020 ;
      LAYER met2 ;
        RECT 298.530 400.180 298.810 404.000 ;
        RECT 298.530 400.000 298.840 400.180 ;
        RECT 298.700 387.590 298.840 400.000 ;
        RECT 298.640 387.270 298.900 387.590 ;
        RECT 306.920 387.270 307.180 387.590 ;
        RECT 306.980 20.050 307.120 387.270 ;
        RECT 306.920 19.730 307.180 20.050 ;
        RECT 327.620 19.730 327.880 20.050 ;
        RECT 327.680 2.400 327.820 19.730 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.590 18.940 304.910 19.000 ;
        RECT 345.530 18.940 345.850 19.000 ;
        RECT 304.590 18.800 345.850 18.940 ;
        RECT 304.590 18.740 304.910 18.800 ;
        RECT 345.530 18.740 345.850 18.800 ;
      LAYER via ;
        RECT 304.620 18.740 304.880 19.000 ;
        RECT 345.560 18.740 345.820 19.000 ;
      LAYER met2 ;
        RECT 304.050 400.250 304.330 404.000 ;
        RECT 304.050 400.110 304.820 400.250 ;
        RECT 304.050 400.000 304.330 400.110 ;
        RECT 304.680 19.030 304.820 400.110 ;
        RECT 304.620 18.710 304.880 19.030 ;
        RECT 345.560 18.710 345.820 19.030 ;
        RECT 345.620 2.400 345.760 18.710 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.130 375.940 304.450 376.000 ;
        RECT 307.810 375.940 308.130 376.000 ;
        RECT 304.130 375.800 308.130 375.940 ;
        RECT 304.130 375.740 304.450 375.800 ;
        RECT 307.810 375.740 308.130 375.800 ;
        RECT 304.130 18.600 304.450 18.660 ;
        RECT 304.130 18.460 320.000 18.600 ;
        RECT 304.130 18.400 304.450 18.460 ;
        RECT 319.860 18.260 320.000 18.460 ;
        RECT 363.010 18.260 363.330 18.320 ;
        RECT 319.860 18.120 363.330 18.260 ;
        RECT 363.010 18.060 363.330 18.120 ;
      LAYER via ;
        RECT 304.160 375.740 304.420 376.000 ;
        RECT 307.840 375.740 308.100 376.000 ;
        RECT 304.160 18.400 304.420 18.660 ;
        RECT 363.040 18.060 363.300 18.320 ;
      LAYER met2 ;
        RECT 309.110 400.250 309.390 404.000 ;
        RECT 307.900 400.110 309.390 400.250 ;
        RECT 307.900 376.030 308.040 400.110 ;
        RECT 309.110 400.000 309.390 400.110 ;
        RECT 304.160 375.710 304.420 376.030 ;
        RECT 307.840 375.710 308.100 376.030 ;
        RECT 304.220 18.690 304.360 375.710 ;
        RECT 304.160 18.370 304.420 18.690 ;
        RECT 363.040 18.030 363.300 18.350 ;
        RECT 363.100 2.400 363.240 18.030 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 314.710 392.600 315.030 392.660 ;
        RECT 379.570 392.600 379.890 392.660 ;
        RECT 314.710 392.460 379.890 392.600 ;
        RECT 314.710 392.400 315.030 392.460 ;
        RECT 379.570 392.400 379.890 392.460 ;
      LAYER via ;
        RECT 314.740 392.400 315.000 392.660 ;
        RECT 379.600 392.400 379.860 392.660 ;
      LAYER met2 ;
        RECT 314.630 400.180 314.910 404.000 ;
        RECT 314.630 400.000 314.940 400.180 ;
        RECT 314.800 392.690 314.940 400.000 ;
        RECT 314.740 392.370 315.000 392.690 ;
        RECT 379.600 392.370 379.860 392.690 ;
        RECT 379.660 1.770 379.800 392.370 ;
        RECT 380.830 1.770 381.390 2.400 ;
        RECT 379.660 1.630 381.390 1.770 ;
        RECT 380.830 -4.800 381.390 1.630 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 319.310 25.400 319.630 25.460 ;
        RECT 398.430 25.400 398.750 25.460 ;
        RECT 319.310 25.260 398.750 25.400 ;
        RECT 319.310 25.200 319.630 25.260 ;
        RECT 398.430 25.200 398.750 25.260 ;
      LAYER via ;
        RECT 319.340 25.200 319.600 25.460 ;
        RECT 398.460 25.200 398.720 25.460 ;
      LAYER met2 ;
        RECT 320.150 400.250 320.430 404.000 ;
        RECT 319.400 400.110 320.430 400.250 ;
        RECT 319.400 25.490 319.540 400.110 ;
        RECT 320.150 400.000 320.430 400.110 ;
        RECT 319.340 25.170 319.600 25.490 ;
        RECT 398.460 25.170 398.720 25.490 ;
        RECT 398.520 2.400 398.660 25.170 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.890 314.060 215.210 314.120 ;
        RECT 215.810 314.060 216.130 314.120 ;
        RECT 214.890 313.920 216.130 314.060 ;
        RECT 214.890 313.860 215.210 313.920 ;
        RECT 215.810 313.860 216.130 313.920 ;
        RECT 61.710 19.280 62.030 19.340 ;
        RECT 61.710 19.140 197.180 19.280 ;
        RECT 61.710 19.080 62.030 19.140 ;
        RECT 197.040 18.940 197.180 19.140 ;
        RECT 214.890 18.940 215.210 19.000 ;
        RECT 197.040 18.800 215.210 18.940 ;
        RECT 214.890 18.740 215.210 18.800 ;
      LAYER via ;
        RECT 214.920 313.860 215.180 314.120 ;
        RECT 215.840 313.860 216.100 314.120 ;
        RECT 61.740 19.080 62.000 19.340 ;
        RECT 214.920 18.740 215.180 19.000 ;
      LAYER met2 ;
        RECT 218.030 400.250 218.310 404.000 ;
        RECT 216.820 400.110 218.310 400.250 ;
        RECT 216.820 351.970 216.960 400.110 ;
        RECT 218.030 400.000 218.310 400.110 ;
        RECT 215.900 351.830 216.960 351.970 ;
        RECT 215.900 314.150 216.040 351.830 ;
        RECT 214.920 313.830 215.180 314.150 ;
        RECT 215.840 313.830 216.100 314.150 ;
        RECT 61.740 19.050 62.000 19.370 ;
        RECT 61.800 2.400 61.940 19.050 ;
        RECT 214.980 19.030 215.120 313.830 ;
        RECT 214.920 18.710 215.180 19.030 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 325.290 25.060 325.610 25.120 ;
        RECT 416.370 25.060 416.690 25.120 ;
        RECT 325.290 24.920 416.690 25.060 ;
        RECT 325.290 24.860 325.610 24.920 ;
        RECT 416.370 24.860 416.690 24.920 ;
      LAYER via ;
        RECT 325.320 24.860 325.580 25.120 ;
        RECT 416.400 24.860 416.660 25.120 ;
      LAYER met2 ;
        RECT 325.210 400.250 325.490 404.000 ;
        RECT 324.460 400.110 325.490 400.250 ;
        RECT 324.460 386.650 324.600 400.110 ;
        RECT 325.210 400.000 325.490 400.110 ;
        RECT 324.460 386.585 325.520 386.650 ;
        RECT 324.460 386.510 325.590 386.585 ;
        RECT 325.310 386.215 325.590 386.510 ;
        RECT 326.230 385.035 326.510 385.405 ;
        RECT 326.300 338.170 326.440 385.035 ;
        RECT 325.380 338.030 326.440 338.170 ;
        RECT 325.380 25.150 325.520 338.030 ;
        RECT 325.320 24.830 325.580 25.150 ;
        RECT 416.400 24.830 416.660 25.150 ;
        RECT 416.460 2.400 416.600 24.830 ;
        RECT 416.250 -4.800 416.810 2.400 ;
      LAYER via2 ;
        RECT 325.310 386.260 325.590 386.540 ;
        RECT 326.230 385.080 326.510 385.360 ;
      LAYER met3 ;
        RECT 325.285 386.550 325.615 386.565 ;
        RECT 325.070 386.235 325.615 386.550 ;
        RECT 325.070 385.370 325.370 386.235 ;
        RECT 326.205 385.370 326.535 385.385 ;
        RECT 325.070 385.070 326.535 385.370 ;
        RECT 326.205 385.055 326.535 385.070 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 325.750 24.720 326.070 24.780 ;
        RECT 434.310 24.720 434.630 24.780 ;
        RECT 325.750 24.580 434.630 24.720 ;
        RECT 325.750 24.520 326.070 24.580 ;
        RECT 434.310 24.520 434.630 24.580 ;
      LAYER via ;
        RECT 325.780 24.520 326.040 24.780 ;
        RECT 434.340 24.520 434.600 24.780 ;
      LAYER met2 ;
        RECT 330.730 400.250 331.010 404.000 ;
        RECT 329.520 400.110 331.010 400.250 ;
        RECT 329.520 324.370 329.660 400.110 ;
        RECT 330.730 400.000 331.010 400.110 ;
        RECT 325.840 324.230 329.660 324.370 ;
        RECT 325.840 24.810 325.980 324.230 ;
        RECT 325.780 24.490 326.040 24.810 ;
        RECT 434.340 24.490 434.600 24.810 ;
        RECT 434.400 2.400 434.540 24.490 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 336.330 392.940 336.650 393.000 ;
        RECT 445.810 392.940 446.130 393.000 ;
        RECT 336.330 392.800 446.130 392.940 ;
        RECT 336.330 392.740 336.650 392.800 ;
        RECT 445.810 392.740 446.130 392.800 ;
        RECT 444.890 17.580 445.210 17.640 ;
        RECT 451.790 17.580 452.110 17.640 ;
        RECT 444.890 17.440 452.110 17.580 ;
        RECT 444.890 17.380 445.210 17.440 ;
        RECT 451.790 17.380 452.110 17.440 ;
      LAYER via ;
        RECT 336.360 392.740 336.620 393.000 ;
        RECT 445.840 392.740 446.100 393.000 ;
        RECT 444.920 17.380 445.180 17.640 ;
        RECT 451.820 17.380 452.080 17.640 ;
      LAYER met2 ;
        RECT 336.250 400.180 336.530 404.000 ;
        RECT 336.250 400.000 336.560 400.180 ;
        RECT 336.420 393.030 336.560 400.000 ;
        RECT 336.360 392.710 336.620 393.030 ;
        RECT 445.840 392.710 446.100 393.030 ;
        RECT 445.900 324.370 446.040 392.710 ;
        RECT 444.980 324.230 446.040 324.370 ;
        RECT 444.980 17.670 445.120 324.230 ;
        RECT 444.920 17.350 445.180 17.670 ;
        RECT 451.820 17.350 452.080 17.670 ;
        RECT 451.880 2.400 452.020 17.350 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 376.350 391.580 376.670 391.640 ;
        RECT 465.590 391.580 465.910 391.640 ;
        RECT 376.350 391.440 465.910 391.580 ;
        RECT 376.350 391.380 376.670 391.440 ;
        RECT 465.590 391.380 465.910 391.440 ;
        RECT 341.390 389.880 341.710 389.940 ;
        RECT 376.350 389.880 376.670 389.940 ;
        RECT 341.390 389.740 376.670 389.880 ;
        RECT 341.390 389.680 341.710 389.740 ;
        RECT 376.350 389.680 376.670 389.740 ;
        RECT 465.590 20.640 465.910 20.700 ;
        RECT 469.730 20.640 470.050 20.700 ;
        RECT 465.590 20.500 470.050 20.640 ;
        RECT 465.590 20.440 465.910 20.500 ;
        RECT 469.730 20.440 470.050 20.500 ;
      LAYER via ;
        RECT 376.380 391.380 376.640 391.640 ;
        RECT 465.620 391.380 465.880 391.640 ;
        RECT 341.420 389.680 341.680 389.940 ;
        RECT 376.380 389.680 376.640 389.940 ;
        RECT 465.620 20.440 465.880 20.700 ;
        RECT 469.760 20.440 470.020 20.700 ;
      LAYER met2 ;
        RECT 341.310 400.180 341.590 404.000 ;
        RECT 341.310 400.000 341.620 400.180 ;
        RECT 341.480 389.970 341.620 400.000 ;
        RECT 376.380 391.350 376.640 391.670 ;
        RECT 465.620 391.350 465.880 391.670 ;
        RECT 376.440 389.970 376.580 391.350 ;
        RECT 341.420 389.650 341.680 389.970 ;
        RECT 376.380 389.650 376.640 389.970 ;
        RECT 465.680 20.730 465.820 391.350 ;
        RECT 465.620 20.410 465.880 20.730 ;
        RECT 469.760 20.410 470.020 20.730 ;
        RECT 469.820 2.400 469.960 20.410 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 24.040 345.390 24.100 ;
        RECT 487.210 24.040 487.530 24.100 ;
        RECT 345.070 23.900 487.530 24.040 ;
        RECT 345.070 23.840 345.390 23.900 ;
        RECT 487.210 23.840 487.530 23.900 ;
      LAYER via ;
        RECT 345.100 23.840 345.360 24.100 ;
        RECT 487.240 23.840 487.500 24.100 ;
      LAYER met2 ;
        RECT 346.830 400.250 347.110 404.000 ;
        RECT 345.620 400.110 347.110 400.250 ;
        RECT 345.620 324.370 345.760 400.110 ;
        RECT 346.830 400.000 347.110 400.110 ;
        RECT 345.160 324.230 345.760 324.370 ;
        RECT 345.160 24.130 345.300 324.230 ;
        RECT 345.100 23.810 345.360 24.130 ;
        RECT 487.240 23.810 487.500 24.130 ;
        RECT 487.300 2.400 487.440 23.810 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.970 393.280 352.290 393.340 ;
        RECT 353.350 393.280 353.670 393.340 ;
        RECT 351.970 393.140 353.670 393.280 ;
        RECT 351.970 393.080 352.290 393.140 ;
        RECT 353.350 393.080 353.670 393.140 ;
        RECT 472.030 391.920 472.350 391.980 ;
        RECT 375.980 391.780 472.350 391.920 ;
        RECT 353.350 391.580 353.670 391.640 ;
        RECT 375.980 391.580 376.120 391.780 ;
        RECT 472.030 391.720 472.350 391.780 ;
        RECT 353.350 391.440 376.120 391.580 ;
        RECT 353.350 391.380 353.670 391.440 ;
        RECT 472.490 15.200 472.810 15.260 ;
        RECT 505.150 15.200 505.470 15.260 ;
        RECT 472.490 15.060 505.470 15.200 ;
        RECT 472.490 15.000 472.810 15.060 ;
        RECT 505.150 15.000 505.470 15.060 ;
      LAYER via ;
        RECT 352.000 393.080 352.260 393.340 ;
        RECT 353.380 393.080 353.640 393.340 ;
        RECT 353.380 391.380 353.640 391.640 ;
        RECT 472.060 391.720 472.320 391.980 ;
        RECT 472.520 15.000 472.780 15.260 ;
        RECT 505.180 15.000 505.440 15.260 ;
      LAYER met2 ;
        RECT 352.350 400.250 352.630 404.000 ;
        RECT 352.060 400.110 352.630 400.250 ;
        RECT 352.060 393.370 352.200 400.110 ;
        RECT 352.350 400.000 352.630 400.110 ;
        RECT 352.000 393.050 352.260 393.370 ;
        RECT 353.380 393.050 353.640 393.370 ;
        RECT 353.440 391.670 353.580 393.050 ;
        RECT 472.060 391.690 472.320 392.010 ;
        RECT 353.380 391.350 353.640 391.670 ;
        RECT 472.120 372.670 472.260 391.690 ;
        RECT 472.120 372.530 472.720 372.670 ;
        RECT 472.580 15.290 472.720 372.530 ;
        RECT 472.520 14.970 472.780 15.290 ;
        RECT 505.180 14.970 505.440 15.290 ;
        RECT 505.240 2.400 505.380 14.970 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.430 23.020 352.750 23.080 ;
        RECT 522.630 23.020 522.950 23.080 ;
        RECT 352.430 22.880 522.950 23.020 ;
        RECT 352.430 22.820 352.750 22.880 ;
        RECT 522.630 22.820 522.950 22.880 ;
      LAYER via ;
        RECT 352.460 22.820 352.720 23.080 ;
        RECT 522.660 22.820 522.920 23.080 ;
      LAYER met2 ;
        RECT 357.410 400.250 357.690 404.000 ;
        RECT 356.200 400.110 357.690 400.250 ;
        RECT 356.200 399.570 356.340 400.110 ;
        RECT 357.410 400.000 357.690 400.110 ;
        RECT 354.820 399.430 356.340 399.570 ;
        RECT 354.820 351.970 354.960 399.430 ;
        RECT 352.520 351.830 354.960 351.970 ;
        RECT 352.520 23.110 352.660 351.830 ;
        RECT 352.460 22.790 352.720 23.110 ;
        RECT 522.660 22.790 522.920 23.110 ;
        RECT 522.720 2.400 522.860 22.790 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 363.010 387.840 363.330 387.900 ;
        RECT 403.490 387.840 403.810 387.900 ;
        RECT 363.010 387.700 403.810 387.840 ;
        RECT 363.010 387.640 363.330 387.700 ;
        RECT 403.490 387.640 403.810 387.700 ;
        RECT 403.490 20.300 403.810 20.360 ;
        RECT 540.570 20.300 540.890 20.360 ;
        RECT 403.490 20.160 540.890 20.300 ;
        RECT 403.490 20.100 403.810 20.160 ;
        RECT 540.570 20.100 540.890 20.160 ;
      LAYER via ;
        RECT 363.040 387.640 363.300 387.900 ;
        RECT 403.520 387.640 403.780 387.900 ;
        RECT 403.520 20.100 403.780 20.360 ;
        RECT 540.600 20.100 540.860 20.360 ;
      LAYER met2 ;
        RECT 362.930 400.180 363.210 404.000 ;
        RECT 362.930 400.000 363.240 400.180 ;
        RECT 363.100 387.930 363.240 400.000 ;
        RECT 363.040 387.610 363.300 387.930 ;
        RECT 403.520 387.610 403.780 387.930 ;
        RECT 403.580 20.390 403.720 387.610 ;
        RECT 403.520 20.070 403.780 20.390 ;
        RECT 540.600 20.070 540.860 20.390 ;
        RECT 540.660 2.400 540.800 20.070 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 18.600 366.090 18.660 ;
        RECT 558.050 18.600 558.370 18.660 ;
        RECT 365.770 18.460 558.370 18.600 ;
        RECT 365.770 18.400 366.090 18.460 ;
        RECT 558.050 18.400 558.370 18.460 ;
      LAYER via ;
        RECT 365.800 18.400 366.060 18.660 ;
        RECT 558.080 18.400 558.340 18.660 ;
      LAYER met2 ;
        RECT 367.990 400.250 368.270 404.000 ;
        RECT 367.240 400.110 368.270 400.250 ;
        RECT 367.240 351.970 367.380 400.110 ;
        RECT 367.990 400.000 368.270 400.110 ;
        RECT 365.860 351.830 367.380 351.970 ;
        RECT 365.860 18.690 366.000 351.830 ;
        RECT 365.800 18.370 366.060 18.690 ;
        RECT 558.080 18.370 558.340 18.690 ;
        RECT 558.140 2.400 558.280 18.370 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 373.590 393.280 373.910 393.340 ;
        RECT 493.190 393.280 493.510 393.340 ;
        RECT 373.590 393.140 493.510 393.280 ;
        RECT 373.590 393.080 373.910 393.140 ;
        RECT 493.190 393.080 493.510 393.140 ;
        RECT 493.190 390.560 493.510 390.620 ;
        RECT 527.690 390.560 528.010 390.620 ;
        RECT 493.190 390.420 528.010 390.560 ;
        RECT 493.190 390.360 493.510 390.420 ;
        RECT 527.690 390.360 528.010 390.420 ;
        RECT 527.690 15.200 528.010 15.260 ;
        RECT 575.990 15.200 576.310 15.260 ;
        RECT 527.690 15.060 576.310 15.200 ;
        RECT 527.690 15.000 528.010 15.060 ;
        RECT 575.990 15.000 576.310 15.060 ;
      LAYER via ;
        RECT 373.620 393.080 373.880 393.340 ;
        RECT 493.220 393.080 493.480 393.340 ;
        RECT 493.220 390.360 493.480 390.620 ;
        RECT 527.720 390.360 527.980 390.620 ;
        RECT 527.720 15.000 527.980 15.260 ;
        RECT 576.020 15.000 576.280 15.260 ;
      LAYER met2 ;
        RECT 373.510 400.180 373.790 404.000 ;
        RECT 373.510 400.000 373.820 400.180 ;
        RECT 373.680 393.370 373.820 400.000 ;
        RECT 373.620 393.050 373.880 393.370 ;
        RECT 493.220 393.050 493.480 393.370 ;
        RECT 493.280 390.650 493.420 393.050 ;
        RECT 493.220 390.330 493.480 390.650 ;
        RECT 527.720 390.330 527.980 390.650 ;
        RECT 527.780 15.290 527.920 390.330 ;
        RECT 527.720 14.970 527.980 15.290 ;
        RECT 576.020 14.970 576.280 15.290 ;
        RECT 576.080 2.400 576.220 14.970 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203.850 20.300 204.170 20.360 ;
        RECT 221.790 20.300 222.110 20.360 ;
        RECT 203.850 20.160 222.110 20.300 ;
        RECT 203.850 20.100 204.170 20.160 ;
        RECT 221.790 20.100 222.110 20.160 ;
        RECT 85.170 19.620 85.490 19.680 ;
        RECT 85.170 19.480 202.700 19.620 ;
        RECT 85.170 19.420 85.490 19.480 ;
        RECT 202.560 19.340 202.700 19.480 ;
        RECT 202.470 19.080 202.790 19.340 ;
      LAYER via ;
        RECT 203.880 20.100 204.140 20.360 ;
        RECT 221.820 20.100 222.080 20.360 ;
        RECT 85.200 19.420 85.460 19.680 ;
        RECT 202.500 19.080 202.760 19.340 ;
      LAYER met2 ;
        RECT 225.390 400.250 225.670 404.000 ;
        RECT 224.180 400.110 225.670 400.250 ;
        RECT 224.180 399.570 224.320 400.110 ;
        RECT 225.390 400.000 225.670 400.110 ;
        RECT 223.720 399.430 224.320 399.570 ;
        RECT 223.720 303.670 223.860 399.430 ;
        RECT 221.880 303.530 223.860 303.670 ;
        RECT 221.880 20.390 222.020 303.530 ;
        RECT 203.880 20.070 204.140 20.390 ;
        RECT 221.820 20.070 222.080 20.390 ;
        RECT 85.200 19.390 85.460 19.710 ;
        RECT 203.940 19.450 204.080 20.070 ;
        RECT 85.260 2.400 85.400 19.390 ;
        RECT 202.560 19.370 204.080 19.450 ;
        RECT 202.500 19.310 204.080 19.370 ;
        RECT 202.500 19.050 202.760 19.310 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 376.280 372.990 376.340 ;
        RECT 377.730 376.280 378.050 376.340 ;
        RECT 372.670 376.140 378.050 376.280 ;
        RECT 372.670 376.080 372.990 376.140 ;
        RECT 377.730 376.080 378.050 376.140 ;
        RECT 372.670 17.920 372.990 17.980 ;
        RECT 593.930 17.920 594.250 17.980 ;
        RECT 372.670 17.780 594.250 17.920 ;
        RECT 372.670 17.720 372.990 17.780 ;
        RECT 593.930 17.720 594.250 17.780 ;
      LAYER via ;
        RECT 372.700 376.080 372.960 376.340 ;
        RECT 377.760 376.080 378.020 376.340 ;
        RECT 372.700 17.720 372.960 17.980 ;
        RECT 593.960 17.720 594.220 17.980 ;
      LAYER met2 ;
        RECT 379.030 400.250 379.310 404.000 ;
        RECT 377.820 400.110 379.310 400.250 ;
        RECT 377.820 376.370 377.960 400.110 ;
        RECT 379.030 400.000 379.310 400.110 ;
        RECT 372.700 376.050 372.960 376.370 ;
        RECT 377.760 376.050 378.020 376.370 ;
        RECT 372.760 18.010 372.900 376.050 ;
        RECT 372.700 17.690 372.960 18.010 ;
        RECT 593.960 17.690 594.220 18.010 ;
        RECT 594.020 2.400 594.160 17.690 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.950 33.220 381.270 33.280 ;
        RECT 532.750 33.220 533.070 33.280 ;
        RECT 380.950 33.080 533.070 33.220 ;
        RECT 380.950 33.020 381.270 33.080 ;
        RECT 532.750 33.020 533.070 33.080 ;
        RECT 532.750 16.900 533.070 16.960 ;
        RECT 611.410 16.900 611.730 16.960 ;
        RECT 532.750 16.760 611.730 16.900 ;
        RECT 532.750 16.700 533.070 16.760 ;
        RECT 611.410 16.700 611.730 16.760 ;
      LAYER via ;
        RECT 380.980 33.020 381.240 33.280 ;
        RECT 532.780 33.020 533.040 33.280 ;
        RECT 532.780 16.700 533.040 16.960 ;
        RECT 611.440 16.700 611.700 16.960 ;
      LAYER met2 ;
        RECT 384.090 400.250 384.370 404.000 ;
        RECT 383.340 400.110 384.370 400.250 ;
        RECT 383.340 324.370 383.480 400.110 ;
        RECT 384.090 400.000 384.370 400.110 ;
        RECT 381.040 324.230 383.480 324.370 ;
        RECT 381.040 33.310 381.180 324.230 ;
        RECT 380.980 32.990 381.240 33.310 ;
        RECT 532.780 32.990 533.040 33.310 ;
        RECT 532.840 16.990 532.980 32.990 ;
        RECT 532.780 16.670 533.040 16.990 ;
        RECT 611.440 16.670 611.700 16.990 ;
        RECT 611.500 2.400 611.640 16.670 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.690 375.940 229.010 376.000 ;
        RECT 231.450 375.940 231.770 376.000 ;
        RECT 228.690 375.800 231.770 375.940 ;
        RECT 228.690 375.740 229.010 375.800 ;
        RECT 231.450 375.740 231.770 375.800 ;
        RECT 109.090 16.900 109.410 16.960 ;
        RECT 228.690 16.900 229.010 16.960 ;
        RECT 109.090 16.760 229.010 16.900 ;
        RECT 109.090 16.700 109.410 16.760 ;
        RECT 228.690 16.700 229.010 16.760 ;
      LAYER via ;
        RECT 228.720 375.740 228.980 376.000 ;
        RECT 231.480 375.740 231.740 376.000 ;
        RECT 109.120 16.700 109.380 16.960 ;
        RECT 228.720 16.700 228.980 16.960 ;
      LAYER met2 ;
        RECT 232.290 400.250 232.570 404.000 ;
        RECT 231.540 400.110 232.570 400.250 ;
        RECT 231.540 376.030 231.680 400.110 ;
        RECT 232.290 400.000 232.570 400.110 ;
        RECT 228.720 375.710 228.980 376.030 ;
        RECT 231.480 375.710 231.740 376.030 ;
        RECT 228.780 16.990 228.920 375.710 ;
        RECT 109.120 16.670 109.380 16.990 ;
        RECT 228.720 16.670 228.980 16.990 ;
        RECT 109.180 2.400 109.320 16.670 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.550 24.040 132.870 24.100 ;
        RECT 235.130 24.040 235.450 24.100 ;
        RECT 132.550 23.900 235.450 24.040 ;
        RECT 132.550 23.840 132.870 23.900 ;
        RECT 235.130 23.840 235.450 23.900 ;
      LAYER via ;
        RECT 132.580 23.840 132.840 24.100 ;
        RECT 235.160 23.840 235.420 24.100 ;
      LAYER met2 ;
        RECT 239.650 400.250 239.930 404.000 ;
        RECT 238.440 400.110 239.930 400.250 ;
        RECT 238.440 351.970 238.580 400.110 ;
        RECT 239.650 400.000 239.930 400.110 ;
        RECT 235.220 351.830 238.580 351.970 ;
        RECT 235.220 24.130 235.360 351.830 ;
        RECT 132.580 23.810 132.840 24.130 ;
        RECT 235.160 23.810 235.420 24.130 ;
        RECT 132.640 2.400 132.780 23.810 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.490 375.940 242.810 376.000 ;
        RECT 243.870 375.940 244.190 376.000 ;
        RECT 242.490 375.800 244.190 375.940 ;
        RECT 242.490 375.740 242.810 375.800 ;
        RECT 243.870 375.740 244.190 375.800 ;
        RECT 150.490 24.380 150.810 24.440 ;
        RECT 242.490 24.380 242.810 24.440 ;
        RECT 150.490 24.240 242.810 24.380 ;
        RECT 150.490 24.180 150.810 24.240 ;
        RECT 242.490 24.180 242.810 24.240 ;
      LAYER via ;
        RECT 242.520 375.740 242.780 376.000 ;
        RECT 243.900 375.740 244.160 376.000 ;
        RECT 150.520 24.180 150.780 24.440 ;
        RECT 242.520 24.180 242.780 24.440 ;
      LAYER met2 ;
        RECT 245.170 400.250 245.450 404.000 ;
        RECT 243.960 400.110 245.450 400.250 ;
        RECT 243.960 376.030 244.100 400.110 ;
        RECT 245.170 400.000 245.450 400.110 ;
        RECT 242.520 375.710 242.780 376.030 ;
        RECT 243.900 375.710 244.160 376.030 ;
        RECT 242.580 24.470 242.720 375.710 ;
        RECT 150.520 24.150 150.780 24.470 ;
        RECT 242.520 24.150 242.780 24.470 ;
        RECT 150.580 2.400 150.720 24.150 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 167.970 24.720 168.290 24.780 ;
        RECT 249.850 24.720 250.170 24.780 ;
        RECT 167.970 24.580 250.170 24.720 ;
        RECT 167.970 24.520 168.290 24.580 ;
        RECT 249.850 24.520 250.170 24.580 ;
      LAYER via ;
        RECT 168.000 24.520 168.260 24.780 ;
        RECT 249.880 24.520 250.140 24.780 ;
      LAYER met2 ;
        RECT 250.230 400.180 250.510 404.000 ;
        RECT 250.230 400.000 250.540 400.180 ;
        RECT 250.400 303.670 250.540 400.000 ;
        RECT 249.940 303.530 250.540 303.670 ;
        RECT 249.940 24.810 250.080 303.530 ;
        RECT 168.000 24.490 168.260 24.810 ;
        RECT 249.880 24.490 250.140 24.810 ;
        RECT 168.060 2.400 168.200 24.490 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 179.470 393.280 179.790 393.340 ;
        RECT 255.830 393.280 256.150 393.340 ;
        RECT 179.470 393.140 256.150 393.280 ;
        RECT 179.470 393.080 179.790 393.140 ;
        RECT 255.830 393.080 256.150 393.140 ;
      LAYER via ;
        RECT 179.500 393.080 179.760 393.340 ;
        RECT 255.860 393.080 256.120 393.340 ;
      LAYER met2 ;
        RECT 255.750 400.180 256.030 404.000 ;
        RECT 255.750 400.000 256.060 400.180 ;
        RECT 255.920 393.370 256.060 400.000 ;
        RECT 179.500 393.050 179.760 393.370 ;
        RECT 255.860 393.050 256.120 393.370 ;
        RECT 179.560 82.870 179.700 393.050 ;
        RECT 179.560 82.730 183.840 82.870 ;
        RECT 183.700 1.770 183.840 82.730 ;
        RECT 185.790 1.770 186.350 2.400 ;
        RECT 183.700 1.630 186.350 1.770 ;
        RECT 185.790 -4.800 186.350 1.630 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203.390 15.200 203.710 15.260 ;
        RECT 255.830 15.200 256.150 15.260 ;
        RECT 203.390 15.060 256.150 15.200 ;
        RECT 203.390 15.000 203.710 15.060 ;
        RECT 255.830 15.000 256.150 15.060 ;
      LAYER via ;
        RECT 203.420 15.000 203.680 15.260 ;
        RECT 255.860 15.000 256.120 15.260 ;
      LAYER met2 ;
        RECT 261.270 400.250 261.550 404.000 ;
        RECT 260.060 400.110 261.550 400.250 ;
        RECT 260.060 388.010 260.200 400.110 ;
        RECT 261.270 400.000 261.550 400.110 ;
        RECT 255.920 387.870 260.200 388.010 ;
        RECT 255.920 15.290 256.060 387.870 ;
        RECT 203.420 14.970 203.680 15.290 ;
        RECT 255.860 14.970 256.120 15.290 ;
        RECT 203.480 2.400 203.620 14.970 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 224.640 17.440 244.560 17.580 ;
        RECT 221.330 17.240 221.650 17.300 ;
        RECT 224.640 17.240 224.780 17.440 ;
        RECT 221.330 17.100 224.780 17.240 ;
        RECT 244.420 17.240 244.560 17.440 ;
        RECT 263.650 17.240 263.970 17.300 ;
        RECT 244.420 17.100 263.970 17.240 ;
        RECT 221.330 17.040 221.650 17.100 ;
        RECT 263.650 17.040 263.970 17.100 ;
      LAYER via ;
        RECT 221.360 17.040 221.620 17.300 ;
        RECT 263.680 17.040 263.940 17.300 ;
      LAYER met2 ;
        RECT 266.330 400.250 266.610 404.000 ;
        RECT 265.120 400.110 266.610 400.250 ;
        RECT 265.120 386.480 265.260 400.110 ;
        RECT 266.330 400.000 266.610 400.110 ;
        RECT 263.740 386.340 265.260 386.480 ;
        RECT 263.740 17.330 263.880 386.340 ;
        RECT 221.360 17.010 221.620 17.330 ;
        RECT 263.680 17.010 263.940 17.330 ;
        RECT 221.420 2.400 221.560 17.010 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.870 389.880 14.190 389.940 ;
        RECT 205.690 389.880 206.010 389.940 ;
        RECT 13.870 389.740 206.010 389.880 ;
        RECT 13.870 389.680 14.190 389.740 ;
        RECT 205.690 389.680 206.010 389.740 ;
      LAYER via ;
        RECT 13.900 389.680 14.160 389.940 ;
        RECT 205.720 389.680 205.980 389.940 ;
      LAYER met2 ;
        RECT 205.610 400.180 205.890 404.000 ;
        RECT 205.610 400.000 205.920 400.180 ;
        RECT 205.780 389.970 205.920 400.000 ;
        RECT 13.900 389.650 14.160 389.970 ;
        RECT 205.720 389.650 205.980 389.970 ;
        RECT 13.960 82.870 14.100 389.650 ;
        RECT 13.960 82.730 18.240 82.870 ;
        RECT 18.100 1.770 18.240 82.730 ;
        RECT 20.190 1.770 20.750 2.400 ;
        RECT 18.100 1.630 20.750 1.770 ;
        RECT 20.190 -4.800 20.750 1.630 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 43.770 18.260 44.090 18.320 ;
        RECT 208.910 18.260 209.230 18.320 ;
        RECT 43.770 18.120 209.230 18.260 ;
        RECT 43.770 18.060 44.090 18.120 ;
        RECT 208.910 18.060 209.230 18.120 ;
      LAYER via ;
        RECT 43.800 18.060 44.060 18.320 ;
        RECT 208.940 18.060 209.200 18.320 ;
      LAYER met2 ;
        RECT 212.970 400.250 213.250 404.000 ;
        RECT 211.760 400.110 213.250 400.250 ;
        RECT 211.760 303.670 211.900 400.110 ;
        RECT 212.970 400.000 213.250 400.110 ;
        RECT 209.000 303.530 211.900 303.670 ;
        RECT 209.000 18.350 209.140 303.530 ;
        RECT 43.800 18.030 44.060 18.350 ;
        RECT 208.940 18.030 209.200 18.350 ;
        RECT 43.860 2.400 44.000 18.030 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.590 387.160 258.910 387.220 ;
        RECT 273.770 387.160 274.090 387.220 ;
        RECT 258.590 387.020 274.090 387.160 ;
        RECT 258.590 386.960 258.910 387.020 ;
        RECT 273.770 386.960 274.090 387.020 ;
        RECT 244.790 17.580 245.110 17.640 ;
        RECT 258.590 17.580 258.910 17.640 ;
        RECT 244.790 17.440 258.910 17.580 ;
        RECT 244.790 17.380 245.110 17.440 ;
        RECT 258.590 17.380 258.910 17.440 ;
      LAYER via ;
        RECT 258.620 386.960 258.880 387.220 ;
        RECT 273.800 386.960 274.060 387.220 ;
        RECT 244.820 17.380 245.080 17.640 ;
        RECT 258.620 17.380 258.880 17.640 ;
      LAYER met2 ;
        RECT 273.690 400.180 273.970 404.000 ;
        RECT 273.690 400.000 274.000 400.180 ;
        RECT 273.860 387.250 274.000 400.000 ;
        RECT 258.620 386.930 258.880 387.250 ;
        RECT 273.800 386.930 274.060 387.250 ;
        RECT 258.680 17.670 258.820 386.930 ;
        RECT 244.820 17.350 245.080 17.670 ;
        RECT 258.620 17.350 258.880 17.670 ;
        RECT 244.880 2.400 245.020 17.350 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 265.490 392.940 265.810 393.000 ;
        RECT 278.830 392.940 279.150 393.000 ;
        RECT 265.490 392.800 279.150 392.940 ;
        RECT 265.490 392.740 265.810 392.800 ;
        RECT 278.830 392.740 279.150 392.800 ;
      LAYER via ;
        RECT 265.520 392.740 265.780 393.000 ;
        RECT 278.860 392.740 279.120 393.000 ;
      LAYER met2 ;
        RECT 278.750 400.180 279.030 404.000 ;
        RECT 278.750 400.000 279.060 400.180 ;
        RECT 278.920 393.030 279.060 400.000 ;
        RECT 265.520 392.710 265.780 393.030 ;
        RECT 278.860 392.710 279.120 393.030 ;
        RECT 265.580 324.370 265.720 392.710 ;
        RECT 264.660 324.230 265.720 324.370 ;
        RECT 262.610 1.770 263.170 2.400 ;
        RECT 264.660 1.770 264.800 324.230 ;
        RECT 262.610 1.630 264.800 1.770 ;
        RECT 262.610 -4.800 263.170 1.630 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.270 400.250 284.550 404.000 ;
        RECT 283.980 400.110 284.550 400.250 ;
        RECT 283.980 373.050 284.120 400.110 ;
        RECT 284.270 400.000 284.550 400.110 ;
        RECT 283.520 372.910 284.120 373.050 ;
        RECT 283.520 14.010 283.660 372.910 ;
        RECT 282.600 13.870 283.660 14.010 ;
        RECT 280.090 1.770 280.650 2.400 ;
        RECT 282.600 1.770 282.740 13.870 ;
        RECT 280.090 1.630 282.740 1.770 ;
        RECT 280.090 -4.800 280.650 1.630 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 291.250 17.580 291.570 17.640 ;
        RECT 298.150 17.580 298.470 17.640 ;
        RECT 291.250 17.440 298.470 17.580 ;
        RECT 291.250 17.380 291.570 17.440 ;
        RECT 298.150 17.380 298.470 17.440 ;
      LAYER via ;
        RECT 291.280 17.380 291.540 17.640 ;
        RECT 298.180 17.380 298.440 17.640 ;
      LAYER met2 ;
        RECT 289.790 400.250 290.070 404.000 ;
        RECT 289.790 400.110 291.480 400.250 ;
        RECT 289.790 400.000 290.070 400.110 ;
        RECT 291.340 17.670 291.480 400.110 ;
        RECT 291.280 17.350 291.540 17.670 ;
        RECT 298.180 17.350 298.440 17.670 ;
        RECT 298.240 2.400 298.380 17.350 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.330 386.480 290.650 386.540 ;
        RECT 293.550 386.480 293.870 386.540 ;
        RECT 290.330 386.340 293.870 386.480 ;
        RECT 290.330 386.280 290.650 386.340 ;
        RECT 293.550 386.280 293.870 386.340 ;
        RECT 290.330 17.920 290.650 17.980 ;
        RECT 316.090 17.920 316.410 17.980 ;
        RECT 290.330 17.780 316.410 17.920 ;
        RECT 290.330 17.720 290.650 17.780 ;
        RECT 316.090 17.720 316.410 17.780 ;
      LAYER via ;
        RECT 290.360 386.280 290.620 386.540 ;
        RECT 293.580 386.280 293.840 386.540 ;
        RECT 290.360 17.720 290.620 17.980 ;
        RECT 316.120 17.720 316.380 17.980 ;
      LAYER met2 ;
        RECT 294.850 400.250 295.130 404.000 ;
        RECT 293.640 400.110 295.130 400.250 ;
        RECT 293.640 386.570 293.780 400.110 ;
        RECT 294.850 400.000 295.130 400.110 ;
        RECT 290.360 386.250 290.620 386.570 ;
        RECT 293.580 386.250 293.840 386.570 ;
        RECT 290.420 18.010 290.560 386.250 ;
        RECT 290.360 17.690 290.620 18.010 ;
        RECT 316.120 17.690 316.380 18.010 ;
        RECT 316.180 2.400 316.320 17.690 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.770 15.540 297.090 15.600 ;
        RECT 333.570 15.540 333.890 15.600 ;
        RECT 296.770 15.400 333.890 15.540 ;
        RECT 296.770 15.340 297.090 15.400 ;
        RECT 333.570 15.340 333.890 15.400 ;
      LAYER via ;
        RECT 296.800 15.340 297.060 15.600 ;
        RECT 333.600 15.340 333.860 15.600 ;
      LAYER met2 ;
        RECT 300.370 400.250 300.650 404.000 ;
        RECT 299.160 400.110 300.650 400.250 ;
        RECT 299.160 324.370 299.300 400.110 ;
        RECT 300.370 400.000 300.650 400.110 ;
        RECT 296.860 324.230 299.300 324.370 ;
        RECT 296.860 15.630 297.000 324.230 ;
        RECT 296.800 15.310 297.060 15.630 ;
        RECT 333.600 15.310 333.860 15.630 ;
        RECT 333.660 2.400 333.800 15.310 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 305.970 386.480 306.290 386.540 ;
        RECT 313.790 386.480 314.110 386.540 ;
        RECT 305.970 386.340 314.110 386.480 ;
        RECT 305.970 386.280 306.290 386.340 ;
        RECT 313.790 386.280 314.110 386.340 ;
        RECT 313.790 19.280 314.110 19.340 ;
        RECT 351.510 19.280 351.830 19.340 ;
        RECT 313.790 19.140 351.830 19.280 ;
        RECT 313.790 19.080 314.110 19.140 ;
        RECT 351.510 19.080 351.830 19.140 ;
      LAYER via ;
        RECT 306.000 386.280 306.260 386.540 ;
        RECT 313.820 386.280 314.080 386.540 ;
        RECT 313.820 19.080 314.080 19.340 ;
        RECT 351.540 19.080 351.800 19.340 ;
      LAYER met2 ;
        RECT 305.890 400.180 306.170 404.000 ;
        RECT 305.890 400.000 306.200 400.180 ;
        RECT 306.060 386.570 306.200 400.000 ;
        RECT 306.000 386.250 306.260 386.570 ;
        RECT 313.820 386.250 314.080 386.570 ;
        RECT 313.880 19.370 314.020 386.250 ;
        RECT 313.820 19.050 314.080 19.370 ;
        RECT 351.540 19.050 351.800 19.370 ;
        RECT 351.600 2.400 351.740 19.050 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.570 18.260 310.890 18.320 ;
        RECT 310.570 18.120 319.540 18.260 ;
        RECT 310.570 18.060 310.890 18.120 ;
        RECT 319.400 17.920 319.540 18.120 ;
        RECT 368.990 17.920 369.310 17.980 ;
        RECT 319.400 17.780 369.310 17.920 ;
        RECT 368.990 17.720 369.310 17.780 ;
      LAYER via ;
        RECT 310.600 18.060 310.860 18.320 ;
        RECT 369.020 17.720 369.280 17.980 ;
      LAYER met2 ;
        RECT 310.950 400.250 311.230 404.000 ;
        RECT 310.660 400.110 311.230 400.250 ;
        RECT 310.660 18.350 310.800 400.110 ;
        RECT 310.950 400.000 311.230 400.110 ;
        RECT 310.600 18.030 310.860 18.350 ;
        RECT 369.020 17.690 369.280 18.010 ;
        RECT 369.080 2.400 369.220 17.690 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.030 20.640 311.350 20.700 ;
        RECT 311.030 20.500 324.370 20.640 ;
        RECT 311.030 20.440 311.350 20.500 ;
        RECT 324.230 20.300 324.370 20.500 ;
        RECT 324.230 20.160 351.970 20.300 ;
        RECT 351.830 19.960 351.970 20.160 ;
        RECT 375.430 19.960 375.750 20.020 ;
        RECT 351.830 19.820 375.750 19.960 ;
        RECT 375.430 19.760 375.750 19.820 ;
        RECT 376.350 19.960 376.670 20.020 ;
        RECT 386.930 19.960 387.250 20.020 ;
        RECT 376.350 19.820 387.250 19.960 ;
        RECT 376.350 19.760 376.670 19.820 ;
        RECT 386.930 19.760 387.250 19.820 ;
      LAYER via ;
        RECT 311.060 20.440 311.320 20.700 ;
        RECT 375.460 19.760 375.720 20.020 ;
        RECT 376.380 19.760 376.640 20.020 ;
        RECT 386.960 19.760 387.220 20.020 ;
      LAYER met2 ;
        RECT 316.470 400.250 316.750 404.000 ;
        RECT 315.260 400.110 316.750 400.250 ;
        RECT 315.260 388.690 315.400 400.110 ;
        RECT 316.470 400.000 316.750 400.110 ;
        RECT 313.420 388.550 315.400 388.690 ;
        RECT 313.420 351.970 313.560 388.550 ;
        RECT 311.120 351.830 313.560 351.970 ;
        RECT 311.120 20.730 311.260 351.830 ;
        RECT 311.060 20.410 311.320 20.730 ;
        RECT 375.520 20.050 376.580 20.130 ;
        RECT 375.460 19.990 376.640 20.050 ;
        RECT 375.460 19.730 375.720 19.990 ;
        RECT 376.380 19.730 376.640 19.990 ;
        RECT 386.960 19.730 387.220 20.050 ;
        RECT 387.020 2.400 387.160 19.730 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.850 376.280 319.170 376.340 ;
        RECT 320.690 376.280 321.010 376.340 ;
        RECT 318.850 376.140 321.010 376.280 ;
        RECT 318.850 376.080 319.170 376.140 ;
        RECT 320.690 376.080 321.010 376.140 ;
        RECT 318.850 17.720 319.170 17.980 ;
        RECT 318.940 17.580 319.080 17.720 ;
        RECT 404.410 17.580 404.730 17.640 ;
        RECT 318.940 17.440 404.730 17.580 ;
        RECT 404.410 17.380 404.730 17.440 ;
      LAYER via ;
        RECT 318.880 376.080 319.140 376.340 ;
        RECT 320.720 376.080 320.980 376.340 ;
        RECT 318.880 17.720 319.140 17.980 ;
        RECT 404.440 17.380 404.700 17.640 ;
      LAYER met2 ;
        RECT 321.990 400.250 322.270 404.000 ;
        RECT 320.780 400.110 322.270 400.250 ;
        RECT 320.780 376.370 320.920 400.110 ;
        RECT 321.990 400.000 322.270 400.110 ;
        RECT 318.880 376.050 319.140 376.370 ;
        RECT 320.720 376.050 320.980 376.370 ;
        RECT 318.940 18.010 319.080 376.050 ;
        RECT 318.880 17.690 319.140 18.010 ;
        RECT 404.440 17.350 404.700 17.670 ;
        RECT 404.500 2.400 404.640 17.350 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.170 390.900 62.490 390.960 ;
        RECT 219.950 390.900 220.270 390.960 ;
        RECT 62.170 390.760 220.270 390.900 ;
        RECT 62.170 390.700 62.490 390.760 ;
        RECT 219.950 390.700 220.270 390.760 ;
      LAYER via ;
        RECT 62.200 390.700 62.460 390.960 ;
        RECT 219.980 390.700 220.240 390.960 ;
      LAYER met2 ;
        RECT 219.870 400.180 220.150 404.000 ;
        RECT 219.870 400.000 220.180 400.180 ;
        RECT 220.040 390.990 220.180 400.000 ;
        RECT 62.200 390.670 62.460 390.990 ;
        RECT 219.980 390.670 220.240 390.990 ;
        RECT 62.260 82.870 62.400 390.670 ;
        RECT 62.260 82.730 67.920 82.870 ;
        RECT 67.780 2.400 67.920 82.730 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.830 16.220 325.150 16.280 ;
        RECT 422.350 16.220 422.670 16.280 ;
        RECT 324.830 16.080 422.670 16.220 ;
        RECT 324.830 16.020 325.150 16.080 ;
        RECT 422.350 16.020 422.670 16.080 ;
      LAYER via ;
        RECT 324.860 16.020 325.120 16.280 ;
        RECT 422.380 16.020 422.640 16.280 ;
      LAYER met2 ;
        RECT 327.050 400.250 327.330 404.000 ;
        RECT 325.840 400.110 327.330 400.250 ;
        RECT 325.840 386.470 325.980 400.110 ;
        RECT 327.050 400.000 327.330 400.110 ;
        RECT 325.840 386.330 326.440 386.470 ;
        RECT 326.300 385.970 326.440 386.330 ;
        RECT 325.840 385.830 326.440 385.970 ;
        RECT 325.840 362.170 325.980 385.830 ;
        RECT 324.920 362.030 325.980 362.170 ;
        RECT 324.920 16.310 325.060 362.030 ;
        RECT 324.860 15.990 325.120 16.310 ;
        RECT 422.380 15.990 422.640 16.310 ;
        RECT 422.440 2.400 422.580 15.990 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.730 16.900 332.050 16.960 ;
        RECT 439.830 16.900 440.150 16.960 ;
        RECT 331.730 16.760 440.150 16.900 ;
        RECT 331.730 16.700 332.050 16.760 ;
        RECT 439.830 16.700 440.150 16.760 ;
      LAYER via ;
        RECT 331.760 16.700 332.020 16.960 ;
        RECT 439.860 16.700 440.120 16.960 ;
      LAYER met2 ;
        RECT 332.570 400.250 332.850 404.000 ;
        RECT 332.280 400.110 332.850 400.250 ;
        RECT 332.280 351.970 332.420 400.110 ;
        RECT 332.570 400.000 332.850 400.110 ;
        RECT 331.820 351.830 332.420 351.970 ;
        RECT 331.820 16.990 331.960 351.830 ;
        RECT 331.760 16.670 332.020 16.990 ;
        RECT 439.860 16.670 440.120 16.990 ;
        RECT 439.920 2.400 440.060 16.670 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 337.710 389.200 338.030 389.260 ;
        RECT 375.890 389.200 376.210 389.260 ;
        RECT 337.710 389.060 376.210 389.200 ;
        RECT 337.710 389.000 338.030 389.060 ;
        RECT 375.890 389.000 376.210 389.060 ;
        RECT 375.890 387.500 376.210 387.560 ;
        RECT 410.390 387.500 410.710 387.560 ;
        RECT 375.890 387.360 410.710 387.500 ;
        RECT 375.890 387.300 376.210 387.360 ;
        RECT 410.390 387.300 410.710 387.360 ;
        RECT 410.850 15.200 411.170 15.260 ;
        RECT 457.770 15.200 458.090 15.260 ;
        RECT 410.850 15.060 458.090 15.200 ;
        RECT 410.850 15.000 411.170 15.060 ;
        RECT 457.770 15.000 458.090 15.060 ;
      LAYER via ;
        RECT 337.740 389.000 338.000 389.260 ;
        RECT 375.920 389.000 376.180 389.260 ;
        RECT 375.920 387.300 376.180 387.560 ;
        RECT 410.420 387.300 410.680 387.560 ;
        RECT 410.880 15.000 411.140 15.260 ;
        RECT 457.800 15.000 458.060 15.260 ;
      LAYER met2 ;
        RECT 337.630 400.180 337.910 404.000 ;
        RECT 337.630 400.000 337.940 400.180 ;
        RECT 337.800 389.290 337.940 400.000 ;
        RECT 337.740 388.970 338.000 389.290 ;
        RECT 375.920 388.970 376.180 389.290 ;
        RECT 375.980 387.590 376.120 388.970 ;
        RECT 375.920 387.270 376.180 387.590 ;
        RECT 410.420 387.270 410.680 387.590 ;
        RECT 410.480 82.870 410.620 387.270 ;
        RECT 410.480 82.730 411.080 82.870 ;
        RECT 410.940 15.290 411.080 82.730 ;
        RECT 410.880 14.970 411.140 15.290 ;
        RECT 457.800 14.970 458.060 15.290 ;
        RECT 457.860 2.400 458.000 14.970 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 391.070 388.520 391.390 388.580 ;
        RECT 376.440 388.380 391.390 388.520 ;
        RECT 343.230 388.180 343.550 388.240 ;
        RECT 376.440 388.180 376.580 388.380 ;
        RECT 391.070 388.320 391.390 388.380 ;
        RECT 343.230 388.040 376.580 388.180 ;
        RECT 343.230 387.980 343.550 388.040 ;
        RECT 475.710 15.880 476.030 15.940 ;
        RECT 420.830 15.740 476.030 15.880 ;
        RECT 390.150 15.540 390.470 15.600 ;
        RECT 420.830 15.540 420.970 15.740 ;
        RECT 475.710 15.680 476.030 15.740 ;
        RECT 390.150 15.400 420.970 15.540 ;
        RECT 390.150 15.340 390.470 15.400 ;
      LAYER via ;
        RECT 343.260 387.980 343.520 388.240 ;
        RECT 391.100 388.320 391.360 388.580 ;
        RECT 390.180 15.340 390.440 15.600 ;
        RECT 475.740 15.680 476.000 15.940 ;
      LAYER met2 ;
        RECT 343.150 400.180 343.430 404.000 ;
        RECT 343.150 400.000 343.460 400.180 ;
        RECT 343.320 388.270 343.460 400.000 ;
        RECT 391.100 388.290 391.360 388.610 ;
        RECT 343.260 387.950 343.520 388.270 ;
        RECT 391.160 324.370 391.300 388.290 ;
        RECT 390.240 324.230 391.300 324.370 ;
        RECT 390.240 15.630 390.380 324.230 ;
        RECT 475.740 15.650 476.000 15.970 ;
        RECT 390.180 15.310 390.440 15.630 ;
        RECT 475.800 2.400 475.940 15.650 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.690 392.260 459.010 392.320 ;
        RECT 352.520 392.120 459.010 392.260 ;
        RECT 348.750 391.580 349.070 391.640 ;
        RECT 352.520 391.580 352.660 392.120 ;
        RECT 458.690 392.060 459.010 392.120 ;
        RECT 348.750 391.440 352.660 391.580 ;
        RECT 348.750 391.380 349.070 391.440 ;
        RECT 458.690 16.220 459.010 16.280 ;
        RECT 493.190 16.220 493.510 16.280 ;
        RECT 458.690 16.080 493.510 16.220 ;
        RECT 458.690 16.020 459.010 16.080 ;
        RECT 493.190 16.020 493.510 16.080 ;
      LAYER via ;
        RECT 348.780 391.380 349.040 391.640 ;
        RECT 458.720 392.060 458.980 392.320 ;
        RECT 458.720 16.020 458.980 16.280 ;
        RECT 493.220 16.020 493.480 16.280 ;
      LAYER met2 ;
        RECT 348.670 400.180 348.950 404.000 ;
        RECT 348.670 400.000 348.980 400.180 ;
        RECT 348.840 391.670 348.980 400.000 ;
        RECT 458.720 392.030 458.980 392.350 ;
        RECT 348.780 391.350 349.040 391.670 ;
        RECT 458.780 16.310 458.920 392.030 ;
        RECT 458.720 15.990 458.980 16.310 ;
        RECT 493.220 15.990 493.480 16.310 ;
        RECT 493.280 2.400 493.420 15.990 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 375.980 20.160 400.270 20.300 ;
        RECT 351.970 19.620 352.290 19.680 ;
        RECT 375.980 19.620 376.120 20.160 ;
        RECT 400.130 19.960 400.270 20.160 ;
        RECT 510.210 19.960 510.530 20.020 ;
        RECT 400.130 19.820 510.530 19.960 ;
        RECT 510.210 19.760 510.530 19.820 ;
        RECT 351.970 19.480 376.120 19.620 ;
        RECT 351.970 19.420 352.290 19.480 ;
      LAYER via ;
        RECT 352.000 19.420 352.260 19.680 ;
        RECT 510.240 19.760 510.500 20.020 ;
      LAYER met2 ;
        RECT 353.730 400.250 354.010 404.000 ;
        RECT 352.980 400.110 354.010 400.250 ;
        RECT 352.980 391.410 353.120 400.110 ;
        RECT 353.730 400.000 354.010 400.110 ;
        RECT 352.060 391.270 353.120 391.410 ;
        RECT 352.060 19.710 352.200 391.270 ;
        RECT 510.240 19.730 510.500 20.050 ;
        RECT 352.000 19.390 352.260 19.710 ;
        RECT 510.300 19.450 510.440 19.730 ;
        RECT 510.300 19.310 511.360 19.450 ;
        RECT 511.220 2.400 511.360 19.310 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.330 389.540 359.650 389.600 ;
        RECT 391.990 389.540 392.310 389.600 ;
        RECT 359.330 389.400 392.310 389.540 ;
        RECT 359.330 389.340 359.650 389.400 ;
        RECT 391.990 389.340 392.310 389.400 ;
        RECT 391.990 388.180 392.310 388.240 ;
        RECT 486.290 388.180 486.610 388.240 ;
        RECT 391.990 388.040 486.610 388.180 ;
        RECT 391.990 387.980 392.310 388.040 ;
        RECT 486.290 387.980 486.610 388.040 ;
        RECT 486.290 16.900 486.610 16.960 ;
        RECT 528.610 16.900 528.930 16.960 ;
        RECT 486.290 16.760 528.930 16.900 ;
        RECT 486.290 16.700 486.610 16.760 ;
        RECT 528.610 16.700 528.930 16.760 ;
      LAYER via ;
        RECT 359.360 389.340 359.620 389.600 ;
        RECT 392.020 389.340 392.280 389.600 ;
        RECT 392.020 387.980 392.280 388.240 ;
        RECT 486.320 387.980 486.580 388.240 ;
        RECT 486.320 16.700 486.580 16.960 ;
        RECT 528.640 16.700 528.900 16.960 ;
      LAYER met2 ;
        RECT 359.250 400.180 359.530 404.000 ;
        RECT 359.250 400.000 359.560 400.180 ;
        RECT 359.420 389.630 359.560 400.000 ;
        RECT 359.360 389.310 359.620 389.630 ;
        RECT 392.020 389.310 392.280 389.630 ;
        RECT 392.080 388.270 392.220 389.310 ;
        RECT 392.020 387.950 392.280 388.270 ;
        RECT 486.320 387.950 486.580 388.270 ;
        RECT 486.380 16.990 486.520 387.950 ;
        RECT 486.320 16.670 486.580 16.990 ;
        RECT 528.640 16.670 528.900 16.990 ;
        RECT 528.700 2.400 528.840 16.670 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.330 24.380 359.650 24.440 ;
        RECT 475.710 24.380 476.030 24.440 ;
        RECT 359.330 24.240 476.030 24.380 ;
        RECT 359.330 24.180 359.650 24.240 ;
        RECT 475.710 24.180 476.030 24.240 ;
        RECT 475.710 20.640 476.030 20.700 ;
        RECT 546.550 20.640 546.870 20.700 ;
        RECT 475.710 20.500 546.870 20.640 ;
        RECT 475.710 20.440 476.030 20.500 ;
        RECT 546.550 20.440 546.870 20.500 ;
      LAYER via ;
        RECT 359.360 24.180 359.620 24.440 ;
        RECT 475.740 24.180 476.000 24.440 ;
        RECT 475.740 20.440 476.000 20.700 ;
        RECT 546.580 20.440 546.840 20.700 ;
      LAYER met2 ;
        RECT 364.770 400.250 365.050 404.000 ;
        RECT 363.560 400.110 365.050 400.250 ;
        RECT 363.560 324.370 363.700 400.110 ;
        RECT 364.770 400.000 365.050 400.110 ;
        RECT 359.420 324.230 363.700 324.370 ;
        RECT 359.420 24.470 359.560 324.230 ;
        RECT 359.360 24.150 359.620 24.470 ;
        RECT 475.740 24.150 476.000 24.470 ;
        RECT 475.800 20.730 475.940 24.150 ;
        RECT 475.740 20.410 476.000 20.730 ;
        RECT 546.580 20.410 546.840 20.730 ;
        RECT 546.640 2.400 546.780 20.410 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 369.910 391.240 370.230 391.300 ;
        RECT 500.090 391.240 500.410 391.300 ;
        RECT 369.910 391.100 500.410 391.240 ;
        RECT 369.910 391.040 370.230 391.100 ;
        RECT 500.090 391.040 500.410 391.100 ;
        RECT 500.090 16.220 500.410 16.280 ;
        RECT 564.030 16.220 564.350 16.280 ;
        RECT 500.090 16.080 564.350 16.220 ;
        RECT 500.090 16.020 500.410 16.080 ;
        RECT 564.030 16.020 564.350 16.080 ;
      LAYER via ;
        RECT 369.940 391.040 370.200 391.300 ;
        RECT 500.120 391.040 500.380 391.300 ;
        RECT 500.120 16.020 500.380 16.280 ;
        RECT 564.060 16.020 564.320 16.280 ;
      LAYER met2 ;
        RECT 369.830 400.180 370.110 404.000 ;
        RECT 369.830 400.000 370.140 400.180 ;
        RECT 370.000 391.330 370.140 400.000 ;
        RECT 369.940 391.010 370.200 391.330 ;
        RECT 500.120 391.010 500.380 391.330 ;
        RECT 500.180 16.310 500.320 391.010 ;
        RECT 500.120 15.990 500.380 16.310 ;
        RECT 564.060 15.990 564.320 16.310 ;
        RECT 564.120 2.400 564.260 15.990 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 373.130 18.260 373.450 18.320 ;
        RECT 581.970 18.260 582.290 18.320 ;
        RECT 373.130 18.120 582.290 18.260 ;
        RECT 373.130 18.060 373.450 18.120 ;
        RECT 581.970 18.060 582.290 18.120 ;
      LAYER via ;
        RECT 373.160 18.060 373.420 18.320 ;
        RECT 582.000 18.060 582.260 18.320 ;
      LAYER met2 ;
        RECT 375.350 400.250 375.630 404.000 ;
        RECT 374.140 400.110 375.630 400.250 ;
        RECT 374.140 324.370 374.280 400.110 ;
        RECT 375.350 400.000 375.630 400.110 ;
        RECT 373.220 324.230 374.280 324.370 ;
        RECT 373.220 18.350 373.360 324.230 ;
        RECT 373.160 18.030 373.420 18.350 ;
        RECT 582.000 18.030 582.260 18.350 ;
        RECT 582.060 2.400 582.200 18.030 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 221.330 376.280 221.650 376.340 ;
        RECT 225.930 376.280 226.250 376.340 ;
        RECT 221.330 376.140 226.250 376.280 ;
        RECT 221.330 376.080 221.650 376.140 ;
        RECT 225.930 376.080 226.250 376.140 ;
        RECT 202.470 20.980 202.790 21.040 ;
        RECT 202.470 20.840 204.080 20.980 ;
        RECT 202.470 20.780 202.790 20.840 ;
        RECT 203.940 20.640 204.080 20.840 ;
        RECT 221.330 20.640 221.650 20.700 ;
        RECT 203.940 20.500 221.650 20.640 ;
        RECT 221.330 20.440 221.650 20.500 ;
        RECT 91.150 19.960 91.470 20.020 ;
        RECT 202.470 19.960 202.790 20.020 ;
        RECT 91.150 19.820 202.790 19.960 ;
        RECT 91.150 19.760 91.470 19.820 ;
        RECT 202.470 19.760 202.790 19.820 ;
      LAYER via ;
        RECT 221.360 376.080 221.620 376.340 ;
        RECT 225.960 376.080 226.220 376.340 ;
        RECT 202.500 20.780 202.760 21.040 ;
        RECT 221.360 20.440 221.620 20.700 ;
        RECT 91.180 19.760 91.440 20.020 ;
        RECT 202.500 19.760 202.760 20.020 ;
      LAYER met2 ;
        RECT 227.230 400.250 227.510 404.000 ;
        RECT 226.020 400.110 227.510 400.250 ;
        RECT 226.020 376.370 226.160 400.110 ;
        RECT 227.230 400.000 227.510 400.110 ;
        RECT 221.360 376.050 221.620 376.370 ;
        RECT 225.960 376.050 226.220 376.370 ;
        RECT 202.500 20.750 202.760 21.070 ;
        RECT 202.560 20.050 202.700 20.750 ;
        RECT 221.420 20.730 221.560 376.050 ;
        RECT 221.360 20.410 221.620 20.730 ;
        RECT 91.180 19.730 91.440 20.050 ;
        RECT 202.500 19.730 202.760 20.050 ;
        RECT 91.240 2.400 91.380 19.730 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.950 392.600 381.270 392.660 ;
        RECT 401.190 392.600 401.510 392.660 ;
        RECT 380.950 392.460 401.510 392.600 ;
        RECT 380.950 392.400 381.270 392.460 ;
        RECT 401.190 392.400 401.510 392.460 ;
        RECT 401.190 389.540 401.510 389.600 ;
        RECT 535.510 389.540 535.830 389.600 ;
        RECT 401.190 389.400 535.830 389.540 ;
        RECT 401.190 389.340 401.510 389.400 ;
        RECT 535.510 389.340 535.830 389.400 ;
        RECT 535.050 15.540 535.370 15.600 ;
        RECT 599.450 15.540 599.770 15.600 ;
        RECT 535.050 15.400 599.770 15.540 ;
        RECT 535.050 15.340 535.370 15.400 ;
        RECT 599.450 15.340 599.770 15.400 ;
      LAYER via ;
        RECT 380.980 392.400 381.240 392.660 ;
        RECT 401.220 392.400 401.480 392.660 ;
        RECT 401.220 389.340 401.480 389.600 ;
        RECT 535.540 389.340 535.800 389.600 ;
        RECT 535.080 15.340 535.340 15.600 ;
        RECT 599.480 15.340 599.740 15.600 ;
      LAYER met2 ;
        RECT 380.870 400.180 381.150 404.000 ;
        RECT 380.870 400.000 381.180 400.180 ;
        RECT 381.040 392.690 381.180 400.000 ;
        RECT 380.980 392.370 381.240 392.690 ;
        RECT 401.220 392.370 401.480 392.690 ;
        RECT 401.280 389.630 401.420 392.370 ;
        RECT 401.220 389.310 401.480 389.630 ;
        RECT 535.540 389.310 535.800 389.630 ;
        RECT 535.600 324.370 535.740 389.310 ;
        RECT 534.680 324.230 535.740 324.370 ;
        RECT 534.680 82.870 534.820 324.230 ;
        RECT 534.680 82.730 535.280 82.870 ;
        RECT 535.140 15.630 535.280 82.730 ;
        RECT 535.080 15.310 535.340 15.630 ;
        RECT 599.480 15.310 599.740 15.630 ;
        RECT 599.540 2.400 599.680 15.310 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.030 376.280 380.350 376.340 ;
        RECT 384.630 376.280 384.950 376.340 ;
        RECT 380.030 376.140 384.950 376.280 ;
        RECT 380.030 376.080 380.350 376.140 ;
        RECT 384.630 376.080 384.950 376.140 ;
        RECT 380.030 18.940 380.350 19.000 ;
        RECT 617.390 18.940 617.710 19.000 ;
        RECT 380.030 18.800 617.710 18.940 ;
        RECT 380.030 18.740 380.350 18.800 ;
        RECT 617.390 18.740 617.710 18.800 ;
      LAYER via ;
        RECT 380.060 376.080 380.320 376.340 ;
        RECT 384.660 376.080 384.920 376.340 ;
        RECT 380.060 18.740 380.320 19.000 ;
        RECT 617.420 18.740 617.680 19.000 ;
      LAYER met2 ;
        RECT 385.930 400.250 386.210 404.000 ;
        RECT 384.720 400.110 386.210 400.250 ;
        RECT 384.720 376.370 384.860 400.110 ;
        RECT 385.930 400.000 386.210 400.110 ;
        RECT 380.060 376.050 380.320 376.370 ;
        RECT 384.660 376.050 384.920 376.370 ;
        RECT 380.120 19.030 380.260 376.050 ;
        RECT 380.060 18.710 380.320 19.030 ;
        RECT 617.420 18.710 617.680 19.030 ;
        RECT 617.480 2.400 617.620 18.710 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 110.470 391.920 110.790 391.980 ;
        RECT 234.210 391.920 234.530 391.980 ;
        RECT 110.470 391.780 234.530 391.920 ;
        RECT 110.470 391.720 110.790 391.780 ;
        RECT 234.210 391.720 234.530 391.780 ;
      LAYER via ;
        RECT 110.500 391.720 110.760 391.980 ;
        RECT 234.240 391.720 234.500 391.980 ;
      LAYER met2 ;
        RECT 234.130 400.180 234.410 404.000 ;
        RECT 234.130 400.000 234.440 400.180 ;
        RECT 234.300 392.010 234.440 400.000 ;
        RECT 110.500 391.690 110.760 392.010 ;
        RECT 234.240 391.690 234.500 392.010 ;
        RECT 110.560 82.870 110.700 391.690 ;
        RECT 110.560 82.730 113.000 82.870 ;
        RECT 112.860 1.770 113.000 82.730 ;
        RECT 114.950 1.770 115.510 2.400 ;
        RECT 112.860 1.630 115.510 1.770 ;
        RECT 114.950 -4.800 115.510 1.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 138.530 16.220 138.850 16.280 ;
        RECT 138.530 16.080 233.060 16.220 ;
        RECT 138.530 16.020 138.850 16.080 ;
        RECT 232.920 15.880 233.060 16.080 ;
        RECT 242.950 15.880 243.270 15.940 ;
        RECT 232.920 15.740 243.270 15.880 ;
        RECT 242.950 15.680 243.270 15.740 ;
      LAYER via ;
        RECT 138.560 16.020 138.820 16.280 ;
        RECT 242.980 15.680 243.240 15.940 ;
      LAYER met2 ;
        RECT 241.490 400.250 241.770 404.000 ;
        RECT 241.490 400.110 243.180 400.250 ;
        RECT 241.490 400.000 241.770 400.110 ;
        RECT 138.560 15.990 138.820 16.310 ;
        RECT 138.620 2.400 138.760 15.990 ;
        RECT 243.040 15.970 243.180 400.110 ;
        RECT 242.980 15.650 243.240 15.970 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 151.870 392.940 152.190 393.000 ;
        RECT 246.630 392.940 246.950 393.000 ;
        RECT 151.870 392.800 246.950 392.940 ;
        RECT 151.870 392.740 152.190 392.800 ;
        RECT 246.630 392.740 246.950 392.800 ;
      LAYER via ;
        RECT 151.900 392.740 152.160 393.000 ;
        RECT 246.660 392.740 246.920 393.000 ;
      LAYER met2 ;
        RECT 246.550 400.180 246.830 404.000 ;
        RECT 246.550 400.000 246.860 400.180 ;
        RECT 246.720 393.030 246.860 400.000 ;
        RECT 151.900 392.710 152.160 393.030 ;
        RECT 246.660 392.710 246.920 393.030 ;
        RECT 151.960 82.870 152.100 392.710 ;
        RECT 151.960 82.730 154.400 82.870 ;
        RECT 154.260 1.770 154.400 82.730 ;
        RECT 156.350 1.770 156.910 2.400 ;
        RECT 154.260 1.630 156.910 1.770 ;
        RECT 156.350 -4.800 156.910 1.630 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 249.390 375.940 249.710 376.000 ;
        RECT 250.770 375.940 251.090 376.000 ;
        RECT 249.390 375.800 251.090 375.940 ;
        RECT 249.390 375.740 249.710 375.800 ;
        RECT 250.770 375.740 251.090 375.800 ;
        RECT 232.370 18.260 232.690 18.320 ;
        RECT 249.390 18.260 249.710 18.320 ;
        RECT 232.370 18.120 249.710 18.260 ;
        RECT 232.370 18.060 232.690 18.120 ;
        RECT 249.390 18.060 249.710 18.120 ;
        RECT 173.950 15.880 174.270 15.940 ;
        RECT 232.370 15.880 232.690 15.940 ;
        RECT 173.950 15.740 232.690 15.880 ;
        RECT 173.950 15.680 174.270 15.740 ;
        RECT 232.370 15.680 232.690 15.740 ;
      LAYER via ;
        RECT 249.420 375.740 249.680 376.000 ;
        RECT 250.800 375.740 251.060 376.000 ;
        RECT 232.400 18.060 232.660 18.320 ;
        RECT 249.420 18.060 249.680 18.320 ;
        RECT 173.980 15.680 174.240 15.940 ;
        RECT 232.400 15.680 232.660 15.940 ;
      LAYER met2 ;
        RECT 252.070 400.250 252.350 404.000 ;
        RECT 250.860 400.110 252.350 400.250 ;
        RECT 250.860 376.030 251.000 400.110 ;
        RECT 252.070 400.000 252.350 400.110 ;
        RECT 249.420 375.710 249.680 376.030 ;
        RECT 250.800 375.710 251.060 376.030 ;
        RECT 249.480 18.350 249.620 375.710 ;
        RECT 232.400 18.030 232.660 18.350 ;
        RECT 249.420 18.030 249.680 18.350 ;
        RECT 232.460 15.970 232.600 18.030 ;
        RECT 173.980 15.650 174.240 15.970 ;
        RECT 232.400 15.650 232.660 15.970 ;
        RECT 174.040 2.400 174.180 15.650 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 186.370 389.540 186.690 389.600 ;
        RECT 257.670 389.540 257.990 389.600 ;
        RECT 186.370 389.400 257.990 389.540 ;
        RECT 186.370 389.340 186.690 389.400 ;
        RECT 257.670 389.340 257.990 389.400 ;
      LAYER via ;
        RECT 186.400 389.340 186.660 389.600 ;
        RECT 257.700 389.340 257.960 389.600 ;
      LAYER met2 ;
        RECT 257.590 400.180 257.870 404.000 ;
        RECT 257.590 400.000 257.900 400.180 ;
        RECT 257.760 389.630 257.900 400.000 ;
        RECT 186.400 389.310 186.660 389.630 ;
        RECT 257.700 389.310 257.960 389.630 ;
        RECT 186.460 82.870 186.600 389.310 ;
        RECT 186.460 82.730 192.120 82.870 ;
        RECT 191.980 2.400 192.120 82.730 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 238.810 387.500 239.130 387.560 ;
        RECT 262.270 387.500 262.590 387.560 ;
        RECT 238.810 387.360 262.590 387.500 ;
        RECT 238.810 387.300 239.130 387.360 ;
        RECT 262.270 387.300 262.590 387.360 ;
        RECT 209.370 19.960 209.690 20.020 ;
        RECT 237.890 19.960 238.210 20.020 ;
        RECT 209.370 19.820 238.210 19.960 ;
        RECT 209.370 19.760 209.690 19.820 ;
        RECT 237.890 19.760 238.210 19.820 ;
      LAYER via ;
        RECT 238.840 387.300 239.100 387.560 ;
        RECT 262.300 387.300 262.560 387.560 ;
        RECT 209.400 19.760 209.660 20.020 ;
        RECT 237.920 19.760 238.180 20.020 ;
      LAYER met2 ;
        RECT 262.650 400.250 262.930 404.000 ;
        RECT 262.360 400.110 262.930 400.250 ;
        RECT 262.360 387.590 262.500 400.110 ;
        RECT 262.650 400.000 262.930 400.110 ;
        RECT 238.840 387.270 239.100 387.590 ;
        RECT 262.300 387.270 262.560 387.590 ;
        RECT 238.900 303.670 239.040 387.270 ;
        RECT 237.980 303.530 239.040 303.670 ;
        RECT 237.980 20.050 238.120 303.530 ;
        RECT 209.400 19.730 209.660 20.050 ;
        RECT 237.920 19.730 238.180 20.050 ;
        RECT 209.460 2.400 209.600 19.730 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 263.190 386.480 263.510 386.540 ;
        RECT 266.870 386.480 267.190 386.540 ;
        RECT 263.190 386.340 267.190 386.480 ;
        RECT 263.190 386.280 263.510 386.340 ;
        RECT 266.870 386.280 267.190 386.340 ;
        RECT 227.310 17.240 227.630 17.300 ;
        RECT 227.310 17.100 244.100 17.240 ;
        RECT 227.310 17.040 227.630 17.100 ;
        RECT 243.960 16.900 244.100 17.100 ;
        RECT 263.190 16.900 263.510 16.960 ;
        RECT 243.960 16.760 263.510 16.900 ;
        RECT 263.190 16.700 263.510 16.760 ;
      LAYER via ;
        RECT 263.220 386.280 263.480 386.540 ;
        RECT 266.900 386.280 267.160 386.540 ;
        RECT 227.340 17.040 227.600 17.300 ;
        RECT 263.220 16.700 263.480 16.960 ;
      LAYER met2 ;
        RECT 268.170 400.250 268.450 404.000 ;
        RECT 266.960 400.110 268.450 400.250 ;
        RECT 266.960 386.570 267.100 400.110 ;
        RECT 268.170 400.000 268.450 400.110 ;
        RECT 263.220 386.250 263.480 386.570 ;
        RECT 266.900 386.250 267.160 386.570 ;
        RECT 227.340 17.010 227.600 17.330 ;
        RECT 227.400 2.400 227.540 17.010 ;
        RECT 263.280 16.990 263.420 386.250 ;
        RECT 263.220 16.670 263.480 16.990 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 49.750 18.600 50.070 18.660 ;
        RECT 196.030 18.600 196.350 18.660 ;
        RECT 49.750 18.460 196.350 18.600 ;
        RECT 49.750 18.400 50.070 18.460 ;
        RECT 196.030 18.400 196.350 18.460 ;
        RECT 196.030 14.860 196.350 14.920 ;
        RECT 215.810 14.860 216.130 14.920 ;
        RECT 196.030 14.720 216.130 14.860 ;
        RECT 196.030 14.660 196.350 14.720 ;
        RECT 215.810 14.660 216.130 14.720 ;
      LAYER via ;
        RECT 49.780 18.400 50.040 18.660 ;
        RECT 196.060 18.400 196.320 18.660 ;
        RECT 196.060 14.660 196.320 14.920 ;
        RECT 215.840 14.660 216.100 14.920 ;
      LAYER met2 ;
        RECT 214.810 400.250 215.090 404.000 ;
        RECT 214.810 400.110 215.580 400.250 ;
        RECT 214.810 400.000 215.090 400.110 ;
        RECT 215.440 338.170 215.580 400.110 ;
        RECT 214.980 338.030 215.580 338.170 ;
        RECT 214.980 314.570 215.120 338.030 ;
        RECT 214.980 314.430 215.580 314.570 ;
        RECT 215.440 82.870 215.580 314.430 ;
        RECT 215.440 82.730 216.040 82.870 ;
        RECT 49.780 18.370 50.040 18.690 ;
        RECT 196.060 18.370 196.320 18.690 ;
        RECT 49.840 2.400 49.980 18.370 ;
        RECT 196.120 14.950 196.260 18.370 ;
        RECT 215.900 14.950 216.040 82.730 ;
        RECT 196.060 14.630 196.320 14.950 ;
        RECT 215.840 14.630 216.100 14.950 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.470 387.840 248.790 387.900 ;
        RECT 275.610 387.840 275.930 387.900 ;
        RECT 248.470 387.700 275.930 387.840 ;
        RECT 248.470 387.640 248.790 387.700 ;
        RECT 275.610 387.640 275.930 387.700 ;
      LAYER via ;
        RECT 248.500 387.640 248.760 387.900 ;
        RECT 275.640 387.640 275.900 387.900 ;
      LAYER met2 ;
        RECT 275.530 400.180 275.810 404.000 ;
        RECT 275.530 400.000 275.840 400.180 ;
        RECT 275.700 387.930 275.840 400.000 ;
        RECT 248.500 387.610 248.760 387.930 ;
        RECT 275.640 387.610 275.900 387.930 ;
        RECT 248.560 14.690 248.700 387.610 ;
        RECT 248.560 14.550 251.000 14.690 ;
        RECT 250.860 2.400 251.000 14.550 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 262.730 392.600 263.050 392.660 ;
        RECT 280.670 392.600 280.990 392.660 ;
        RECT 262.730 392.460 280.990 392.600 ;
        RECT 262.730 392.400 263.050 392.460 ;
        RECT 280.670 392.400 280.990 392.460 ;
        RECT 262.730 17.580 263.050 17.640 ;
        RECT 266.870 17.580 267.190 17.640 ;
        RECT 262.730 17.440 267.190 17.580 ;
        RECT 262.730 17.380 263.050 17.440 ;
        RECT 266.870 17.380 267.190 17.440 ;
      LAYER via ;
        RECT 262.760 392.400 263.020 392.660 ;
        RECT 280.700 392.400 280.960 392.660 ;
        RECT 262.760 17.380 263.020 17.640 ;
        RECT 266.900 17.380 267.160 17.640 ;
      LAYER met2 ;
        RECT 280.590 400.180 280.870 404.000 ;
        RECT 280.590 400.000 280.900 400.180 ;
        RECT 280.760 392.690 280.900 400.000 ;
        RECT 262.760 392.370 263.020 392.690 ;
        RECT 280.700 392.370 280.960 392.690 ;
        RECT 262.820 17.670 262.960 392.370 ;
        RECT 262.760 17.350 263.020 17.670 ;
        RECT 266.900 17.350 267.160 17.670 ;
        RECT 266.960 1.770 267.100 17.350 ;
        RECT 268.590 1.770 269.150 2.400 ;
        RECT 266.960 1.630 269.150 1.770 ;
        RECT 268.590 -4.800 269.150 1.630 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.970 386.480 283.290 386.540 ;
        RECT 284.810 386.480 285.130 386.540 ;
        RECT 282.970 386.340 285.130 386.480 ;
        RECT 282.970 386.280 283.290 386.340 ;
        RECT 284.810 386.280 285.130 386.340 ;
        RECT 282.970 17.580 283.290 17.640 ;
        RECT 284.350 17.580 284.670 17.640 ;
        RECT 282.970 17.440 284.670 17.580 ;
        RECT 282.970 17.380 283.290 17.440 ;
        RECT 284.350 17.380 284.670 17.440 ;
      LAYER via ;
        RECT 283.000 386.280 283.260 386.540 ;
        RECT 284.840 386.280 285.100 386.540 ;
        RECT 283.000 17.380 283.260 17.640 ;
        RECT 284.380 17.380 284.640 17.640 ;
      LAYER met2 ;
        RECT 286.110 400.250 286.390 404.000 ;
        RECT 284.900 400.110 286.390 400.250 ;
        RECT 284.900 386.570 285.040 400.110 ;
        RECT 286.110 400.000 286.390 400.110 ;
        RECT 283.000 386.250 283.260 386.570 ;
        RECT 284.840 386.250 285.100 386.570 ;
        RECT 283.060 17.670 283.200 386.250 ;
        RECT 283.000 17.350 283.260 17.670 ;
        RECT 284.380 17.350 284.640 17.670 ;
        RECT 284.440 1.770 284.580 17.350 ;
        RECT 286.070 1.770 286.630 2.400 ;
        RECT 284.440 1.630 286.630 1.770 ;
        RECT 286.070 -4.800 286.630 1.630 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 291.710 387.160 292.030 387.220 ;
        RECT 299.990 387.160 300.310 387.220 ;
        RECT 291.710 387.020 300.310 387.160 ;
        RECT 291.710 386.960 292.030 387.020 ;
        RECT 299.990 386.960 300.310 387.020 ;
        RECT 299.990 17.580 300.310 17.640 ;
        RECT 304.130 17.580 304.450 17.640 ;
        RECT 299.990 17.440 304.450 17.580 ;
        RECT 299.990 17.380 300.310 17.440 ;
        RECT 304.130 17.380 304.450 17.440 ;
      LAYER via ;
        RECT 291.740 386.960 292.000 387.220 ;
        RECT 300.020 386.960 300.280 387.220 ;
        RECT 300.020 17.380 300.280 17.640 ;
        RECT 304.160 17.380 304.420 17.640 ;
      LAYER met2 ;
        RECT 291.630 400.180 291.910 404.000 ;
        RECT 291.630 400.000 291.940 400.180 ;
        RECT 291.800 387.250 291.940 400.000 ;
        RECT 291.740 386.930 292.000 387.250 ;
        RECT 300.020 386.930 300.280 387.250 ;
        RECT 300.080 17.670 300.220 386.930 ;
        RECT 300.020 17.350 300.280 17.670 ;
        RECT 304.160 17.350 304.420 17.670 ;
        RECT 304.220 2.400 304.360 17.350 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.770 387.840 297.090 387.900 ;
        RECT 317.470 387.840 317.790 387.900 ;
        RECT 296.770 387.700 317.790 387.840 ;
        RECT 296.770 387.640 297.090 387.700 ;
        RECT 317.470 387.640 317.790 387.700 ;
      LAYER via ;
        RECT 296.800 387.640 297.060 387.900 ;
        RECT 317.500 387.640 317.760 387.900 ;
      LAYER met2 ;
        RECT 296.690 400.180 296.970 404.000 ;
        RECT 296.690 400.000 297.000 400.180 ;
        RECT 296.860 387.930 297.000 400.000 ;
        RECT 296.800 387.610 297.060 387.930 ;
        RECT 317.500 387.610 317.760 387.930 ;
        RECT 317.560 17.410 317.700 387.610 ;
        RECT 317.560 17.270 321.840 17.410 ;
        RECT 321.700 2.400 321.840 17.270 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 302.290 389.880 302.610 389.940 ;
        RECT 338.170 389.880 338.490 389.940 ;
        RECT 302.290 389.740 338.490 389.880 ;
        RECT 302.290 389.680 302.610 389.740 ;
        RECT 338.170 389.680 338.490 389.740 ;
      LAYER via ;
        RECT 302.320 389.680 302.580 389.940 ;
        RECT 338.200 389.680 338.460 389.940 ;
      LAYER met2 ;
        RECT 302.210 400.180 302.490 404.000 ;
        RECT 302.210 400.000 302.520 400.180 ;
        RECT 302.380 389.970 302.520 400.000 ;
        RECT 302.320 389.650 302.580 389.970 ;
        RECT 338.200 389.650 338.460 389.970 ;
        RECT 338.260 1.770 338.400 389.650 ;
        RECT 339.430 1.770 339.990 2.400 ;
        RECT 338.260 1.630 339.990 1.770 ;
        RECT 339.430 -4.800 339.990 1.630 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.670 376.280 303.990 376.340 ;
        RECT 306.430 376.280 306.750 376.340 ;
        RECT 303.670 376.140 306.750 376.280 ;
        RECT 303.670 376.080 303.990 376.140 ;
        RECT 306.430 376.080 306.750 376.140 ;
        RECT 303.670 19.620 303.990 19.680 ;
        RECT 320.230 19.620 320.550 19.680 ;
        RECT 303.670 19.480 320.550 19.620 ;
        RECT 303.670 19.420 303.990 19.480 ;
        RECT 320.230 19.420 320.550 19.480 ;
        RECT 320.230 18.600 320.550 18.660 ;
        RECT 357.490 18.600 357.810 18.660 ;
        RECT 320.230 18.460 357.810 18.600 ;
        RECT 320.230 18.400 320.550 18.460 ;
        RECT 357.490 18.400 357.810 18.460 ;
      LAYER via ;
        RECT 303.700 376.080 303.960 376.340 ;
        RECT 306.460 376.080 306.720 376.340 ;
        RECT 303.700 19.420 303.960 19.680 ;
        RECT 320.260 19.420 320.520 19.680 ;
        RECT 320.260 18.400 320.520 18.660 ;
        RECT 357.520 18.400 357.780 18.660 ;
      LAYER met2 ;
        RECT 307.270 400.250 307.550 404.000 ;
        RECT 306.520 400.110 307.550 400.250 ;
        RECT 306.520 376.370 306.660 400.110 ;
        RECT 307.270 400.000 307.550 400.110 ;
        RECT 303.700 376.050 303.960 376.370 ;
        RECT 306.460 376.050 306.720 376.370 ;
        RECT 303.760 19.710 303.900 376.050 ;
        RECT 303.700 19.390 303.960 19.710 ;
        RECT 320.260 19.390 320.520 19.710 ;
        RECT 320.320 18.690 320.460 19.390 ;
        RECT 320.260 18.370 320.520 18.690 ;
        RECT 357.520 18.370 357.780 18.690 ;
        RECT 357.580 2.400 357.720 18.370 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 312.870 390.560 313.190 390.620 ;
        RECT 355.190 390.560 355.510 390.620 ;
        RECT 312.870 390.420 355.510 390.560 ;
        RECT 312.870 390.360 313.190 390.420 ;
        RECT 355.190 390.360 355.510 390.420 ;
        RECT 355.190 20.300 355.510 20.360 ;
        RECT 374.970 20.300 375.290 20.360 ;
        RECT 355.190 20.160 375.290 20.300 ;
        RECT 355.190 20.100 355.510 20.160 ;
        RECT 374.970 20.100 375.290 20.160 ;
      LAYER via ;
        RECT 312.900 390.360 313.160 390.620 ;
        RECT 355.220 390.360 355.480 390.620 ;
        RECT 355.220 20.100 355.480 20.360 ;
        RECT 375.000 20.100 375.260 20.360 ;
      LAYER met2 ;
        RECT 312.790 400.180 313.070 404.000 ;
        RECT 312.790 400.000 313.100 400.180 ;
        RECT 312.960 390.650 313.100 400.000 ;
        RECT 312.900 390.330 313.160 390.650 ;
        RECT 355.220 390.330 355.480 390.650 ;
        RECT 355.280 20.390 355.420 390.330 ;
        RECT 355.220 20.070 355.480 20.390 ;
        RECT 375.000 20.070 375.260 20.390 ;
        RECT 375.060 2.400 375.200 20.070 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.390 20.300 318.710 20.360 ;
        RECT 322.070 20.300 322.390 20.360 ;
        RECT 318.390 20.160 322.390 20.300 ;
        RECT 318.390 20.100 318.710 20.160 ;
        RECT 322.070 20.100 322.390 20.160 ;
        RECT 322.070 15.880 322.390 15.940 ;
        RECT 392.910 15.880 393.230 15.940 ;
        RECT 322.070 15.740 393.230 15.880 ;
        RECT 322.070 15.680 322.390 15.740 ;
        RECT 392.910 15.680 393.230 15.740 ;
      LAYER via ;
        RECT 318.420 20.100 318.680 20.360 ;
        RECT 322.100 20.100 322.360 20.360 ;
        RECT 322.100 15.680 322.360 15.940 ;
        RECT 392.940 15.680 393.200 15.940 ;
      LAYER met2 ;
        RECT 318.310 400.180 318.590 404.000 ;
        RECT 318.310 400.000 318.620 400.180 ;
        RECT 318.480 20.390 318.620 400.000 ;
        RECT 318.420 20.070 318.680 20.390 ;
        RECT 322.100 20.070 322.360 20.390 ;
        RECT 322.160 15.970 322.300 20.070 ;
        RECT 322.100 15.650 322.360 15.970 ;
        RECT 392.940 15.650 393.200 15.970 ;
        RECT 393.000 2.400 393.140 15.650 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.930 375.940 318.250 376.000 ;
        RECT 322.530 375.940 322.850 376.000 ;
        RECT 317.930 375.800 322.850 375.940 ;
        RECT 317.930 375.740 318.250 375.800 ;
        RECT 322.530 375.740 322.850 375.800 ;
        RECT 317.930 17.920 318.250 17.980 ;
        RECT 317.930 17.780 318.620 17.920 ;
        RECT 317.930 17.720 318.250 17.780 ;
        RECT 318.480 17.240 318.620 17.780 ;
        RECT 410.390 17.240 410.710 17.300 ;
        RECT 318.480 17.100 410.710 17.240 ;
        RECT 410.390 17.040 410.710 17.100 ;
      LAYER via ;
        RECT 317.960 375.740 318.220 376.000 ;
        RECT 322.560 375.740 322.820 376.000 ;
        RECT 317.960 17.720 318.220 17.980 ;
        RECT 410.420 17.040 410.680 17.300 ;
      LAYER met2 ;
        RECT 323.370 400.250 323.650 404.000 ;
        RECT 322.620 400.110 323.650 400.250 ;
        RECT 322.620 376.030 322.760 400.110 ;
        RECT 323.370 400.000 323.650 400.110 ;
        RECT 317.960 375.710 318.220 376.030 ;
        RECT 322.560 375.710 322.820 376.030 ;
        RECT 318.020 18.010 318.160 375.710 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 410.420 17.010 410.680 17.330 ;
        RECT 410.480 2.400 410.620 17.010 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 69.070 390.560 69.390 390.620 ;
        RECT 221.790 390.560 222.110 390.620 ;
        RECT 69.070 390.420 222.110 390.560 ;
        RECT 69.070 390.360 69.390 390.420 ;
        RECT 221.790 390.360 222.110 390.420 ;
      LAYER via ;
        RECT 69.100 390.360 69.360 390.620 ;
        RECT 221.820 390.360 222.080 390.620 ;
      LAYER met2 ;
        RECT 221.710 400.180 221.990 404.000 ;
        RECT 221.710 400.000 222.020 400.180 ;
        RECT 221.880 390.650 222.020 400.000 ;
        RECT 69.100 390.330 69.360 390.650 ;
        RECT 221.820 390.330 222.080 390.650 ;
        RECT 69.160 82.870 69.300 390.330 ;
        RECT 69.160 82.730 71.600 82.870 ;
        RECT 71.460 1.770 71.600 82.730 ;
        RECT 73.550 1.770 74.110 2.400 ;
        RECT 71.460 1.630 74.110 1.770 ;
        RECT 73.550 -4.800 74.110 1.630 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 376.280 324.690 376.340 ;
        RECT 327.590 376.280 327.910 376.340 ;
        RECT 324.370 376.140 327.910 376.280 ;
        RECT 324.370 376.080 324.690 376.140 ;
        RECT 327.590 376.080 327.910 376.140 ;
        RECT 324.370 16.560 324.690 16.620 ;
        RECT 428.330 16.560 428.650 16.620 ;
        RECT 324.370 16.420 428.650 16.560 ;
        RECT 324.370 16.360 324.690 16.420 ;
        RECT 428.330 16.360 428.650 16.420 ;
      LAYER via ;
        RECT 324.400 376.080 324.660 376.340 ;
        RECT 327.620 376.080 327.880 376.340 ;
        RECT 324.400 16.360 324.660 16.620 ;
        RECT 428.360 16.360 428.620 16.620 ;
      LAYER met2 ;
        RECT 328.890 400.250 329.170 404.000 ;
        RECT 327.680 400.110 329.170 400.250 ;
        RECT 327.680 376.370 327.820 400.110 ;
        RECT 328.890 400.000 329.170 400.110 ;
        RECT 324.400 376.050 324.660 376.370 ;
        RECT 327.620 376.050 327.880 376.370 ;
        RECT 324.460 16.650 324.600 376.050 ;
        RECT 324.400 16.330 324.660 16.650 ;
        RECT 428.360 16.330 428.620 16.650 ;
        RECT 428.420 2.400 428.560 16.330 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 376.280 331.590 376.340 ;
        RECT 333.110 376.280 333.430 376.340 ;
        RECT 331.270 376.140 333.430 376.280 ;
        RECT 331.270 376.080 331.590 376.140 ;
        RECT 333.110 376.080 333.430 376.140 ;
        RECT 331.270 20.640 331.590 20.700 ;
        RECT 445.810 20.640 446.130 20.700 ;
        RECT 331.270 20.500 446.130 20.640 ;
        RECT 331.270 20.440 331.590 20.500 ;
        RECT 445.810 20.440 446.130 20.500 ;
      LAYER via ;
        RECT 331.300 376.080 331.560 376.340 ;
        RECT 333.140 376.080 333.400 376.340 ;
        RECT 331.300 20.440 331.560 20.700 ;
        RECT 445.840 20.440 446.100 20.700 ;
      LAYER met2 ;
        RECT 334.410 400.250 334.690 404.000 ;
        RECT 333.200 400.110 334.690 400.250 ;
        RECT 333.200 376.370 333.340 400.110 ;
        RECT 334.410 400.000 334.690 400.110 ;
        RECT 331.300 376.050 331.560 376.370 ;
        RECT 333.140 376.050 333.400 376.370 ;
        RECT 331.360 20.730 331.500 376.050 ;
        RECT 331.300 20.410 331.560 20.730 ;
        RECT 445.840 20.410 446.100 20.730 ;
        RECT 445.900 2.400 446.040 20.410 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 339.550 387.160 339.870 387.220 ;
        RECT 389.690 387.160 390.010 387.220 ;
        RECT 339.550 387.020 390.010 387.160 ;
        RECT 339.550 386.960 339.870 387.020 ;
        RECT 389.690 386.960 390.010 387.020 ;
        RECT 389.690 14.860 390.010 14.920 ;
        RECT 463.750 14.860 464.070 14.920 ;
        RECT 389.690 14.720 464.070 14.860 ;
        RECT 389.690 14.660 390.010 14.720 ;
        RECT 463.750 14.660 464.070 14.720 ;
      LAYER via ;
        RECT 339.580 386.960 339.840 387.220 ;
        RECT 389.720 386.960 389.980 387.220 ;
        RECT 389.720 14.660 389.980 14.920 ;
        RECT 463.780 14.660 464.040 14.920 ;
      LAYER met2 ;
        RECT 339.470 400.180 339.750 404.000 ;
        RECT 339.470 400.000 339.780 400.180 ;
        RECT 339.640 387.250 339.780 400.000 ;
        RECT 339.580 386.930 339.840 387.250 ;
        RECT 389.720 386.930 389.980 387.250 ;
        RECT 389.780 14.950 389.920 386.930 ;
        RECT 389.720 14.630 389.980 14.950 ;
        RECT 463.780 14.630 464.040 14.950 ;
        RECT 463.840 2.400 463.980 14.630 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 472.950 389.880 473.270 389.940 ;
        RECT 400.130 389.740 473.270 389.880 ;
        RECT 400.130 389.200 400.270 389.740 ;
        RECT 472.950 389.680 473.270 389.740 ;
        RECT 376.440 389.060 400.270 389.200 ;
        RECT 345.070 388.860 345.390 388.920 ;
        RECT 376.440 388.860 376.580 389.060 ;
        RECT 345.070 388.720 376.580 388.860 ;
        RECT 345.070 388.660 345.390 388.720 ;
        RECT 472.950 16.900 473.270 16.960 ;
        RECT 481.230 16.900 481.550 16.960 ;
        RECT 472.950 16.760 481.550 16.900 ;
        RECT 472.950 16.700 473.270 16.760 ;
        RECT 481.230 16.700 481.550 16.760 ;
      LAYER via ;
        RECT 472.980 389.680 473.240 389.940 ;
        RECT 345.100 388.660 345.360 388.920 ;
        RECT 472.980 16.700 473.240 16.960 ;
        RECT 481.260 16.700 481.520 16.960 ;
      LAYER met2 ;
        RECT 344.990 400.180 345.270 404.000 ;
        RECT 344.990 400.000 345.300 400.180 ;
        RECT 345.160 388.950 345.300 400.000 ;
        RECT 472.980 389.650 473.240 389.970 ;
        RECT 345.100 388.630 345.360 388.950 ;
        RECT 473.040 16.990 473.180 389.650 ;
        RECT 472.980 16.670 473.240 16.990 ;
        RECT 481.260 16.670 481.520 16.990 ;
        RECT 481.320 2.400 481.460 16.670 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 350.590 390.900 350.910 390.960 ;
        RECT 479.850 390.900 480.170 390.960 ;
        RECT 350.590 390.760 480.170 390.900 ;
        RECT 350.590 390.700 350.910 390.760 ;
        RECT 479.850 390.700 480.170 390.760 ;
        RECT 479.390 16.560 479.710 16.620 ;
        RECT 499.170 16.560 499.490 16.620 ;
        RECT 479.390 16.420 499.490 16.560 ;
        RECT 479.390 16.360 479.710 16.420 ;
        RECT 499.170 16.360 499.490 16.420 ;
      LAYER via ;
        RECT 350.620 390.700 350.880 390.960 ;
        RECT 479.880 390.700 480.140 390.960 ;
        RECT 479.420 16.360 479.680 16.620 ;
        RECT 499.200 16.360 499.460 16.620 ;
      LAYER met2 ;
        RECT 350.510 400.180 350.790 404.000 ;
        RECT 350.510 400.000 350.820 400.180 ;
        RECT 350.680 390.990 350.820 400.000 ;
        RECT 350.620 390.670 350.880 390.990 ;
        RECT 479.880 390.670 480.140 390.990 ;
        RECT 479.940 324.370 480.080 390.670 ;
        RECT 479.480 324.230 480.080 324.370 ;
        RECT 479.480 16.650 479.620 324.230 ;
        RECT 479.420 16.330 479.680 16.650 ;
        RECT 499.200 16.330 499.460 16.650 ;
        RECT 499.260 2.400 499.400 16.330 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 354.270 390.220 354.590 390.280 ;
        RECT 500.550 390.220 500.870 390.280 ;
        RECT 354.270 390.080 500.870 390.220 ;
        RECT 354.270 390.020 354.590 390.080 ;
        RECT 500.550 390.020 500.870 390.080 ;
        RECT 500.550 15.540 500.870 15.600 ;
        RECT 516.650 15.540 516.970 15.600 ;
        RECT 500.550 15.400 516.970 15.540 ;
        RECT 500.550 15.340 500.870 15.400 ;
        RECT 516.650 15.340 516.970 15.400 ;
      LAYER via ;
        RECT 354.300 390.020 354.560 390.280 ;
        RECT 500.580 390.020 500.840 390.280 ;
        RECT 500.580 15.340 500.840 15.600 ;
        RECT 516.680 15.340 516.940 15.600 ;
      LAYER met2 ;
        RECT 355.570 400.250 355.850 404.000 ;
        RECT 354.360 400.110 355.850 400.250 ;
        RECT 354.360 390.310 354.500 400.110 ;
        RECT 355.570 400.000 355.850 400.110 ;
        RECT 354.300 389.990 354.560 390.310 ;
        RECT 500.580 389.990 500.840 390.310 ;
        RECT 500.640 15.630 500.780 389.990 ;
        RECT 500.580 15.310 500.840 15.630 ;
        RECT 516.680 15.310 516.940 15.630 ;
        RECT 516.740 2.400 516.880 15.310 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 19.280 359.190 19.340 ;
        RECT 534.590 19.280 534.910 19.340 ;
        RECT 358.870 19.140 534.910 19.280 ;
        RECT 358.870 19.080 359.190 19.140 ;
        RECT 534.590 19.080 534.910 19.140 ;
      LAYER via ;
        RECT 358.900 19.080 359.160 19.340 ;
        RECT 534.620 19.080 534.880 19.340 ;
      LAYER met2 ;
        RECT 361.090 400.250 361.370 404.000 ;
        RECT 359.880 400.110 361.370 400.250 ;
        RECT 359.880 351.970 360.020 400.110 ;
        RECT 361.090 400.000 361.370 400.110 ;
        RECT 358.960 351.830 360.020 351.970 ;
        RECT 358.960 19.370 359.100 351.830 ;
        RECT 358.900 19.050 359.160 19.370 ;
        RECT 534.620 19.050 534.880 19.370 ;
        RECT 534.680 2.400 534.820 19.050 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.990 390.900 507.310 390.960 ;
        RECT 488.220 390.760 507.310 390.900 ;
        RECT 366.690 390.560 367.010 390.620 ;
        RECT 488.220 390.560 488.360 390.760 ;
        RECT 506.990 390.700 507.310 390.760 ;
        RECT 366.690 390.420 488.360 390.560 ;
        RECT 366.690 390.360 367.010 390.420 ;
        RECT 506.990 16.560 507.310 16.620 ;
        RECT 552.530 16.560 552.850 16.620 ;
        RECT 506.990 16.420 552.850 16.560 ;
        RECT 506.990 16.360 507.310 16.420 ;
        RECT 552.530 16.360 552.850 16.420 ;
      LAYER via ;
        RECT 366.720 390.360 366.980 390.620 ;
        RECT 507.020 390.700 507.280 390.960 ;
        RECT 507.020 16.360 507.280 16.620 ;
        RECT 552.560 16.360 552.820 16.620 ;
      LAYER met2 ;
        RECT 366.610 400.180 366.890 404.000 ;
        RECT 366.610 400.000 366.920 400.180 ;
        RECT 366.780 390.650 366.920 400.000 ;
        RECT 507.020 390.670 507.280 390.990 ;
        RECT 366.720 390.330 366.980 390.650 ;
        RECT 507.080 16.650 507.220 390.670 ;
        RECT 507.020 16.330 507.280 16.650 ;
        RECT 552.560 16.330 552.820 16.650 ;
        RECT 552.620 2.400 552.760 16.330 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.230 22.340 366.550 22.400 ;
        RECT 510.670 22.340 510.990 22.400 ;
        RECT 366.230 22.200 510.990 22.340 ;
        RECT 366.230 22.140 366.550 22.200 ;
        RECT 510.670 22.140 510.990 22.200 ;
        RECT 510.670 19.960 510.990 20.020 ;
        RECT 570.010 19.960 570.330 20.020 ;
        RECT 510.670 19.820 570.330 19.960 ;
        RECT 510.670 19.760 510.990 19.820 ;
        RECT 570.010 19.760 570.330 19.820 ;
      LAYER via ;
        RECT 366.260 22.140 366.520 22.400 ;
        RECT 510.700 22.140 510.960 22.400 ;
        RECT 510.700 19.760 510.960 20.020 ;
        RECT 570.040 19.760 570.300 20.020 ;
      LAYER met2 ;
        RECT 371.670 400.250 371.950 404.000 ;
        RECT 370.460 400.110 371.950 400.250 ;
        RECT 370.460 324.370 370.600 400.110 ;
        RECT 371.670 400.000 371.950 400.110 ;
        RECT 366.320 324.230 370.600 324.370 ;
        RECT 366.320 22.430 366.460 324.230 ;
        RECT 366.260 22.110 366.520 22.430 ;
        RECT 510.700 22.110 510.960 22.430 ;
        RECT 510.760 20.050 510.900 22.110 ;
        RECT 510.700 19.730 510.960 20.050 ;
        RECT 570.040 19.730 570.300 20.050 ;
        RECT 570.100 2.400 570.240 19.730 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.490 19.280 541.810 19.340 ;
        RECT 587.950 19.280 588.270 19.340 ;
        RECT 541.490 19.140 588.270 19.280 ;
        RECT 541.490 19.080 541.810 19.140 ;
        RECT 587.950 19.080 588.270 19.140 ;
      LAYER via ;
        RECT 541.520 19.080 541.780 19.340 ;
        RECT 587.980 19.080 588.240 19.340 ;
      LAYER met2 ;
        RECT 377.190 400.180 377.470 404.000 ;
        RECT 377.190 400.000 377.500 400.180 ;
        RECT 377.360 389.485 377.500 400.000 ;
        RECT 377.290 389.115 377.570 389.485 ;
        RECT 541.510 389.115 541.790 389.485 ;
        RECT 541.580 19.370 541.720 389.115 ;
        RECT 541.520 19.050 541.780 19.370 ;
        RECT 587.980 19.050 588.240 19.370 ;
        RECT 588.040 2.400 588.180 19.050 ;
        RECT 587.830 -4.800 588.390 2.400 ;
      LAYER via2 ;
        RECT 377.290 389.160 377.570 389.440 ;
        RECT 541.510 389.160 541.790 389.440 ;
      LAYER met3 ;
        RECT 377.265 389.450 377.595 389.465 ;
        RECT 541.485 389.450 541.815 389.465 ;
        RECT 377.265 389.150 541.815 389.450 ;
        RECT 377.265 389.135 377.595 389.150 ;
        RECT 541.485 389.135 541.815 389.150 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 97.130 20.300 97.450 20.360 ;
        RECT 97.130 20.160 203.160 20.300 ;
        RECT 97.130 20.100 97.450 20.160 ;
        RECT 203.020 19.280 203.160 20.160 ;
        RECT 229.150 19.280 229.470 19.340 ;
        RECT 203.020 19.140 229.470 19.280 ;
        RECT 229.150 19.080 229.470 19.140 ;
      LAYER via ;
        RECT 97.160 20.100 97.420 20.360 ;
        RECT 229.180 19.080 229.440 19.340 ;
      LAYER met2 ;
        RECT 229.070 400.250 229.350 404.000 ;
        RECT 229.070 400.110 230.300 400.250 ;
        RECT 229.070 400.000 229.350 400.110 ;
        RECT 230.160 303.670 230.300 400.110 ;
        RECT 229.240 303.530 230.300 303.670 ;
        RECT 97.160 20.070 97.420 20.390 ;
        RECT 97.220 2.400 97.360 20.070 ;
        RECT 229.240 19.370 229.380 303.530 ;
        RECT 229.180 19.050 229.440 19.370 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.490 19.620 380.810 19.680 ;
        RECT 605.430 19.620 605.750 19.680 ;
        RECT 380.490 19.480 605.750 19.620 ;
        RECT 380.490 19.420 380.810 19.480 ;
        RECT 605.430 19.420 605.750 19.480 ;
      LAYER via ;
        RECT 380.520 19.420 380.780 19.680 ;
        RECT 605.460 19.420 605.720 19.680 ;
      LAYER met2 ;
        RECT 382.710 400.250 382.990 404.000 ;
        RECT 381.500 400.110 382.990 400.250 ;
        RECT 381.500 351.970 381.640 400.110 ;
        RECT 382.710 400.000 382.990 400.110 ;
        RECT 380.580 351.830 381.640 351.970 ;
        RECT 380.580 19.710 380.720 351.830 ;
        RECT 380.520 19.390 380.780 19.710 ;
        RECT 605.460 19.390 605.720 19.710 ;
        RECT 605.520 2.400 605.660 19.390 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 444.890 392.600 445.210 392.660 ;
        RECT 548.390 392.600 548.710 392.660 ;
        RECT 444.890 392.460 548.710 392.600 ;
        RECT 444.890 392.400 445.210 392.460 ;
        RECT 548.390 392.400 548.710 392.460 ;
        RECT 444.890 388.520 445.210 388.580 ;
        RECT 391.620 388.380 445.210 388.520 ;
        RECT 387.850 388.180 388.170 388.240 ;
        RECT 391.620 388.180 391.760 388.380 ;
        RECT 444.890 388.320 445.210 388.380 ;
        RECT 387.850 388.040 391.760 388.180 ;
        RECT 387.850 387.980 388.170 388.040 ;
        RECT 548.390 20.640 548.710 20.700 ;
        RECT 623.370 20.640 623.690 20.700 ;
        RECT 548.390 20.500 623.690 20.640 ;
        RECT 548.390 20.440 548.710 20.500 ;
        RECT 623.370 20.440 623.690 20.500 ;
      LAYER via ;
        RECT 444.920 392.400 445.180 392.660 ;
        RECT 548.420 392.400 548.680 392.660 ;
        RECT 387.880 387.980 388.140 388.240 ;
        RECT 444.920 388.320 445.180 388.580 ;
        RECT 548.420 20.440 548.680 20.700 ;
        RECT 623.400 20.440 623.660 20.700 ;
      LAYER met2 ;
        RECT 387.770 400.180 388.050 404.000 ;
        RECT 387.770 400.000 388.080 400.180 ;
        RECT 387.940 388.270 388.080 400.000 ;
        RECT 444.920 392.370 445.180 392.690 ;
        RECT 548.420 392.370 548.680 392.690 ;
        RECT 444.980 388.610 445.120 392.370 ;
        RECT 444.920 388.290 445.180 388.610 ;
        RECT 387.880 387.950 388.140 388.270 ;
        RECT 548.480 20.730 548.620 392.370 ;
        RECT 548.420 20.410 548.680 20.730 ;
        RECT 623.400 20.410 623.660 20.730 ;
        RECT 623.460 2.400 623.600 20.410 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 117.370 391.580 117.690 391.640 ;
        RECT 236.050 391.580 236.370 391.640 ;
        RECT 117.370 391.440 236.370 391.580 ;
        RECT 117.370 391.380 117.690 391.440 ;
        RECT 236.050 391.380 236.370 391.440 ;
      LAYER via ;
        RECT 117.400 391.380 117.660 391.640 ;
        RECT 236.080 391.380 236.340 391.640 ;
      LAYER met2 ;
        RECT 235.970 400.180 236.250 404.000 ;
        RECT 235.970 400.000 236.280 400.180 ;
        RECT 236.140 391.670 236.280 400.000 ;
        RECT 117.400 391.350 117.660 391.670 ;
        RECT 236.080 391.350 236.340 391.670 ;
        RECT 117.460 82.870 117.600 391.350 ;
        RECT 117.460 82.730 121.280 82.870 ;
        RECT 121.140 2.400 121.280 82.730 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.030 376.280 242.350 376.340 ;
        RECT 243.410 376.280 243.730 376.340 ;
        RECT 242.030 376.140 243.730 376.280 ;
        RECT 242.030 376.080 242.350 376.140 ;
        RECT 243.410 376.080 243.730 376.140 ;
        RECT 144.510 16.560 144.830 16.620 ;
        RECT 242.030 16.560 242.350 16.620 ;
        RECT 144.510 16.420 242.350 16.560 ;
        RECT 144.510 16.360 144.830 16.420 ;
        RECT 242.030 16.360 242.350 16.420 ;
      LAYER via ;
        RECT 242.060 376.080 242.320 376.340 ;
        RECT 243.440 376.080 243.700 376.340 ;
        RECT 144.540 16.360 144.800 16.620 ;
        RECT 242.060 16.360 242.320 16.620 ;
      LAYER met2 ;
        RECT 243.330 400.180 243.610 404.000 ;
        RECT 243.330 400.000 243.640 400.180 ;
        RECT 243.500 376.370 243.640 400.000 ;
        RECT 242.060 376.050 242.320 376.370 ;
        RECT 243.440 376.050 243.700 376.370 ;
        RECT 242.120 16.650 242.260 376.050 ;
        RECT 144.540 16.330 144.800 16.650 ;
        RECT 242.060 16.330 242.320 16.650 ;
        RECT 144.600 2.400 144.740 16.330 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.770 392.600 159.090 392.660 ;
        RECT 248.470 392.600 248.790 392.660 ;
        RECT 158.770 392.460 248.790 392.600 ;
        RECT 158.770 392.400 159.090 392.460 ;
        RECT 248.470 392.400 248.790 392.460 ;
      LAYER via ;
        RECT 158.800 392.400 159.060 392.660 ;
        RECT 248.500 392.400 248.760 392.660 ;
      LAYER met2 ;
        RECT 248.390 400.180 248.670 404.000 ;
        RECT 248.390 400.000 248.700 400.180 ;
        RECT 248.560 392.690 248.700 400.000 ;
        RECT 158.800 392.370 159.060 392.690 ;
        RECT 248.500 392.370 248.760 392.690 ;
        RECT 158.860 82.870 159.000 392.370 ;
        RECT 158.860 82.730 159.920 82.870 ;
        RECT 159.780 1.770 159.920 82.730 ;
        RECT 161.870 1.770 162.430 2.400 ;
        RECT 159.780 1.630 162.430 1.770 ;
        RECT 161.870 -4.800 162.430 1.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.930 376.280 249.250 376.340 ;
        RECT 252.610 376.280 252.930 376.340 ;
        RECT 248.930 376.140 252.930 376.280 ;
        RECT 248.930 376.080 249.250 376.140 ;
        RECT 252.610 376.080 252.930 376.140 ;
        RECT 179.930 15.540 180.250 15.600 ;
        RECT 248.930 15.540 249.250 15.600 ;
        RECT 179.930 15.400 249.250 15.540 ;
        RECT 179.930 15.340 180.250 15.400 ;
        RECT 248.930 15.340 249.250 15.400 ;
      LAYER via ;
        RECT 248.960 376.080 249.220 376.340 ;
        RECT 252.640 376.080 252.900 376.340 ;
        RECT 179.960 15.340 180.220 15.600 ;
        RECT 248.960 15.340 249.220 15.600 ;
      LAYER met2 ;
        RECT 253.910 400.250 254.190 404.000 ;
        RECT 252.700 400.110 254.190 400.250 ;
        RECT 252.700 376.370 252.840 400.110 ;
        RECT 253.910 400.000 254.190 400.110 ;
        RECT 248.960 376.050 249.220 376.370 ;
        RECT 252.640 376.050 252.900 376.370 ;
        RECT 249.020 15.630 249.160 376.050 ;
        RECT 179.960 15.310 180.220 15.630 ;
        RECT 248.960 15.310 249.220 15.630 ;
        RECT 180.020 2.400 180.160 15.310 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 193.270 388.860 193.590 388.920 ;
        RECT 259.510 388.860 259.830 388.920 ;
        RECT 193.270 388.720 259.830 388.860 ;
        RECT 193.270 388.660 193.590 388.720 ;
        RECT 259.510 388.660 259.830 388.720 ;
      LAYER via ;
        RECT 193.300 388.660 193.560 388.920 ;
        RECT 259.540 388.660 259.800 388.920 ;
      LAYER met2 ;
        RECT 259.430 400.180 259.710 404.000 ;
        RECT 259.430 400.000 259.740 400.180 ;
        RECT 259.600 388.950 259.740 400.000 ;
        RECT 193.300 388.630 193.560 388.950 ;
        RECT 259.540 388.630 259.800 388.950 ;
        RECT 193.360 82.870 193.500 388.630 ;
        RECT 193.360 82.730 195.800 82.870 ;
        RECT 195.660 1.770 195.800 82.730 ;
        RECT 197.750 1.770 198.310 2.400 ;
        RECT 195.660 1.630 198.310 1.770 ;
        RECT 197.750 -4.800 198.310 1.630 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 224.090 389.200 224.410 389.260 ;
        RECT 264.570 389.200 264.890 389.260 ;
        RECT 224.090 389.060 264.890 389.200 ;
        RECT 224.090 389.000 224.410 389.060 ;
        RECT 264.570 389.000 264.890 389.060 ;
        RECT 215.350 17.580 215.670 17.640 ;
        RECT 224.090 17.580 224.410 17.640 ;
        RECT 215.350 17.440 224.410 17.580 ;
        RECT 215.350 17.380 215.670 17.440 ;
        RECT 224.090 17.380 224.410 17.440 ;
      LAYER via ;
        RECT 224.120 389.000 224.380 389.260 ;
        RECT 264.600 389.000 264.860 389.260 ;
        RECT 215.380 17.380 215.640 17.640 ;
        RECT 224.120 17.380 224.380 17.640 ;
      LAYER met2 ;
        RECT 264.490 400.180 264.770 404.000 ;
        RECT 264.490 400.000 264.800 400.180 ;
        RECT 264.660 389.290 264.800 400.000 ;
        RECT 224.120 388.970 224.380 389.290 ;
        RECT 264.600 388.970 264.860 389.290 ;
        RECT 224.180 17.670 224.320 388.970 ;
        RECT 215.380 17.350 215.640 17.670 ;
        RECT 224.120 17.350 224.380 17.670 ;
        RECT 215.440 2.400 215.580 17.350 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 251.690 386.820 252.010 386.880 ;
        RECT 270.090 386.820 270.410 386.880 ;
        RECT 251.690 386.680 270.410 386.820 ;
        RECT 251.690 386.620 252.010 386.680 ;
        RECT 270.090 386.620 270.410 386.680 ;
        RECT 233.290 16.220 233.610 16.280 ;
        RECT 251.690 16.220 252.010 16.280 ;
        RECT 233.290 16.080 252.010 16.220 ;
        RECT 233.290 16.020 233.610 16.080 ;
        RECT 251.690 16.020 252.010 16.080 ;
      LAYER via ;
        RECT 251.720 386.620 251.980 386.880 ;
        RECT 270.120 386.620 270.380 386.880 ;
        RECT 233.320 16.020 233.580 16.280 ;
        RECT 251.720 16.020 251.980 16.280 ;
      LAYER met2 ;
        RECT 270.010 400.180 270.290 404.000 ;
        RECT 270.010 400.000 270.320 400.180 ;
        RECT 270.180 386.910 270.320 400.000 ;
        RECT 251.720 386.590 251.980 386.910 ;
        RECT 270.120 386.590 270.380 386.910 ;
        RECT 251.780 16.310 251.920 386.590 ;
        RECT 233.320 15.990 233.580 16.310 ;
        RECT 251.720 15.990 251.980 16.310 ;
        RECT 233.380 2.400 233.520 15.990 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 214.430 376.280 214.750 376.340 ;
        RECT 215.810 376.280 216.130 376.340 ;
        RECT 214.430 376.140 216.130 376.280 ;
        RECT 214.430 376.080 214.750 376.140 ;
        RECT 215.810 376.080 216.130 376.140 ;
        RECT 55.730 18.940 56.050 19.000 ;
        RECT 55.730 18.800 196.720 18.940 ;
        RECT 55.730 18.740 56.050 18.800 ;
        RECT 196.580 18.600 196.720 18.800 ;
        RECT 214.430 18.600 214.750 18.660 ;
        RECT 196.580 18.460 214.750 18.600 ;
        RECT 214.430 18.400 214.750 18.460 ;
      LAYER via ;
        RECT 214.460 376.080 214.720 376.340 ;
        RECT 215.840 376.080 216.100 376.340 ;
        RECT 55.760 18.740 56.020 19.000 ;
        RECT 214.460 18.400 214.720 18.660 ;
      LAYER met2 ;
        RECT 216.190 400.250 216.470 404.000 ;
        RECT 215.900 400.110 216.470 400.250 ;
        RECT 215.900 376.370 216.040 400.110 ;
        RECT 216.190 400.000 216.470 400.110 ;
        RECT 214.460 376.050 214.720 376.370 ;
        RECT 215.840 376.050 216.100 376.370 ;
        RECT 55.760 18.710 56.020 19.030 ;
        RECT 55.820 2.400 55.960 18.710 ;
        RECT 214.520 18.690 214.660 376.050 ;
        RECT 214.460 18.370 214.720 18.690 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 75.970 391.240 76.290 391.300 ;
        RECT 222.250 391.240 222.570 391.300 ;
        RECT 75.970 391.100 222.570 391.240 ;
        RECT 75.970 391.040 76.290 391.100 ;
        RECT 222.250 391.040 222.570 391.100 ;
      LAYER via ;
        RECT 76.000 391.040 76.260 391.300 ;
        RECT 222.280 391.040 222.540 391.300 ;
      LAYER met2 ;
        RECT 223.550 400.250 223.830 404.000 ;
        RECT 222.340 400.110 223.830 400.250 ;
        RECT 222.340 391.330 222.480 400.110 ;
        RECT 223.550 400.000 223.830 400.110 ;
        RECT 76.000 391.010 76.260 391.330 ;
        RECT 222.280 391.010 222.540 391.330 ;
        RECT 76.060 82.870 76.200 391.010 ;
        RECT 76.060 82.730 79.880 82.870 ;
        RECT 79.740 2.400 79.880 82.730 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.230 376.280 228.550 376.340 ;
        RECT 230.530 376.280 230.850 376.340 ;
        RECT 228.230 376.140 230.850 376.280 ;
        RECT 228.230 376.080 228.550 376.140 ;
        RECT 230.530 376.080 230.850 376.140 ;
        RECT 103.110 20.640 103.430 20.700 ;
        RECT 103.110 20.500 203.620 20.640 ;
        RECT 103.110 20.440 103.430 20.500 ;
        RECT 203.480 19.620 203.620 20.500 ;
        RECT 228.230 19.620 228.550 19.680 ;
        RECT 203.480 19.480 228.550 19.620 ;
        RECT 228.230 19.420 228.550 19.480 ;
      LAYER via ;
        RECT 228.260 376.080 228.520 376.340 ;
        RECT 230.560 376.080 230.820 376.340 ;
        RECT 103.140 20.440 103.400 20.700 ;
        RECT 228.260 19.420 228.520 19.680 ;
      LAYER met2 ;
        RECT 230.910 400.250 231.190 404.000 ;
        RECT 230.620 400.110 231.190 400.250 ;
        RECT 230.620 376.370 230.760 400.110 ;
        RECT 230.910 400.000 231.190 400.110 ;
        RECT 228.260 376.050 228.520 376.370 ;
        RECT 230.560 376.050 230.820 376.370 ;
        RECT 103.140 20.410 103.400 20.730 ;
        RECT 103.200 2.400 103.340 20.410 ;
        RECT 228.320 19.710 228.460 376.050 ;
        RECT 228.260 19.390 228.520 19.710 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.270 392.260 124.590 392.320 ;
        RECT 237.890 392.260 238.210 392.320 ;
        RECT 124.270 392.120 238.210 392.260 ;
        RECT 124.270 392.060 124.590 392.120 ;
        RECT 237.890 392.060 238.210 392.120 ;
      LAYER via ;
        RECT 124.300 392.060 124.560 392.320 ;
        RECT 237.920 392.060 238.180 392.320 ;
      LAYER met2 ;
        RECT 237.810 400.180 238.090 404.000 ;
        RECT 237.810 400.000 238.120 400.180 ;
        RECT 237.980 392.350 238.120 400.000 ;
        RECT 124.300 392.030 124.560 392.350 ;
        RECT 237.920 392.030 238.180 392.350 ;
        RECT 124.360 82.870 124.500 392.030 ;
        RECT 124.360 82.730 126.800 82.870 ;
        RECT 126.660 2.400 126.800 82.730 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 207.990 17.240 208.310 17.300 ;
        RECT 26.290 17.100 208.310 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 207.990 17.040 208.310 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 208.020 17.040 208.280 17.300 ;
      LAYER met2 ;
        RECT 207.450 400.250 207.730 404.000 ;
        RECT 207.450 400.110 208.220 400.250 ;
        RECT 207.450 400.000 207.730 400.110 ;
        RECT 208.080 17.330 208.220 400.110 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 208.020 17.010 208.280 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.670 390.220 27.990 390.280 ;
        RECT 209.370 390.220 209.690 390.280 ;
        RECT 27.670 390.080 209.690 390.220 ;
        RECT 27.670 390.020 27.990 390.080 ;
        RECT 209.370 390.020 209.690 390.080 ;
      LAYER via ;
        RECT 27.700 390.020 27.960 390.280 ;
        RECT 209.400 390.020 209.660 390.280 ;
      LAYER met2 ;
        RECT 209.290 400.180 209.570 404.000 ;
        RECT 209.290 400.000 209.600 400.180 ;
        RECT 209.460 390.310 209.600 400.000 ;
        RECT 27.700 389.990 27.960 390.310 ;
        RECT 209.400 389.990 209.660 390.310 ;
        RECT 27.760 82.870 27.900 389.990 ;
        RECT 27.760 82.730 30.200 82.870 ;
        RECT 30.060 1.770 30.200 82.730 ;
        RECT 32.150 1.770 32.710 2.400 ;
        RECT 30.060 1.630 32.710 1.770 ;
        RECT 32.150 -4.800 32.710 1.630 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 205.520 410.795 1094.240 987.605 ;
      LAYER met1 ;
        RECT 203.750 410.640 1094.240 990.880 ;
      LAYER met2 ;
        RECT 204.330 995.720 210.850 996.770 ;
        RECT 211.690 995.720 218.210 996.770 ;
        RECT 219.050 995.720 225.570 996.770 ;
        RECT 226.410 995.720 232.930 996.770 ;
        RECT 233.770 995.720 240.290 996.770 ;
        RECT 241.130 995.720 247.650 996.770 ;
        RECT 248.490 995.720 255.010 996.770 ;
        RECT 255.850 995.720 262.370 996.770 ;
        RECT 263.210 995.720 269.730 996.770 ;
        RECT 270.570 995.720 277.090 996.770 ;
        RECT 277.930 995.720 284.450 996.770 ;
        RECT 285.290 995.720 291.810 996.770 ;
        RECT 292.650 995.720 299.170 996.770 ;
        RECT 300.010 995.720 306.530 996.770 ;
        RECT 307.370 995.720 313.890 996.770 ;
        RECT 314.730 995.720 321.250 996.770 ;
        RECT 322.090 995.720 328.610 996.770 ;
        RECT 329.450 995.720 335.970 996.770 ;
        RECT 336.810 995.720 343.330 996.770 ;
        RECT 344.170 995.720 350.690 996.770 ;
        RECT 351.530 995.720 358.050 996.770 ;
        RECT 358.890 995.720 365.410 996.770 ;
        RECT 366.250 995.720 372.770 996.770 ;
        RECT 373.610 995.720 380.130 996.770 ;
        RECT 380.970 995.720 387.950 996.770 ;
        RECT 388.790 995.720 395.310 996.770 ;
        RECT 396.150 995.720 402.670 996.770 ;
        RECT 403.510 995.720 410.030 996.770 ;
        RECT 410.870 995.720 417.390 996.770 ;
        RECT 418.230 995.720 424.750 996.770 ;
        RECT 425.590 995.720 432.110 996.770 ;
        RECT 432.950 995.720 439.470 996.770 ;
        RECT 440.310 995.720 446.830 996.770 ;
        RECT 447.670 995.720 454.190 996.770 ;
        RECT 455.030 995.720 461.550 996.770 ;
        RECT 462.390 995.720 468.910 996.770 ;
        RECT 469.750 995.720 476.270 996.770 ;
        RECT 477.110 995.720 483.630 996.770 ;
        RECT 484.470 995.720 490.990 996.770 ;
        RECT 491.830 995.720 498.350 996.770 ;
        RECT 499.190 995.720 505.710 996.770 ;
        RECT 506.550 995.720 513.070 996.770 ;
        RECT 513.910 995.720 520.430 996.770 ;
        RECT 521.270 995.720 527.790 996.770 ;
        RECT 528.630 995.720 535.150 996.770 ;
        RECT 535.990 995.720 542.510 996.770 ;
        RECT 543.350 995.720 549.870 996.770 ;
        RECT 550.710 995.720 557.230 996.770 ;
        RECT 558.070 995.720 565.050 996.770 ;
        RECT 565.890 995.720 572.410 996.770 ;
        RECT 573.250 995.720 579.770 996.770 ;
        RECT 580.610 995.720 587.130 996.770 ;
        RECT 587.970 995.720 594.490 996.770 ;
        RECT 595.330 995.720 601.850 996.770 ;
        RECT 602.690 995.720 609.210 996.770 ;
        RECT 610.050 995.720 616.570 996.770 ;
        RECT 617.410 995.720 623.930 996.770 ;
        RECT 624.770 995.720 631.290 996.770 ;
        RECT 632.130 995.720 638.650 996.770 ;
        RECT 639.490 995.720 646.010 996.770 ;
        RECT 646.850 995.720 653.370 996.770 ;
        RECT 654.210 995.720 660.730 996.770 ;
        RECT 661.570 995.720 668.090 996.770 ;
        RECT 668.930 995.720 675.450 996.770 ;
        RECT 676.290 995.720 682.810 996.770 ;
        RECT 683.650 995.720 690.170 996.770 ;
        RECT 691.010 995.720 697.530 996.770 ;
        RECT 698.370 995.720 704.890 996.770 ;
        RECT 705.730 995.720 712.250 996.770 ;
        RECT 713.090 995.720 719.610 996.770 ;
        RECT 720.450 995.720 726.970 996.770 ;
        RECT 727.810 995.720 734.330 996.770 ;
        RECT 735.170 995.720 741.690 996.770 ;
        RECT 742.530 995.720 749.510 996.770 ;
        RECT 750.350 995.720 756.870 996.770 ;
        RECT 757.710 995.720 764.230 996.770 ;
        RECT 765.070 995.720 771.590 996.770 ;
        RECT 772.430 995.720 778.950 996.770 ;
        RECT 779.790 995.720 786.310 996.770 ;
        RECT 787.150 995.720 793.670 996.770 ;
        RECT 794.510 995.720 801.030 996.770 ;
        RECT 801.870 995.720 808.390 996.770 ;
        RECT 809.230 995.720 815.750 996.770 ;
        RECT 816.590 995.720 823.110 996.770 ;
        RECT 823.950 995.720 830.470 996.770 ;
        RECT 831.310 995.720 837.830 996.770 ;
        RECT 838.670 995.720 845.190 996.770 ;
        RECT 846.030 995.720 852.550 996.770 ;
        RECT 853.390 995.720 859.910 996.770 ;
        RECT 860.750 995.720 867.270 996.770 ;
        RECT 868.110 995.720 874.630 996.770 ;
        RECT 875.470 995.720 881.990 996.770 ;
        RECT 882.830 995.720 889.350 996.770 ;
        RECT 890.190 995.720 896.710 996.770 ;
        RECT 897.550 995.720 904.070 996.770 ;
        RECT 904.910 995.720 911.430 996.770 ;
        RECT 912.270 995.720 918.790 996.770 ;
        RECT 919.630 995.720 926.610 996.770 ;
        RECT 927.450 995.720 933.970 996.770 ;
        RECT 934.810 995.720 941.330 996.770 ;
        RECT 942.170 995.720 948.690 996.770 ;
        RECT 949.530 995.720 956.050 996.770 ;
        RECT 956.890 995.720 963.410 996.770 ;
        RECT 964.250 995.720 970.770 996.770 ;
        RECT 971.610 995.720 978.130 996.770 ;
        RECT 978.970 995.720 985.490 996.770 ;
        RECT 986.330 995.720 992.850 996.770 ;
        RECT 993.690 995.720 1000.210 996.770 ;
        RECT 1001.050 995.720 1007.570 996.770 ;
        RECT 1008.410 995.720 1014.930 996.770 ;
        RECT 1015.770 995.720 1022.290 996.770 ;
        RECT 1023.130 995.720 1029.650 996.770 ;
        RECT 1030.490 995.720 1037.010 996.770 ;
        RECT 1037.850 995.720 1044.370 996.770 ;
        RECT 1045.210 995.720 1051.730 996.770 ;
        RECT 1052.570 995.720 1059.090 996.770 ;
        RECT 1059.930 995.720 1066.450 996.770 ;
        RECT 1067.290 995.720 1073.810 996.770 ;
        RECT 1074.650 995.720 1081.170 996.770 ;
        RECT 1082.010 995.720 1088.530 996.770 ;
        RECT 1089.370 995.720 1090.930 996.770 ;
        RECT 203.780 404.280 1090.930 995.720 ;
        RECT 204.330 404.000 205.330 404.280 ;
        RECT 206.170 404.000 207.170 404.280 ;
        RECT 208.010 404.000 209.010 404.280 ;
        RECT 209.850 404.000 210.850 404.280 ;
        RECT 211.690 404.000 212.690 404.280 ;
        RECT 213.530 404.000 214.530 404.280 ;
        RECT 215.370 404.000 215.910 404.280 ;
        RECT 216.750 404.000 217.750 404.280 ;
        RECT 218.590 404.000 219.590 404.280 ;
        RECT 220.430 404.000 221.430 404.280 ;
        RECT 222.270 404.000 223.270 404.280 ;
        RECT 224.110 404.000 225.110 404.280 ;
        RECT 225.950 404.000 226.950 404.280 ;
        RECT 227.790 404.000 228.790 404.280 ;
        RECT 229.630 404.000 230.630 404.280 ;
        RECT 231.470 404.000 232.010 404.280 ;
        RECT 232.850 404.000 233.850 404.280 ;
        RECT 234.690 404.000 235.690 404.280 ;
        RECT 236.530 404.000 237.530 404.280 ;
        RECT 238.370 404.000 239.370 404.280 ;
        RECT 240.210 404.000 241.210 404.280 ;
        RECT 242.050 404.000 243.050 404.280 ;
        RECT 243.890 404.000 244.890 404.280 ;
        RECT 245.730 404.000 246.270 404.280 ;
        RECT 247.110 404.000 248.110 404.280 ;
        RECT 248.950 404.000 249.950 404.280 ;
        RECT 250.790 404.000 251.790 404.280 ;
        RECT 252.630 404.000 253.630 404.280 ;
        RECT 254.470 404.000 255.470 404.280 ;
        RECT 256.310 404.000 257.310 404.280 ;
        RECT 258.150 404.000 259.150 404.280 ;
        RECT 259.990 404.000 260.990 404.280 ;
        RECT 261.830 404.000 262.370 404.280 ;
        RECT 263.210 404.000 264.210 404.280 ;
        RECT 265.050 404.000 266.050 404.280 ;
        RECT 266.890 404.000 267.890 404.280 ;
        RECT 268.730 404.000 269.730 404.280 ;
        RECT 270.570 404.000 271.570 404.280 ;
        RECT 272.410 404.000 273.410 404.280 ;
        RECT 274.250 404.000 275.250 404.280 ;
        RECT 276.090 404.000 276.630 404.280 ;
        RECT 277.470 404.000 278.470 404.280 ;
        RECT 279.310 404.000 280.310 404.280 ;
        RECT 281.150 404.000 282.150 404.280 ;
        RECT 282.990 404.000 283.990 404.280 ;
        RECT 284.830 404.000 285.830 404.280 ;
        RECT 286.670 404.000 287.670 404.280 ;
        RECT 288.510 404.000 289.510 404.280 ;
        RECT 290.350 404.000 291.350 404.280 ;
        RECT 292.190 404.000 292.730 404.280 ;
        RECT 293.570 404.000 294.570 404.280 ;
        RECT 295.410 404.000 296.410 404.280 ;
        RECT 297.250 404.000 298.250 404.280 ;
        RECT 299.090 404.000 300.090 404.280 ;
        RECT 300.930 404.000 301.930 404.280 ;
        RECT 302.770 404.000 303.770 404.280 ;
        RECT 304.610 404.000 305.610 404.280 ;
        RECT 306.450 404.000 306.990 404.280 ;
        RECT 307.830 404.000 308.830 404.280 ;
        RECT 309.670 404.000 310.670 404.280 ;
        RECT 311.510 404.000 312.510 404.280 ;
        RECT 313.350 404.000 314.350 404.280 ;
        RECT 315.190 404.000 316.190 404.280 ;
        RECT 317.030 404.000 318.030 404.280 ;
        RECT 318.870 404.000 319.870 404.280 ;
        RECT 320.710 404.000 321.710 404.280 ;
        RECT 322.550 404.000 323.090 404.280 ;
        RECT 323.930 404.000 324.930 404.280 ;
        RECT 325.770 404.000 326.770 404.280 ;
        RECT 327.610 404.000 328.610 404.280 ;
        RECT 329.450 404.000 330.450 404.280 ;
        RECT 331.290 404.000 332.290 404.280 ;
        RECT 333.130 404.000 334.130 404.280 ;
        RECT 334.970 404.000 335.970 404.280 ;
        RECT 336.810 404.000 337.350 404.280 ;
        RECT 338.190 404.000 339.190 404.280 ;
        RECT 340.030 404.000 341.030 404.280 ;
        RECT 341.870 404.000 342.870 404.280 ;
        RECT 343.710 404.000 344.710 404.280 ;
        RECT 345.550 404.000 346.550 404.280 ;
        RECT 347.390 404.000 348.390 404.280 ;
        RECT 349.230 404.000 350.230 404.280 ;
        RECT 351.070 404.000 352.070 404.280 ;
        RECT 352.910 404.000 353.450 404.280 ;
        RECT 354.290 404.000 355.290 404.280 ;
        RECT 356.130 404.000 357.130 404.280 ;
        RECT 357.970 404.000 358.970 404.280 ;
        RECT 359.810 404.000 360.810 404.280 ;
        RECT 361.650 404.000 362.650 404.280 ;
        RECT 363.490 404.000 364.490 404.280 ;
        RECT 365.330 404.000 366.330 404.280 ;
        RECT 367.170 404.000 367.710 404.280 ;
        RECT 368.550 404.000 369.550 404.280 ;
        RECT 370.390 404.000 371.390 404.280 ;
        RECT 372.230 404.000 373.230 404.280 ;
        RECT 374.070 404.000 375.070 404.280 ;
        RECT 375.910 404.000 376.910 404.280 ;
        RECT 377.750 404.000 378.750 404.280 ;
        RECT 379.590 404.000 380.590 404.280 ;
        RECT 381.430 404.000 382.430 404.280 ;
        RECT 383.270 404.000 383.810 404.280 ;
        RECT 384.650 404.000 385.650 404.280 ;
        RECT 386.490 404.000 387.490 404.280 ;
        RECT 388.330 404.000 389.330 404.280 ;
        RECT 390.170 404.000 391.170 404.280 ;
        RECT 392.010 404.000 393.010 404.280 ;
        RECT 393.850 404.000 394.850 404.280 ;
        RECT 395.690 404.000 396.690 404.280 ;
        RECT 397.530 404.000 398.530 404.280 ;
        RECT 399.370 404.000 399.910 404.280 ;
        RECT 400.750 404.000 401.750 404.280 ;
        RECT 402.590 404.000 403.590 404.280 ;
        RECT 404.430 404.000 405.430 404.280 ;
        RECT 406.270 404.000 407.270 404.280 ;
        RECT 408.110 404.000 409.110 404.280 ;
        RECT 409.950 404.000 410.950 404.280 ;
        RECT 411.790 404.000 412.790 404.280 ;
        RECT 413.630 404.000 414.170 404.280 ;
        RECT 415.010 404.000 416.010 404.280 ;
        RECT 416.850 404.000 417.850 404.280 ;
        RECT 418.690 404.000 419.690 404.280 ;
        RECT 420.530 404.000 421.530 404.280 ;
        RECT 422.370 404.000 423.370 404.280 ;
        RECT 424.210 404.000 425.210 404.280 ;
        RECT 426.050 404.000 427.050 404.280 ;
        RECT 427.890 404.000 428.890 404.280 ;
        RECT 429.730 404.000 430.270 404.280 ;
        RECT 431.110 404.000 432.110 404.280 ;
        RECT 432.950 404.000 433.950 404.280 ;
        RECT 434.790 404.000 435.790 404.280 ;
        RECT 436.630 404.000 437.630 404.280 ;
        RECT 438.470 404.000 439.470 404.280 ;
        RECT 440.310 404.000 441.310 404.280 ;
        RECT 442.150 404.000 443.150 404.280 ;
        RECT 443.990 404.000 444.530 404.280 ;
        RECT 445.370 404.000 446.370 404.280 ;
        RECT 447.210 404.000 448.210 404.280 ;
        RECT 449.050 404.000 450.050 404.280 ;
        RECT 450.890 404.000 451.890 404.280 ;
        RECT 452.730 404.000 453.730 404.280 ;
        RECT 454.570 404.000 455.570 404.280 ;
        RECT 456.410 404.000 457.410 404.280 ;
        RECT 458.250 404.000 459.250 404.280 ;
        RECT 460.090 404.000 460.630 404.280 ;
        RECT 461.470 404.000 462.470 404.280 ;
        RECT 463.310 404.000 464.310 404.280 ;
        RECT 465.150 404.000 466.150 404.280 ;
        RECT 466.990 404.000 467.990 404.280 ;
        RECT 468.830 404.000 469.830 404.280 ;
        RECT 470.670 404.000 471.670 404.280 ;
        RECT 472.510 404.000 473.510 404.280 ;
        RECT 474.350 404.000 474.890 404.280 ;
        RECT 475.730 404.000 476.730 404.280 ;
        RECT 477.570 404.000 478.570 404.280 ;
        RECT 479.410 404.000 480.410 404.280 ;
        RECT 481.250 404.000 482.250 404.280 ;
        RECT 483.090 404.000 484.090 404.280 ;
        RECT 484.930 404.000 485.930 404.280 ;
        RECT 486.770 404.000 487.770 404.280 ;
        RECT 488.610 404.000 489.610 404.280 ;
        RECT 490.450 404.000 490.990 404.280 ;
        RECT 491.830 404.000 492.830 404.280 ;
        RECT 493.670 404.000 494.670 404.280 ;
        RECT 495.510 404.000 496.510 404.280 ;
        RECT 497.350 404.000 498.350 404.280 ;
        RECT 499.190 404.000 500.190 404.280 ;
        RECT 501.030 404.000 502.030 404.280 ;
        RECT 502.870 404.000 503.870 404.280 ;
        RECT 504.710 404.000 505.250 404.280 ;
        RECT 506.090 404.000 507.090 404.280 ;
        RECT 507.930 404.000 508.930 404.280 ;
        RECT 509.770 404.000 510.770 404.280 ;
        RECT 511.610 404.000 512.610 404.280 ;
        RECT 513.450 404.000 514.450 404.280 ;
        RECT 515.290 404.000 516.290 404.280 ;
        RECT 517.130 404.000 518.130 404.280 ;
        RECT 518.970 404.000 519.970 404.280 ;
        RECT 520.810 404.000 521.350 404.280 ;
        RECT 522.190 404.000 523.190 404.280 ;
        RECT 524.030 404.000 525.030 404.280 ;
        RECT 525.870 404.000 526.870 404.280 ;
        RECT 527.710 404.000 528.710 404.280 ;
        RECT 529.550 404.000 530.550 404.280 ;
        RECT 531.390 404.000 532.390 404.280 ;
        RECT 533.230 404.000 534.230 404.280 ;
        RECT 535.070 404.000 535.610 404.280 ;
        RECT 536.450 404.000 537.450 404.280 ;
        RECT 538.290 404.000 539.290 404.280 ;
        RECT 540.130 404.000 541.130 404.280 ;
        RECT 541.970 404.000 542.970 404.280 ;
        RECT 543.810 404.000 544.810 404.280 ;
        RECT 545.650 404.000 546.650 404.280 ;
        RECT 547.490 404.000 548.490 404.280 ;
        RECT 549.330 404.000 550.330 404.280 ;
        RECT 551.170 404.000 551.710 404.280 ;
        RECT 552.550 404.000 553.550 404.280 ;
        RECT 554.390 404.000 555.390 404.280 ;
        RECT 556.230 404.000 557.230 404.280 ;
        RECT 558.070 404.000 559.070 404.280 ;
        RECT 559.910 404.000 560.910 404.280 ;
        RECT 561.750 404.000 562.750 404.280 ;
        RECT 563.590 404.000 564.590 404.280 ;
        RECT 565.430 404.000 566.430 404.280 ;
        RECT 567.270 404.000 567.810 404.280 ;
        RECT 568.650 404.000 569.650 404.280 ;
        RECT 570.490 404.000 571.490 404.280 ;
        RECT 572.330 404.000 573.330 404.280 ;
        RECT 574.170 404.000 575.170 404.280 ;
        RECT 576.010 404.000 577.010 404.280 ;
        RECT 577.850 404.000 578.850 404.280 ;
        RECT 579.690 404.000 580.690 404.280 ;
        RECT 581.530 404.000 582.070 404.280 ;
        RECT 582.910 404.000 583.910 404.280 ;
        RECT 584.750 404.000 585.750 404.280 ;
        RECT 586.590 404.000 587.590 404.280 ;
        RECT 588.430 404.000 589.430 404.280 ;
        RECT 590.270 404.000 591.270 404.280 ;
        RECT 592.110 404.000 593.110 404.280 ;
        RECT 593.950 404.000 594.950 404.280 ;
        RECT 595.790 404.000 596.790 404.280 ;
        RECT 597.630 404.000 598.170 404.280 ;
        RECT 599.010 404.000 600.010 404.280 ;
        RECT 600.850 404.000 601.850 404.280 ;
        RECT 602.690 404.000 603.690 404.280 ;
        RECT 604.530 404.000 605.530 404.280 ;
        RECT 606.370 404.000 607.370 404.280 ;
        RECT 608.210 404.000 609.210 404.280 ;
        RECT 610.050 404.000 611.050 404.280 ;
        RECT 611.890 404.000 612.430 404.280 ;
        RECT 613.270 404.000 614.270 404.280 ;
        RECT 615.110 404.000 616.110 404.280 ;
        RECT 616.950 404.000 617.950 404.280 ;
        RECT 618.790 404.000 619.790 404.280 ;
        RECT 620.630 404.000 621.630 404.280 ;
        RECT 622.470 404.000 623.470 404.280 ;
        RECT 624.310 404.000 625.310 404.280 ;
        RECT 626.150 404.000 627.150 404.280 ;
        RECT 627.990 404.000 628.530 404.280 ;
        RECT 629.370 404.000 630.370 404.280 ;
        RECT 631.210 404.000 632.210 404.280 ;
        RECT 633.050 404.000 634.050 404.280 ;
        RECT 634.890 404.000 635.890 404.280 ;
        RECT 636.730 404.000 637.730 404.280 ;
        RECT 638.570 404.000 639.570 404.280 ;
        RECT 640.410 404.000 641.410 404.280 ;
        RECT 642.250 404.000 642.790 404.280 ;
        RECT 643.630 404.000 644.630 404.280 ;
        RECT 645.470 404.000 646.470 404.280 ;
        RECT 647.310 404.000 648.310 404.280 ;
        RECT 649.150 404.000 650.150 404.280 ;
        RECT 650.990 404.000 651.990 404.280 ;
        RECT 652.830 404.000 653.830 404.280 ;
        RECT 654.670 404.000 655.670 404.280 ;
        RECT 656.510 404.000 657.510 404.280 ;
        RECT 658.350 404.000 658.890 404.280 ;
        RECT 659.730 404.000 660.730 404.280 ;
        RECT 661.570 404.000 662.570 404.280 ;
        RECT 663.410 404.000 664.410 404.280 ;
        RECT 665.250 404.000 666.250 404.280 ;
        RECT 667.090 404.000 668.090 404.280 ;
        RECT 668.930 404.000 669.930 404.280 ;
        RECT 670.770 404.000 671.770 404.280 ;
        RECT 672.610 404.000 673.150 404.280 ;
        RECT 673.990 404.000 674.990 404.280 ;
        RECT 675.830 404.000 676.830 404.280 ;
        RECT 677.670 404.000 678.670 404.280 ;
        RECT 679.510 404.000 680.510 404.280 ;
        RECT 681.350 404.000 682.350 404.280 ;
        RECT 683.190 404.000 684.190 404.280 ;
        RECT 685.030 404.000 686.030 404.280 ;
        RECT 686.870 404.000 687.870 404.280 ;
        RECT 688.710 404.000 689.250 404.280 ;
        RECT 690.090 404.000 691.090 404.280 ;
        RECT 691.930 404.000 692.930 404.280 ;
        RECT 693.770 404.000 694.770 404.280 ;
        RECT 695.610 404.000 696.610 404.280 ;
        RECT 697.450 404.000 698.450 404.280 ;
        RECT 699.290 404.000 700.290 404.280 ;
        RECT 701.130 404.000 702.130 404.280 ;
        RECT 702.970 404.000 703.510 404.280 ;
        RECT 704.350 404.000 705.350 404.280 ;
        RECT 706.190 404.000 707.190 404.280 ;
        RECT 708.030 404.000 709.030 404.280 ;
        RECT 709.870 404.000 710.870 404.280 ;
        RECT 711.710 404.000 712.710 404.280 ;
        RECT 713.550 404.000 714.550 404.280 ;
        RECT 715.390 404.000 716.390 404.280 ;
        RECT 717.230 404.000 718.230 404.280 ;
        RECT 719.070 404.000 719.610 404.280 ;
        RECT 720.450 404.000 721.450 404.280 ;
        RECT 722.290 404.000 723.290 404.280 ;
        RECT 724.130 404.000 725.130 404.280 ;
        RECT 725.970 404.000 726.970 404.280 ;
        RECT 727.810 404.000 728.810 404.280 ;
        RECT 729.650 404.000 730.650 404.280 ;
        RECT 731.490 404.000 732.490 404.280 ;
        RECT 733.330 404.000 733.870 404.280 ;
        RECT 734.710 404.000 735.710 404.280 ;
        RECT 736.550 404.000 737.550 404.280 ;
        RECT 738.390 404.000 739.390 404.280 ;
        RECT 740.230 404.000 741.230 404.280 ;
        RECT 742.070 404.000 743.070 404.280 ;
        RECT 743.910 404.000 744.910 404.280 ;
        RECT 745.750 404.000 746.750 404.280 ;
        RECT 747.590 404.000 748.590 404.280 ;
        RECT 749.430 404.000 749.970 404.280 ;
        RECT 750.810 404.000 751.810 404.280 ;
        RECT 752.650 404.000 753.650 404.280 ;
        RECT 754.490 404.000 755.490 404.280 ;
        RECT 756.330 404.000 757.330 404.280 ;
        RECT 758.170 404.000 759.170 404.280 ;
        RECT 760.010 404.000 761.010 404.280 ;
        RECT 761.850 404.000 762.850 404.280 ;
        RECT 763.690 404.000 764.690 404.280 ;
        RECT 765.530 404.000 766.070 404.280 ;
        RECT 766.910 404.000 767.910 404.280 ;
        RECT 768.750 404.000 769.750 404.280 ;
        RECT 770.590 404.000 771.590 404.280 ;
        RECT 772.430 404.000 773.430 404.280 ;
        RECT 774.270 404.000 775.270 404.280 ;
        RECT 776.110 404.000 777.110 404.280 ;
        RECT 777.950 404.000 778.950 404.280 ;
        RECT 779.790 404.000 780.330 404.280 ;
        RECT 781.170 404.000 782.170 404.280 ;
        RECT 783.010 404.000 784.010 404.280 ;
        RECT 784.850 404.000 785.850 404.280 ;
        RECT 786.690 404.000 787.690 404.280 ;
        RECT 788.530 404.000 789.530 404.280 ;
        RECT 790.370 404.000 791.370 404.280 ;
        RECT 792.210 404.000 793.210 404.280 ;
        RECT 794.050 404.000 795.050 404.280 ;
        RECT 795.890 404.000 796.430 404.280 ;
        RECT 797.270 404.000 798.270 404.280 ;
        RECT 799.110 404.000 800.110 404.280 ;
        RECT 800.950 404.000 801.950 404.280 ;
        RECT 802.790 404.000 803.790 404.280 ;
        RECT 804.630 404.000 805.630 404.280 ;
        RECT 806.470 404.000 807.470 404.280 ;
        RECT 808.310 404.000 809.310 404.280 ;
        RECT 810.150 404.000 810.690 404.280 ;
        RECT 811.530 404.000 812.530 404.280 ;
        RECT 813.370 404.000 814.370 404.280 ;
        RECT 815.210 404.000 816.210 404.280 ;
        RECT 817.050 404.000 818.050 404.280 ;
        RECT 818.890 404.000 819.890 404.280 ;
        RECT 820.730 404.000 821.730 404.280 ;
        RECT 822.570 404.000 823.570 404.280 ;
        RECT 824.410 404.000 825.410 404.280 ;
        RECT 826.250 404.000 826.790 404.280 ;
        RECT 827.630 404.000 828.630 404.280 ;
        RECT 829.470 404.000 830.470 404.280 ;
        RECT 831.310 404.000 832.310 404.280 ;
        RECT 833.150 404.000 834.150 404.280 ;
        RECT 834.990 404.000 835.990 404.280 ;
        RECT 836.830 404.000 837.830 404.280 ;
        RECT 838.670 404.000 839.670 404.280 ;
        RECT 840.510 404.000 841.050 404.280 ;
        RECT 841.890 404.000 842.890 404.280 ;
        RECT 843.730 404.000 844.730 404.280 ;
        RECT 845.570 404.000 846.570 404.280 ;
        RECT 847.410 404.000 848.410 404.280 ;
        RECT 849.250 404.000 850.250 404.280 ;
        RECT 851.090 404.000 852.090 404.280 ;
        RECT 852.930 404.000 853.930 404.280 ;
        RECT 854.770 404.000 855.770 404.280 ;
        RECT 856.610 404.000 857.150 404.280 ;
        RECT 857.990 404.000 858.990 404.280 ;
        RECT 859.830 404.000 860.830 404.280 ;
        RECT 861.670 404.000 862.670 404.280 ;
        RECT 863.510 404.000 864.510 404.280 ;
        RECT 865.350 404.000 866.350 404.280 ;
        RECT 867.190 404.000 868.190 404.280 ;
        RECT 869.030 404.000 870.030 404.280 ;
        RECT 870.870 404.000 871.410 404.280 ;
        RECT 872.250 404.000 873.250 404.280 ;
        RECT 874.090 404.000 875.090 404.280 ;
        RECT 875.930 404.000 876.930 404.280 ;
        RECT 877.770 404.000 878.770 404.280 ;
        RECT 879.610 404.000 880.610 404.280 ;
        RECT 881.450 404.000 882.450 404.280 ;
        RECT 883.290 404.000 884.290 404.280 ;
        RECT 885.130 404.000 886.130 404.280 ;
        RECT 886.970 404.000 887.510 404.280 ;
        RECT 888.350 404.000 889.350 404.280 ;
        RECT 890.190 404.000 891.190 404.280 ;
        RECT 892.030 404.000 893.030 404.280 ;
        RECT 893.870 404.000 894.870 404.280 ;
        RECT 895.710 404.000 896.710 404.280 ;
        RECT 897.550 404.000 898.550 404.280 ;
        RECT 899.390 404.000 900.390 404.280 ;
        RECT 901.230 404.000 901.770 404.280 ;
        RECT 902.610 404.000 903.610 404.280 ;
        RECT 904.450 404.000 905.450 404.280 ;
        RECT 906.290 404.000 907.290 404.280 ;
        RECT 908.130 404.000 909.130 404.280 ;
        RECT 909.970 404.000 910.970 404.280 ;
        RECT 911.810 404.000 912.810 404.280 ;
        RECT 913.650 404.000 914.650 404.280 ;
        RECT 915.490 404.000 916.490 404.280 ;
        RECT 917.330 404.000 917.870 404.280 ;
        RECT 918.710 404.000 919.710 404.280 ;
        RECT 920.550 404.000 921.550 404.280 ;
        RECT 922.390 404.000 923.390 404.280 ;
        RECT 924.230 404.000 925.230 404.280 ;
        RECT 926.070 404.000 927.070 404.280 ;
        RECT 927.910 404.000 928.910 404.280 ;
        RECT 929.750 404.000 930.750 404.280 ;
        RECT 931.590 404.000 932.590 404.280 ;
        RECT 933.430 404.000 933.970 404.280 ;
        RECT 934.810 404.000 935.810 404.280 ;
        RECT 936.650 404.000 937.650 404.280 ;
        RECT 938.490 404.000 939.490 404.280 ;
        RECT 940.330 404.000 941.330 404.280 ;
        RECT 942.170 404.000 943.170 404.280 ;
        RECT 944.010 404.000 945.010 404.280 ;
        RECT 945.850 404.000 946.850 404.280 ;
        RECT 947.690 404.000 948.230 404.280 ;
        RECT 949.070 404.000 950.070 404.280 ;
        RECT 950.910 404.000 951.910 404.280 ;
        RECT 952.750 404.000 953.750 404.280 ;
        RECT 954.590 404.000 955.590 404.280 ;
        RECT 956.430 404.000 957.430 404.280 ;
        RECT 958.270 404.000 959.270 404.280 ;
        RECT 960.110 404.000 961.110 404.280 ;
        RECT 961.950 404.000 962.950 404.280 ;
        RECT 963.790 404.000 964.330 404.280 ;
        RECT 965.170 404.000 966.170 404.280 ;
        RECT 967.010 404.000 968.010 404.280 ;
        RECT 968.850 404.000 969.850 404.280 ;
        RECT 970.690 404.000 971.690 404.280 ;
        RECT 972.530 404.000 973.530 404.280 ;
        RECT 974.370 404.000 975.370 404.280 ;
        RECT 976.210 404.000 977.210 404.280 ;
        RECT 978.050 404.000 978.590 404.280 ;
        RECT 979.430 404.000 980.430 404.280 ;
        RECT 981.270 404.000 982.270 404.280 ;
        RECT 983.110 404.000 984.110 404.280 ;
        RECT 984.950 404.000 985.950 404.280 ;
        RECT 986.790 404.000 987.790 404.280 ;
        RECT 988.630 404.000 989.630 404.280 ;
        RECT 990.470 404.000 991.470 404.280 ;
        RECT 992.310 404.000 993.310 404.280 ;
        RECT 994.150 404.000 994.690 404.280 ;
        RECT 995.530 404.000 996.530 404.280 ;
        RECT 997.370 404.000 998.370 404.280 ;
        RECT 999.210 404.000 1000.210 404.280 ;
        RECT 1001.050 404.000 1002.050 404.280 ;
        RECT 1002.890 404.000 1003.890 404.280 ;
        RECT 1004.730 404.000 1005.730 404.280 ;
        RECT 1006.570 404.000 1007.570 404.280 ;
        RECT 1008.410 404.000 1008.950 404.280 ;
        RECT 1009.790 404.000 1010.790 404.280 ;
        RECT 1011.630 404.000 1012.630 404.280 ;
        RECT 1013.470 404.000 1014.470 404.280 ;
        RECT 1015.310 404.000 1016.310 404.280 ;
        RECT 1017.150 404.000 1018.150 404.280 ;
        RECT 1018.990 404.000 1019.990 404.280 ;
        RECT 1020.830 404.000 1021.830 404.280 ;
        RECT 1022.670 404.000 1023.670 404.280 ;
        RECT 1024.510 404.000 1025.050 404.280 ;
        RECT 1025.890 404.000 1026.890 404.280 ;
        RECT 1027.730 404.000 1028.730 404.280 ;
        RECT 1029.570 404.000 1030.570 404.280 ;
        RECT 1031.410 404.000 1032.410 404.280 ;
        RECT 1033.250 404.000 1034.250 404.280 ;
        RECT 1035.090 404.000 1036.090 404.280 ;
        RECT 1036.930 404.000 1037.930 404.280 ;
        RECT 1038.770 404.000 1039.310 404.280 ;
        RECT 1040.150 404.000 1041.150 404.280 ;
        RECT 1041.990 404.000 1042.990 404.280 ;
        RECT 1043.830 404.000 1044.830 404.280 ;
        RECT 1045.670 404.000 1046.670 404.280 ;
        RECT 1047.510 404.000 1048.510 404.280 ;
        RECT 1049.350 404.000 1050.350 404.280 ;
        RECT 1051.190 404.000 1052.190 404.280 ;
        RECT 1053.030 404.000 1054.030 404.280 ;
        RECT 1054.870 404.000 1055.410 404.280 ;
        RECT 1056.250 404.000 1057.250 404.280 ;
        RECT 1058.090 404.000 1059.090 404.280 ;
        RECT 1059.930 404.000 1060.930 404.280 ;
        RECT 1061.770 404.000 1062.770 404.280 ;
        RECT 1063.610 404.000 1064.610 404.280 ;
        RECT 1065.450 404.000 1066.450 404.280 ;
        RECT 1067.290 404.000 1068.290 404.280 ;
        RECT 1069.130 404.000 1069.670 404.280 ;
        RECT 1070.510 404.000 1071.510 404.280 ;
        RECT 1072.350 404.000 1073.350 404.280 ;
        RECT 1074.190 404.000 1075.190 404.280 ;
        RECT 1076.030 404.000 1077.030 404.280 ;
        RECT 1077.870 404.000 1078.870 404.280 ;
        RECT 1079.710 404.000 1080.710 404.280 ;
        RECT 1081.550 404.000 1082.550 404.280 ;
        RECT 1083.390 404.000 1084.390 404.280 ;
        RECT 1085.230 404.000 1085.770 404.280 ;
        RECT 1086.610 404.000 1087.610 404.280 ;
        RECT 1088.450 404.000 1089.450 404.280 ;
        RECT 1090.290 404.000 1090.930 404.280 ;
      LAYER met2 ;
        RECT 200.550 400.000 200.830 404.000 ;
      LAYER met3 ;
        RECT 204.000 957.960 1096.000 988.705 ;
        RECT 204.400 956.560 1096.000 957.960 ;
        RECT 204.000 940.280 1096.000 956.560 ;
        RECT 204.000 938.880 1095.600 940.280 ;
        RECT 204.000 872.280 1096.000 938.880 ;
        RECT 204.400 870.880 1096.000 872.280 ;
        RECT 204.000 820.600 1096.000 870.880 ;
        RECT 204.000 819.200 1095.600 820.600 ;
        RECT 204.000 786.600 1096.000 819.200 ;
        RECT 204.400 785.200 1096.000 786.600 ;
        RECT 204.000 700.920 1096.000 785.200 ;
        RECT 204.400 700.240 1096.000 700.920 ;
        RECT 204.400 699.520 1095.600 700.240 ;
        RECT 204.000 698.840 1095.600 699.520 ;
        RECT 204.000 615.240 1096.000 698.840 ;
        RECT 204.400 613.840 1096.000 615.240 ;
        RECT 204.000 580.560 1096.000 613.840 ;
        RECT 204.000 579.160 1095.600 580.560 ;
        RECT 204.000 529.560 1096.000 579.160 ;
        RECT 204.400 528.160 1096.000 529.560 ;
        RECT 204.000 460.880 1096.000 528.160 ;
        RECT 204.000 459.480 1095.600 460.880 ;
        RECT 204.000 443.880 1096.000 459.480 ;
        RECT 204.400 442.480 1096.000 443.880 ;
        RECT 204.000 410.715 1096.000 442.480 ;
      LAYER met4 ;
        RECT 640.975 430.775 681.440 987.345 ;
        RECT 683.840 430.775 684.545 987.345 ;
  END
END user_project_wrapper
END LIBRARY

