



`default_nettype none
/*
*  *-------------------------------------------------------------
*  *
*  * user_project_wrapper also incorporating an analog block
*  *
*  * This wrapper enumerates all of the pins available to
*    the
*  * user for the user project.
*  *
*  * An example user project is provided in
*    this wrapper.  The
*  * example should be removed and replaced
*    with the actual
*  * user project.
*  *
*  *-------------------------------------------------------------
*  *              */
`ifndef MPRJ_IO_PADS
	`define MPRJ_IO_PADS 38
`endif

module user_project_wrapper (
	`ifdef USE_POWER_PINS
		inout vdda1,	// User area 1 3.3V supply
		inout vdda2,	// User area 2 3.3V supply
		inout vssa1,	// User area 1 analog ground
		inout vssa2,	// User area 2 analog ground
		inout vccd1,	// User area 1 1.8V supply
		inout vccd2,	// User area 2 1.8v supply
		inout vssd1,	// User area 1 digital ground
		inout vssd2,	// User area 2 digital ground
	`endif

// Wishbone Slave ports (WB MI A)
 input wb_clk_i,
 input wb_rst_i,
 input wbs_stb_i,
 input wbs_cyc_i,
 input wbs_we_i,
 input [3:0] wbs_sel_i,
 input [31:0] wbs_dat_i,
 input [31:0] wbs_adr_i,

 output wbs_ack_o,
 output [31:0] wbs_dat_o,

// Logic Analyzer Signals
input  [127:0] la_data_in,
output [127:0] la_data_out,
input  [127:0] la_oenb,

// IOs
input  [`MPRJ_IO_PADS-1:0] io_in,
output [`MPRJ_IO_PADS-1:0] io_out,
output [`MPRJ_IO_PADS-1:0] io_oeb,

// Analog (direct connection to GPIO pad---use with caution)
// Note that analog I/O is not available on the 7 lowest-numbered
// GPIO pads, and so the analog_io indexing is offset from the
// GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
 inout [`MPRJ_IO_PADS-10:0] analog_io,

// Independent clock (on independent integer divider)
 input   user_clock2,

// User maskable interrupt signals
 output [2:0] user_irq
 );

 /*--------------------------------------*/
 /* User project is instantiated  here   */
 /*--------------------------------------*/

   // `include "gl/macro_10.v"
  //  `include "gl/macro_13.v"
macro_13 u_macro_13 (
	 
	`ifdef USE_POWER_PINS
	        .vdda1(vdda1),	// User area 1 3.3V supply
		.vdda2(vdda2),	// User area 2 3.3V supply
		.vssa1(vssa1),	// User area 1 analog ground
		.vssa2(vssa2),	// User area 2 analog ground
		.vccd1(vccd1),	// User area 1 1.8V supply
		.vccd2(vccd2),	// User area 2 1.8v supply
		.vssd1(vssd1),	// User area 1 digital ground
		.vssd2(vssd2),	// User area 2 digital ground
	 `endif
	 .wb_rst_i(wb_rst_i),
	 .wbs_stb_i(wbs_stb_i),
	 .wbs_cyc_i(wbs_cyc_i),
	 .wbs_we_i(wbs_we_i),
	 .wbs_sel_i(wbs_sel_i),
	 .wbs_dat_i(wbs_dat_i),
	 .wbs_adr_i(wbs_adr_i),
	 .wbs_ack_o(wbs_ack_o),
	 .wbs_dat_o(wbs_dat_o),
	 .la_data_in(la_data_in),
         .la_data_out(la_data_out),
	 .la_oenb(la_oenb),
	 .io_in(io_in),
	 .io_out(io_out),
	 .io_oeb(io_oeb),
	 .user_irq(user_irq),
	 .user_clock2(user_clock2),
	 .analog_io(analog_io)
 );

 macro_7 u_macro_7 (

	 `ifdef USE_POWER_PINS
		 .vdda1(vdda1),  // User area 1 3.3V supply
			 .vdda2(vdda2),  // User area 2 3.3V supply
			 .vssa1(vssa1),  // User area 1 analog ground
			 .vssa2(vssa2),  // User area 2 analog ground
			 .vccd1(vccd1),  // User area 1 1.8V supply
			 .vccd2(vccd2),  // User area 2 1.8v supply
			 .vssd1(vssd1),  // User area 1 digital ground
			 .vssd2(vssd2),  // User area 2 digital ground
		 `endif
		 .wb_rst_i(wb_rst_i),
			 .wbs_stb_i(wbs_stb_i),
			 .wbs_cyc_i(wbs_cyc_i),
			 .wbs_we_i(wbs_we_i),
			 .wbs_sel_i(wbs_sel_i),
			 .wbs_dat_i(wbs_dat_i),
			 .wbs_adr_i(wbs_adr_i),
			 .wbs_ack_o(wbs_ack_o),
			 .wbs_dat_o(wbs_dat_o),
			 .la_data_in(la_data_in),
			 .la_data_out(la_data_out),
			 .la_oenb(la_oenb),
			 .io_in(io_in),
			 .io_out(io_out),
			 .io_oeb(io_oeb),
			 .user_irq(user_irq),
			 .user_clock2(user_clock2),
			 .analog_io(analog_io)
		 );

macro_10 u_macro_10 (

`ifdef USE_POWER_PINS
.vdda1(vdda1),  // User area 1 3.3V supply
.vdda2(vdda2),  // User area 2 3.3V supply
.vssa1(vssa1),  // User area 1 analog ground
.vssa2(vssa2),  // User area 2 analog ground
.vccd1(vccd1),  // User area 1 1.8V supply
.vccd2(vccd2),  // User area 2 1.8v supply
.vssd1(vssd1),  // User area 1 digital ground
.vssd2(vssd2),  // User area 2 digital ground
`endif
.wb_rst_i(wb_rst_i),
	.wbs_stb_i(wbs_stb_i),
	.wbs_cyc_i(wbs_cyc_i),
	.wbs_we_i(wbs_we_i),
	.wbs_sel_i(wbs_sel_i),
	.wbs_dat_i(wbs_dat_i),
	.wbs_adr_i(wbs_adr_i),
	.wbs_ack_o(wbs_ack_o),
	.wbs_dat_o(wbs_dat_o),
	.la_data_in(la_data_in),
	.la_data_out(la_data_out),
	.la_oenb(la_oenb),
	.io_in(io_in),
	.io_out(io_out),
	.io_oeb(io_oeb),
	.user_irq(user_irq),
	.user_clock2(user_clock2),
	.analog_io(analog_io)
);

 endmodule	// user_project_wrapper

 `default_nettype wire
