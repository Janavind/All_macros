magic
tech sky130A
magscale 1 2
timestamp 1654527384
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 198 1844 49022 47864
<< metal2 >>
rect 202 49200 258 50000
rect 570 49200 626 50000
rect 938 49200 994 50000
rect 1398 49200 1454 50000
rect 1766 49200 1822 50000
rect 2226 49200 2282 50000
rect 2594 49200 2650 50000
rect 3054 49200 3110 50000
rect 3422 49200 3478 50000
rect 3882 49200 3938 50000
rect 4250 49200 4306 50000
rect 4618 49200 4674 50000
rect 5078 49200 5134 50000
rect 5446 49200 5502 50000
rect 5906 49200 5962 50000
rect 6274 49200 6330 50000
rect 6734 49200 6790 50000
rect 7102 49200 7158 50000
rect 7562 49200 7618 50000
rect 7930 49200 7986 50000
rect 8390 49200 8446 50000
rect 8758 49200 8814 50000
rect 9126 49200 9182 50000
rect 9586 49200 9642 50000
rect 9954 49200 10010 50000
rect 10414 49200 10470 50000
rect 10782 49200 10838 50000
rect 11242 49200 11298 50000
rect 11610 49200 11666 50000
rect 12070 49200 12126 50000
rect 12438 49200 12494 50000
rect 12806 49200 12862 50000
rect 13266 49200 13322 50000
rect 13634 49200 13690 50000
rect 14094 49200 14150 50000
rect 14462 49200 14518 50000
rect 14922 49200 14978 50000
rect 15290 49200 15346 50000
rect 15750 49200 15806 50000
rect 16118 49200 16174 50000
rect 16578 49200 16634 50000
rect 16946 49200 17002 50000
rect 17314 49200 17370 50000
rect 17774 49200 17830 50000
rect 18142 49200 18198 50000
rect 18602 49200 18658 50000
rect 18970 49200 19026 50000
rect 19430 49200 19486 50000
rect 19798 49200 19854 50000
rect 20258 49200 20314 50000
rect 20626 49200 20682 50000
rect 20994 49200 21050 50000
rect 21454 49200 21510 50000
rect 21822 49200 21878 50000
rect 22282 49200 22338 50000
rect 22650 49200 22706 50000
rect 23110 49200 23166 50000
rect 23478 49200 23534 50000
rect 23938 49200 23994 50000
rect 24306 49200 24362 50000
rect 24766 49200 24822 50000
rect 25134 49200 25190 50000
rect 25502 49200 25558 50000
rect 25962 49200 26018 50000
rect 26330 49200 26386 50000
rect 26790 49200 26846 50000
rect 27158 49200 27214 50000
rect 27618 49200 27674 50000
rect 27986 49200 28042 50000
rect 28446 49200 28502 50000
rect 28814 49200 28870 50000
rect 29274 49200 29330 50000
rect 29642 49200 29698 50000
rect 30010 49200 30066 50000
rect 30470 49200 30526 50000
rect 30838 49200 30894 50000
rect 31298 49200 31354 50000
rect 31666 49200 31722 50000
rect 32126 49200 32182 50000
rect 32494 49200 32550 50000
rect 32954 49200 33010 50000
rect 33322 49200 33378 50000
rect 33690 49200 33746 50000
rect 34150 49200 34206 50000
rect 34518 49200 34574 50000
rect 34978 49200 35034 50000
rect 35346 49200 35402 50000
rect 35806 49200 35862 50000
rect 36174 49200 36230 50000
rect 36634 49200 36690 50000
rect 37002 49200 37058 50000
rect 37462 49200 37518 50000
rect 37830 49200 37886 50000
rect 38198 49200 38254 50000
rect 38658 49200 38714 50000
rect 39026 49200 39082 50000
rect 39486 49200 39542 50000
rect 39854 49200 39910 50000
rect 40314 49200 40370 50000
rect 40682 49200 40738 50000
rect 41142 49200 41198 50000
rect 41510 49200 41566 50000
rect 41878 49200 41934 50000
rect 42338 49200 42394 50000
rect 42706 49200 42762 50000
rect 43166 49200 43222 50000
rect 43534 49200 43590 50000
rect 43994 49200 44050 50000
rect 44362 49200 44418 50000
rect 44822 49200 44878 50000
rect 45190 49200 45246 50000
rect 45650 49200 45706 50000
rect 46018 49200 46074 50000
rect 46386 49200 46442 50000
rect 46846 49200 46902 50000
rect 47214 49200 47270 50000
rect 47674 49200 47730 50000
rect 48042 49200 48098 50000
rect 48502 49200 48558 50000
rect 48870 49200 48926 50000
rect 49330 49200 49386 50000
rect 49698 49200 49754 50000
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 294 0 350 800
rect 386 0 442 800
rect 478 0 534 800
rect 570 0 626 800
rect 662 0 718 800
rect 754 0 810 800
rect 846 0 902 800
rect 938 0 994 800
rect 1030 0 1086 800
rect 1214 0 1270 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1490 0 1546 800
rect 1582 0 1638 800
rect 1674 0 1730 800
rect 1766 0 1822 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2134 0 2190 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2686 0 2742 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3054 0 3110 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3330 0 3386 800
rect 3422 0 3478 800
rect 3606 0 3662 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 3974 0 4030 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4250 0 4306 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4526 0 4582 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4894 0 4950 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5170 0 5226 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5446 0 5502 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
<< obsm2 >>
rect 314 49144 514 49314
rect 682 49144 882 49314
rect 1050 49144 1342 49314
rect 1510 49144 1710 49314
rect 1878 49144 2170 49314
rect 2338 49144 2538 49314
rect 2706 49144 2998 49314
rect 3166 49144 3366 49314
rect 3534 49144 3826 49314
rect 3994 49144 4194 49314
rect 4362 49144 4562 49314
rect 4730 49144 5022 49314
rect 5190 49144 5390 49314
rect 5558 49144 5850 49314
rect 6018 49144 6218 49314
rect 6386 49144 6678 49314
rect 6846 49144 7046 49314
rect 7214 49144 7506 49314
rect 7674 49144 7874 49314
rect 8042 49144 8334 49314
rect 8502 49144 8702 49314
rect 8870 49144 9070 49314
rect 9238 49144 9530 49314
rect 9698 49144 9898 49314
rect 10066 49144 10358 49314
rect 10526 49144 10726 49314
rect 10894 49144 11186 49314
rect 11354 49144 11554 49314
rect 11722 49144 12014 49314
rect 12182 49144 12382 49314
rect 12550 49144 12750 49314
rect 12918 49144 13210 49314
rect 13378 49144 13578 49314
rect 13746 49144 14038 49314
rect 14206 49144 14406 49314
rect 14574 49144 14866 49314
rect 15034 49144 15234 49314
rect 15402 49144 15694 49314
rect 15862 49144 16062 49314
rect 16230 49144 16522 49314
rect 16690 49144 16890 49314
rect 17058 49144 17258 49314
rect 17426 49144 17718 49314
rect 17886 49144 18086 49314
rect 18254 49144 18546 49314
rect 18714 49144 18914 49314
rect 19082 49144 19374 49314
rect 19542 49144 19742 49314
rect 19910 49144 20202 49314
rect 20370 49144 20570 49314
rect 20738 49144 20938 49314
rect 21106 49144 21398 49314
rect 21566 49144 21766 49314
rect 21934 49144 22226 49314
rect 22394 49144 22594 49314
rect 22762 49144 23054 49314
rect 23222 49144 23422 49314
rect 23590 49144 23882 49314
rect 24050 49144 24250 49314
rect 24418 49144 24710 49314
rect 24878 49144 25078 49314
rect 25246 49144 25446 49314
rect 25614 49144 25906 49314
rect 26074 49144 26274 49314
rect 26442 49144 26734 49314
rect 26902 49144 27102 49314
rect 27270 49144 27562 49314
rect 27730 49144 27930 49314
rect 28098 49144 28390 49314
rect 28558 49144 28758 49314
rect 28926 49144 29218 49314
rect 29386 49144 29586 49314
rect 29754 49144 29954 49314
rect 30122 49144 30414 49314
rect 30582 49144 30782 49314
rect 30950 49144 31242 49314
rect 31410 49144 31610 49314
rect 31778 49144 32070 49314
rect 32238 49144 32438 49314
rect 32606 49144 32898 49314
rect 33066 49144 33266 49314
rect 33434 49144 33634 49314
rect 33802 49144 34094 49314
rect 34262 49144 34462 49314
rect 34630 49144 34922 49314
rect 35090 49144 35290 49314
rect 35458 49144 35750 49314
rect 35918 49144 36118 49314
rect 36286 49144 36578 49314
rect 36746 49144 36946 49314
rect 37114 49144 37406 49314
rect 37574 49144 37774 49314
rect 37942 49144 38142 49314
rect 38310 49144 38602 49314
rect 38770 49144 38970 49314
rect 39138 49144 39430 49314
rect 39598 49144 39798 49314
rect 39966 49144 40258 49314
rect 40426 49144 40626 49314
rect 40794 49144 41086 49314
rect 41254 49144 41454 49314
rect 41622 49144 41822 49314
rect 41990 49144 42282 49314
rect 42450 49144 42650 49314
rect 42818 49144 43110 49314
rect 43278 49144 43478 49314
rect 43646 49144 43938 49314
rect 44106 49144 44306 49314
rect 44474 49144 44766 49314
rect 44934 49144 45134 49314
rect 45302 49144 45594 49314
rect 45762 49144 45962 49314
rect 46130 49144 46330 49314
rect 46498 49144 46790 49314
rect 46958 49144 47158 49314
rect 47326 49144 47618 49314
rect 47786 49144 47986 49314
rect 48154 49144 48446 49314
rect 48614 49144 48814 49314
rect 48982 49144 49016 49314
rect 204 856 49016 49144
rect 1142 800 1158 856
rect 2338 800 2354 856
rect 3534 800 3550 856
rect 4730 800 4746 856
rect 5926 800 5942 856
rect 7122 800 7138 856
rect 8318 800 8334 856
rect 9514 800 9530 856
rect 10710 800 10726 856
rect 11906 800 11922 856
rect 13102 800 13118 856
rect 14298 800 14314 856
rect 15494 800 15510 856
rect 16598 800 16614 856
rect 17794 800 17810 856
rect 18990 800 19006 856
rect 20186 800 20202 856
rect 21382 800 21398 856
rect 22578 800 22594 856
rect 23774 800 23790 856
rect 24970 800 24986 856
rect 26166 800 26182 856
rect 27362 800 27378 856
rect 28558 800 28574 856
rect 29754 800 29770 856
rect 30950 800 30966 856
rect 32146 800 32162 856
rect 33250 800 33266 856
rect 34446 800 34462 856
rect 35642 800 35658 856
rect 36838 800 36854 856
rect 38034 800 38050 856
rect 39230 800 39246 856
rect 40426 800 40442 856
rect 41622 800 41638 856
rect 42818 800 42834 856
rect 44014 800 44030 856
rect 45210 800 45226 856
rect 46406 800 46422 856
rect 47602 800 47618 856
rect 48798 800 48814 856
<< metal3 >>
rect 0 47472 800 47592
rect 49200 44888 50000 45008
rect 0 42440 800 42560
rect 0 37408 800 37528
rect 49200 34824 50000 34944
rect 0 32376 800 32496
rect 0 27480 800 27600
rect 49200 24896 50000 25016
rect 0 22448 800 22568
rect 0 17416 800 17536
rect 49200 14832 50000 14952
rect 0 12384 800 12504
rect 0 7352 800 7472
rect 49200 4904 50000 5024
rect 0 2456 800 2576
<< obsm3 >>
rect 1853 45088 49200 47565
rect 1853 44808 49120 45088
rect 1853 35024 49200 44808
rect 1853 34744 49120 35024
rect 1853 25096 49200 34744
rect 1853 24816 49120 25096
rect 1853 15032 49200 24816
rect 1853 14752 49120 15032
rect 1853 5104 49200 14752
rect 1853 4824 49120 5104
rect 1853 2143 49200 4824
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 20851 4115 31037 47565
<< labels >>
rlabel metal3 s 49200 4904 50000 5024 6 active
port 1 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal2 s 49054 0 49110 800 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal2 s 48502 49200 48558 50000 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal2 s 49146 0 49202 800 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal3 s 0 37408 800 37528 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 48870 49200 48926 50000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal3 s 49200 24896 50000 25016 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 49330 49200 49386 50000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal2 s 49238 0 49294 800 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal3 s 0 42440 800 42560 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 49200 34824 50000 34944 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal3 s 0 12384 800 12504 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 49330 0 49386 800 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 49698 49200 49754 50000 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal2 s 49422 0 49478 800 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal2 s 49514 0 49570 800 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 49606 0 49662 800 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 49698 0 49754 800 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal2 s 49790 0 49846 800 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal3 s 49200 44888 50000 45008 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal3 s 0 47472 800 47592 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal3 s 0 17416 800 17536 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 49200 14832 50000 14952 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 0 22448 800 22568 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal2 s 47214 49200 47270 50000 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 0 27480 800 27600 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal2 s 47674 49200 47730 50000 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 0 32376 800 32496 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 48042 49200 48098 50000 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 202 49200 258 50000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 12438 49200 12494 50000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 13634 49200 13690 50000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 14922 49200 14978 50000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 16118 49200 16174 50000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 17314 49200 17370 50000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 18602 49200 18658 50000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 19798 49200 19854 50000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 20994 49200 21050 50000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 22282 49200 22338 50000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 23478 49200 23534 50000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 1398 49200 1454 50000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 24766 49200 24822 50000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 25962 49200 26018 50000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 27158 49200 27214 50000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 28446 49200 28502 50000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 29642 49200 29698 50000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 30838 49200 30894 50000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 32126 49200 32182 50000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 33322 49200 33378 50000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 34518 49200 34574 50000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 35806 49200 35862 50000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 2594 49200 2650 50000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 37002 49200 37058 50000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 38198 49200 38254 50000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 39486 49200 39542 50000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 40682 49200 40738 50000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 41878 49200 41934 50000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 43166 49200 43222 50000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 44362 49200 44418 50000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 45650 49200 45706 50000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 3882 49200 3938 50000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 5078 49200 5134 50000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 6274 49200 6330 50000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 7562 49200 7618 50000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 8758 49200 8814 50000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 9954 49200 10010 50000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 11242 49200 11298 50000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 570 49200 626 50000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 12806 49200 12862 50000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 14094 49200 14150 50000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 15290 49200 15346 50000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 16578 49200 16634 50000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 17774 49200 17830 50000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 18970 49200 19026 50000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 20258 49200 20314 50000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 21454 49200 21510 50000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 22650 49200 22706 50000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 23938 49200 23994 50000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 1766 49200 1822 50000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 25134 49200 25190 50000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 26330 49200 26386 50000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 27618 49200 27674 50000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 28814 49200 28870 50000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 30010 49200 30066 50000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 31298 49200 31354 50000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 32494 49200 32550 50000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 33690 49200 33746 50000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 34978 49200 35034 50000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 36174 49200 36230 50000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 3054 49200 3110 50000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 37462 49200 37518 50000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 38658 49200 38714 50000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 39854 49200 39910 50000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 41142 49200 41198 50000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 42338 49200 42394 50000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 43534 49200 43590 50000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 44822 49200 44878 50000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 46018 49200 46074 50000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 4250 49200 4306 50000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 5446 49200 5502 50000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 6734 49200 6790 50000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 7930 49200 7986 50000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 9126 49200 9182 50000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 10414 49200 10470 50000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 11610 49200 11666 50000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 938 49200 994 50000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 13266 49200 13322 50000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 14462 49200 14518 50000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 15750 49200 15806 50000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 16946 49200 17002 50000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 18142 49200 18198 50000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 19430 49200 19486 50000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 20626 49200 20682 50000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 21822 49200 21878 50000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 23110 49200 23166 50000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 24306 49200 24362 50000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 2226 49200 2282 50000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 25502 49200 25558 50000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 26790 49200 26846 50000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 27986 49200 28042 50000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 29274 49200 29330 50000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 30470 49200 30526 50000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 31666 49200 31722 50000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 32954 49200 33010 50000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 34150 49200 34206 50000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 35346 49200 35402 50000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 36634 49200 36690 50000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 3422 49200 3478 50000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 37830 49200 37886 50000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 39026 49200 39082 50000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 40314 49200 40370 50000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 41510 49200 41566 50000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 42706 49200 42762 50000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 43994 49200 44050 50000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 45190 49200 45246 50000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 46386 49200 46442 50000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 4618 49200 4674 50000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 5906 49200 5962 50000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 7102 49200 7158 50000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 8390 49200 8446 50000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 9586 49200 9642 50000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 10782 49200 10838 50000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 12070 49200 12126 50000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 user_clock2
port 529 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 46846 49200 46902 50000 6 user_irq[1]
port 531 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 534 nsew ground input
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 570 0 626 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 294 0 350 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 1214 0 1270 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 846 0 902 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1758010
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_decap_3.magic.gds
string GDS_START 222892
<< end >>

