magic
tech sky130A
magscale 1 2
timestamp 1654044043
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 750 2128 178848 118176
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9586 119200 9642 120000
rect 11058 119200 11114 120000
rect 12530 119200 12586 120000
rect 14002 119200 14058 120000
rect 15474 119200 15530 120000
rect 16946 119200 17002 120000
rect 18418 119200 18474 120000
rect 19890 119200 19946 120000
rect 21362 119200 21418 120000
rect 22834 119200 22890 120000
rect 24306 119200 24362 120000
rect 25778 119200 25834 120000
rect 27250 119200 27306 120000
rect 28722 119200 28778 120000
rect 30194 119200 30250 120000
rect 31666 119200 31722 120000
rect 33138 119200 33194 120000
rect 34610 119200 34666 120000
rect 36082 119200 36138 120000
rect 37646 119200 37702 120000
rect 39118 119200 39174 120000
rect 40590 119200 40646 120000
rect 42062 119200 42118 120000
rect 43534 119200 43590 120000
rect 45006 119200 45062 120000
rect 46478 119200 46534 120000
rect 47950 119200 48006 120000
rect 49422 119200 49478 120000
rect 50894 119200 50950 120000
rect 52366 119200 52422 120000
rect 53838 119200 53894 120000
rect 55310 119200 55366 120000
rect 56782 119200 56838 120000
rect 58254 119200 58310 120000
rect 59726 119200 59782 120000
rect 61198 119200 61254 120000
rect 62670 119200 62726 120000
rect 64142 119200 64198 120000
rect 65614 119200 65670 120000
rect 67086 119200 67142 120000
rect 68558 119200 68614 120000
rect 70030 119200 70086 120000
rect 71502 119200 71558 120000
rect 73066 119200 73122 120000
rect 74538 119200 74594 120000
rect 76010 119200 76066 120000
rect 77482 119200 77538 120000
rect 78954 119200 79010 120000
rect 80426 119200 80482 120000
rect 81898 119200 81954 120000
rect 83370 119200 83426 120000
rect 84842 119200 84898 120000
rect 86314 119200 86370 120000
rect 87786 119200 87842 120000
rect 89258 119200 89314 120000
rect 90730 119200 90786 120000
rect 92202 119200 92258 120000
rect 93674 119200 93730 120000
rect 95146 119200 95202 120000
rect 96618 119200 96674 120000
rect 98090 119200 98146 120000
rect 99562 119200 99618 120000
rect 101034 119200 101090 120000
rect 102506 119200 102562 120000
rect 103978 119200 104034 120000
rect 105450 119200 105506 120000
rect 106922 119200 106978 120000
rect 108394 119200 108450 120000
rect 109958 119200 110014 120000
rect 111430 119200 111486 120000
rect 112902 119200 112958 120000
rect 114374 119200 114430 120000
rect 115846 119200 115902 120000
rect 117318 119200 117374 120000
rect 118790 119200 118846 120000
rect 120262 119200 120318 120000
rect 121734 119200 121790 120000
rect 123206 119200 123262 120000
rect 124678 119200 124734 120000
rect 126150 119200 126206 120000
rect 127622 119200 127678 120000
rect 129094 119200 129150 120000
rect 130566 119200 130622 120000
rect 132038 119200 132094 120000
rect 133510 119200 133566 120000
rect 134982 119200 135038 120000
rect 136454 119200 136510 120000
rect 137926 119200 137982 120000
rect 139398 119200 139454 120000
rect 140870 119200 140926 120000
rect 142342 119200 142398 120000
rect 143814 119200 143870 120000
rect 145378 119200 145434 120000
rect 146850 119200 146906 120000
rect 148322 119200 148378 120000
rect 149794 119200 149850 120000
rect 151266 119200 151322 120000
rect 152738 119200 152794 120000
rect 154210 119200 154266 120000
rect 155682 119200 155738 120000
rect 157154 119200 157210 120000
rect 158626 119200 158682 120000
rect 160098 119200 160154 120000
rect 161570 119200 161626 120000
rect 163042 119200 163098 120000
rect 164514 119200 164570 120000
rect 165986 119200 166042 120000
rect 167458 119200 167514 120000
rect 168930 119200 168986 120000
rect 170402 119200 170458 120000
rect 171874 119200 171930 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15750 0 15806 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26514 0 26570 800
rect 26882 0 26938 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31114 0 31170 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 43994 0 44050 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54390 0 54446 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57978 0 58034 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61474 0 61530 800
rect 61842 0 61898 800
rect 62210 0 62266 800
rect 62578 0 62634 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66166 0 66222 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 69018 0 69074 800
rect 69386 0 69442 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73618 0 73674 800
rect 73986 0 74042 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76838 0 76894 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78678 0 78734 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79690 0 79746 800
rect 80058 0 80114 800
rect 80426 0 80482 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86866 0 86922 800
rect 87234 0 87290 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90454 0 90510 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92938 0 92994 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100114 0 100170 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101494 0 101550 800
rect 101862 0 101918 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110786 0 110842 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112258 0 112314 800
rect 112626 0 112682 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114742 0 114798 800
rect 115110 0 115166 800
rect 115478 0 115534 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116490 0 116546 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118698 0 118754 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121182 0 121238 800
rect 121550 0 121606 800
rect 121918 0 121974 800
rect 122194 0 122250 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124402 0 124458 800
rect 124770 0 124826 800
rect 125138 0 125194 800
rect 125414 0 125470 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128266 0 128322 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130106 0 130162 800
rect 130474 0 130530 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132590 0 132646 800
rect 132958 0 133014 800
rect 133326 0 133382 800
rect 133694 0 133750 800
rect 134062 0 134118 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136178 0 136234 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139766 0 139822 800
rect 140134 0 140190 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142618 0 142674 800
rect 142986 0 143042 800
rect 143354 0 143410 800
rect 143630 0 143686 800
rect 143998 0 144054 800
rect 144366 0 144422 800
rect 144734 0 144790 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146850 0 146906 800
rect 147218 0 147274 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149426 0 149482 800
rect 149702 0 149758 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152646 0 152702 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153658 0 153714 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155130 0 155186 800
rect 155498 0 155554 800
rect 155774 0 155830 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156878 0 156934 800
rect 157246 0 157302 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158350 0 158406 800
rect 158718 0 158774 800
rect 158994 0 159050 800
rect 159362 0 159418 800
rect 159730 0 159786 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161846 0 161902 800
rect 162214 0 162270 800
rect 162582 0 162638 800
rect 162950 0 163006 800
rect 163318 0 163374 800
rect 163686 0 163742 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165066 0 165122 800
rect 165434 0 165490 800
rect 165802 0 165858 800
rect 166170 0 166226 800
rect 166538 0 166594 800
rect 166906 0 166962 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 167918 0 167974 800
rect 168286 0 168342 800
rect 168654 0 168710 800
rect 169022 0 169078 800
rect 169390 0 169446 800
rect 169758 0 169814 800
rect 170126 0 170182 800
rect 170494 0 170550 800
rect 170862 0 170918 800
rect 171138 0 171194 800
rect 171506 0 171562 800
rect 171874 0 171930 800
rect 172242 0 172298 800
rect 172610 0 172666 800
rect 172978 0 173034 800
rect 173346 0 173402 800
rect 173714 0 173770 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175094 0 175150 800
rect 175462 0 175518 800
rect 175830 0 175886 800
rect 176198 0 176254 800
rect 176566 0 176622 800
rect 176934 0 176990 800
rect 177210 0 177266 800
rect 177578 0 177634 800
rect 177946 0 178002 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
<< obsm2 >>
rect 866 119144 2170 119354
rect 2338 119144 3642 119354
rect 3810 119144 5114 119354
rect 5282 119144 6586 119354
rect 6754 119144 8058 119354
rect 8226 119144 9530 119354
rect 9698 119144 11002 119354
rect 11170 119144 12474 119354
rect 12642 119144 13946 119354
rect 14114 119144 15418 119354
rect 15586 119144 16890 119354
rect 17058 119144 18362 119354
rect 18530 119144 19834 119354
rect 20002 119144 21306 119354
rect 21474 119144 22778 119354
rect 22946 119144 24250 119354
rect 24418 119144 25722 119354
rect 25890 119144 27194 119354
rect 27362 119144 28666 119354
rect 28834 119144 30138 119354
rect 30306 119144 31610 119354
rect 31778 119144 33082 119354
rect 33250 119144 34554 119354
rect 34722 119144 36026 119354
rect 36194 119144 37590 119354
rect 37758 119144 39062 119354
rect 39230 119144 40534 119354
rect 40702 119144 42006 119354
rect 42174 119144 43478 119354
rect 43646 119144 44950 119354
rect 45118 119144 46422 119354
rect 46590 119144 47894 119354
rect 48062 119144 49366 119354
rect 49534 119144 50838 119354
rect 51006 119144 52310 119354
rect 52478 119144 53782 119354
rect 53950 119144 55254 119354
rect 55422 119144 56726 119354
rect 56894 119144 58198 119354
rect 58366 119144 59670 119354
rect 59838 119144 61142 119354
rect 61310 119144 62614 119354
rect 62782 119144 64086 119354
rect 64254 119144 65558 119354
rect 65726 119144 67030 119354
rect 67198 119144 68502 119354
rect 68670 119144 69974 119354
rect 70142 119144 71446 119354
rect 71614 119144 73010 119354
rect 73178 119144 74482 119354
rect 74650 119144 75954 119354
rect 76122 119144 77426 119354
rect 77594 119144 78898 119354
rect 79066 119144 80370 119354
rect 80538 119144 81842 119354
rect 82010 119144 83314 119354
rect 83482 119144 84786 119354
rect 84954 119144 86258 119354
rect 86426 119144 87730 119354
rect 87898 119144 89202 119354
rect 89370 119144 90674 119354
rect 90842 119144 92146 119354
rect 92314 119144 93618 119354
rect 93786 119144 95090 119354
rect 95258 119144 96562 119354
rect 96730 119144 98034 119354
rect 98202 119144 99506 119354
rect 99674 119144 100978 119354
rect 101146 119144 102450 119354
rect 102618 119144 103922 119354
rect 104090 119144 105394 119354
rect 105562 119144 106866 119354
rect 107034 119144 108338 119354
rect 108506 119144 109902 119354
rect 110070 119144 111374 119354
rect 111542 119144 112846 119354
rect 113014 119144 114318 119354
rect 114486 119144 115790 119354
rect 115958 119144 117262 119354
rect 117430 119144 118734 119354
rect 118902 119144 120206 119354
rect 120374 119144 121678 119354
rect 121846 119144 123150 119354
rect 123318 119144 124622 119354
rect 124790 119144 126094 119354
rect 126262 119144 127566 119354
rect 127734 119144 129038 119354
rect 129206 119144 130510 119354
rect 130678 119144 131982 119354
rect 132150 119144 133454 119354
rect 133622 119144 134926 119354
rect 135094 119144 136398 119354
rect 136566 119144 137870 119354
rect 138038 119144 139342 119354
rect 139510 119144 140814 119354
rect 140982 119144 142286 119354
rect 142454 119144 143758 119354
rect 143926 119144 145322 119354
rect 145490 119144 146794 119354
rect 146962 119144 148266 119354
rect 148434 119144 149738 119354
rect 149906 119144 151210 119354
rect 151378 119144 152682 119354
rect 152850 119144 154154 119354
rect 154322 119144 155626 119354
rect 155794 119144 157098 119354
rect 157266 119144 158570 119354
rect 158738 119144 160042 119354
rect 160210 119144 161514 119354
rect 161682 119144 162986 119354
rect 163154 119144 164458 119354
rect 164626 119144 165930 119354
rect 166098 119144 167402 119354
rect 167570 119144 168874 119354
rect 169042 119144 170346 119354
rect 170514 119144 171818 119354
rect 171986 119144 173290 119354
rect 173458 119144 174762 119354
rect 174930 119144 176234 119354
rect 176402 119144 177706 119354
rect 177874 119144 178186 119354
rect 756 856 178186 119144
rect 866 800 1066 856
rect 1234 800 1434 856
rect 1602 800 1802 856
rect 1970 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3918 856
rect 4086 800 4286 856
rect 4454 800 4654 856
rect 4822 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6126 856
rect 6294 800 6402 856
rect 6570 800 6770 856
rect 6938 800 7138 856
rect 7306 800 7506 856
rect 7674 800 7874 856
rect 8042 800 8242 856
rect 8410 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9254 856
rect 9422 800 9622 856
rect 9790 800 9990 856
rect 10158 800 10358 856
rect 10526 800 10726 856
rect 10894 800 11094 856
rect 11262 800 11462 856
rect 11630 800 11830 856
rect 11998 800 12198 856
rect 12366 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13578 856
rect 13746 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14682 856
rect 14850 800 15050 856
rect 15218 800 15326 856
rect 15494 800 15694 856
rect 15862 800 16062 856
rect 16230 800 16430 856
rect 16598 800 16798 856
rect 16966 800 17166 856
rect 17334 800 17534 856
rect 17702 800 17902 856
rect 18070 800 18270 856
rect 18438 800 18546 856
rect 18714 800 18914 856
rect 19082 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20754 856
rect 20922 800 21122 856
rect 21290 800 21398 856
rect 21566 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22502 856
rect 22670 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23606 856
rect 23774 800 23974 856
rect 24142 800 24342 856
rect 24510 800 24618 856
rect 24786 800 24986 856
rect 25154 800 25354 856
rect 25522 800 25722 856
rect 25890 800 26090 856
rect 26258 800 26458 856
rect 26626 800 26826 856
rect 26994 800 27194 856
rect 27362 800 27470 856
rect 27638 800 27838 856
rect 28006 800 28206 856
rect 28374 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29310 856
rect 29478 800 29678 856
rect 29846 800 30046 856
rect 30214 800 30414 856
rect 30582 800 30690 856
rect 30858 800 31058 856
rect 31226 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34278 856
rect 34446 800 34646 856
rect 34814 800 35014 856
rect 35182 800 35382 856
rect 35550 800 35750 856
rect 35918 800 36118 856
rect 36286 800 36486 856
rect 36654 800 36762 856
rect 36930 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38234 856
rect 38402 800 38602 856
rect 38770 800 38970 856
rect 39138 800 39338 856
rect 39506 800 39706 856
rect 39874 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42558 856
rect 42726 800 42834 856
rect 43002 800 43202 856
rect 43370 800 43570 856
rect 43738 800 43938 856
rect 44106 800 44306 856
rect 44474 800 44674 856
rect 44842 800 45042 856
rect 45210 800 45410 856
rect 45578 800 45778 856
rect 45946 800 46054 856
rect 46222 800 46422 856
rect 46590 800 46790 856
rect 46958 800 47158 856
rect 47326 800 47526 856
rect 47694 800 47894 856
rect 48062 800 48262 856
rect 48430 800 48630 856
rect 48798 800 48906 856
rect 49074 800 49274 856
rect 49442 800 49642 856
rect 49810 800 50010 856
rect 50178 800 50378 856
rect 50546 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51482 856
rect 51650 800 51850 856
rect 52018 800 52126 856
rect 52294 800 52494 856
rect 52662 800 52862 856
rect 53030 800 53230 856
rect 53398 800 53598 856
rect 53766 800 53966 856
rect 54134 800 54334 856
rect 54502 800 54702 856
rect 54870 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55714 856
rect 55882 800 56082 856
rect 56250 800 56450 856
rect 56618 800 56818 856
rect 56986 800 57186 856
rect 57354 800 57554 856
rect 57722 800 57922 856
rect 58090 800 58198 856
rect 58366 800 58566 856
rect 58734 800 58934 856
rect 59102 800 59302 856
rect 59470 800 59670 856
rect 59838 800 60038 856
rect 60206 800 60406 856
rect 60574 800 60774 856
rect 60942 800 61050 856
rect 61218 800 61418 856
rect 61586 800 61786 856
rect 61954 800 62154 856
rect 62322 800 62522 856
rect 62690 800 62890 856
rect 63058 800 63258 856
rect 63426 800 63626 856
rect 63794 800 63994 856
rect 64162 800 64270 856
rect 64438 800 64638 856
rect 64806 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65742 856
rect 65910 800 66110 856
rect 66278 800 66478 856
rect 66646 800 66846 856
rect 67014 800 67122 856
rect 67290 800 67490 856
rect 67658 800 67858 856
rect 68026 800 68226 856
rect 68394 800 68594 856
rect 68762 800 68962 856
rect 69130 800 69330 856
rect 69498 800 69698 856
rect 69866 800 70066 856
rect 70234 800 70342 856
rect 70510 800 70710 856
rect 70878 800 71078 856
rect 71246 800 71446 856
rect 71614 800 71814 856
rect 71982 800 72182 856
rect 72350 800 72550 856
rect 72718 800 72918 856
rect 73086 800 73286 856
rect 73454 800 73562 856
rect 73730 800 73930 856
rect 74098 800 74298 856
rect 74466 800 74666 856
rect 74834 800 75034 856
rect 75202 800 75402 856
rect 75570 800 75770 856
rect 75938 800 76138 856
rect 76306 800 76414 856
rect 76582 800 76782 856
rect 76950 800 77150 856
rect 77318 800 77518 856
rect 77686 800 77886 856
rect 78054 800 78254 856
rect 78422 800 78622 856
rect 78790 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79634 856
rect 79802 800 80002 856
rect 80170 800 80370 856
rect 80538 800 80738 856
rect 80906 800 81106 856
rect 81274 800 81474 856
rect 81642 800 81842 856
rect 82010 800 82210 856
rect 82378 800 82486 856
rect 82654 800 82854 856
rect 83022 800 83222 856
rect 83390 800 83590 856
rect 83758 800 83958 856
rect 84126 800 84326 856
rect 84494 800 84694 856
rect 84862 800 85062 856
rect 85230 800 85430 856
rect 85598 800 85706 856
rect 85874 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86810 856
rect 86978 800 87178 856
rect 87346 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88282 856
rect 88450 800 88558 856
rect 88726 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89662 856
rect 89830 800 90030 856
rect 90198 800 90398 856
rect 90566 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91502 856
rect 91670 800 91778 856
rect 91946 800 92146 856
rect 92314 800 92514 856
rect 92682 800 92882 856
rect 93050 800 93250 856
rect 93418 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94630 856
rect 94798 800 94998 856
rect 95166 800 95366 856
rect 95534 800 95734 856
rect 95902 800 96102 856
rect 96270 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97206 856
rect 97374 800 97574 856
rect 97742 800 97850 856
rect 98018 800 98218 856
rect 98386 800 98586 856
rect 98754 800 98954 856
rect 99122 800 99322 856
rect 99490 800 99690 856
rect 99858 800 100058 856
rect 100226 800 100426 856
rect 100594 800 100702 856
rect 100870 800 101070 856
rect 101238 800 101438 856
rect 101606 800 101806 856
rect 101974 800 102174 856
rect 102342 800 102542 856
rect 102710 800 102910 856
rect 103078 800 103278 856
rect 103446 800 103646 856
rect 103814 800 103922 856
rect 104090 800 104290 856
rect 104458 800 104658 856
rect 104826 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105762 856
rect 105930 800 106130 856
rect 106298 800 106498 856
rect 106666 800 106774 856
rect 106942 800 107142 856
rect 107310 800 107510 856
rect 107678 800 107878 856
rect 108046 800 108246 856
rect 108414 800 108614 856
rect 108782 800 108982 856
rect 109150 800 109350 856
rect 109518 800 109718 856
rect 109886 800 109994 856
rect 110162 800 110362 856
rect 110530 800 110730 856
rect 110898 800 111098 856
rect 111266 800 111466 856
rect 111634 800 111834 856
rect 112002 800 112202 856
rect 112370 800 112570 856
rect 112738 800 112938 856
rect 113106 800 113214 856
rect 113382 800 113582 856
rect 113750 800 113950 856
rect 114118 800 114318 856
rect 114486 800 114686 856
rect 114854 800 115054 856
rect 115222 800 115422 856
rect 115590 800 115790 856
rect 115958 800 116066 856
rect 116234 800 116434 856
rect 116602 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117538 856
rect 117706 800 117906 856
rect 118074 800 118274 856
rect 118442 800 118642 856
rect 118810 800 119010 856
rect 119178 800 119286 856
rect 119454 800 119654 856
rect 119822 800 120022 856
rect 120190 800 120390 856
rect 120558 800 120758 856
rect 120926 800 121126 856
rect 121294 800 121494 856
rect 121662 800 121862 856
rect 122030 800 122138 856
rect 122306 800 122506 856
rect 122674 800 122874 856
rect 123042 800 123242 856
rect 123410 800 123610 856
rect 123778 800 123978 856
rect 124146 800 124346 856
rect 124514 800 124714 856
rect 124882 800 125082 856
rect 125250 800 125358 856
rect 125526 800 125726 856
rect 125894 800 126094 856
rect 126262 800 126462 856
rect 126630 800 126830 856
rect 126998 800 127198 856
rect 127366 800 127566 856
rect 127734 800 127934 856
rect 128102 800 128210 856
rect 128378 800 128578 856
rect 128746 800 128946 856
rect 129114 800 129314 856
rect 129482 800 129682 856
rect 129850 800 130050 856
rect 130218 800 130418 856
rect 130586 800 130786 856
rect 130954 800 131154 856
rect 131322 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132166 856
rect 132334 800 132534 856
rect 132702 800 132902 856
rect 133070 800 133270 856
rect 133438 800 133638 856
rect 133806 800 134006 856
rect 134174 800 134282 856
rect 134450 800 134650 856
rect 134818 800 135018 856
rect 135186 800 135386 856
rect 135554 800 135754 856
rect 135922 800 136122 856
rect 136290 800 136490 856
rect 136658 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137502 856
rect 137670 800 137870 856
rect 138038 800 138238 856
rect 138406 800 138606 856
rect 138774 800 138974 856
rect 139142 800 139342 856
rect 139510 800 139710 856
rect 139878 800 140078 856
rect 140246 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141090 856
rect 141258 800 141458 856
rect 141626 800 141826 856
rect 141994 800 142194 856
rect 142362 800 142562 856
rect 142730 800 142930 856
rect 143098 800 143298 856
rect 143466 800 143574 856
rect 143742 800 143942 856
rect 144110 800 144310 856
rect 144478 800 144678 856
rect 144846 800 145046 856
rect 145214 800 145414 856
rect 145582 800 145782 856
rect 145950 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146794 856
rect 146962 800 147162 856
rect 147330 800 147530 856
rect 147698 800 147898 856
rect 148066 800 148266 856
rect 148434 800 148634 856
rect 148802 800 149002 856
rect 149170 800 149370 856
rect 149538 800 149646 856
rect 149814 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150750 856
rect 150918 800 151118 856
rect 151286 800 151486 856
rect 151654 800 151854 856
rect 152022 800 152222 856
rect 152390 800 152590 856
rect 152758 800 152866 856
rect 153034 800 153234 856
rect 153402 800 153602 856
rect 153770 800 153970 856
rect 154138 800 154338 856
rect 154506 800 154706 856
rect 154874 800 155074 856
rect 155242 800 155442 856
rect 155610 800 155718 856
rect 155886 800 156086 856
rect 156254 800 156454 856
rect 156622 800 156822 856
rect 156990 800 157190 856
rect 157358 800 157558 856
rect 157726 800 157926 856
rect 158094 800 158294 856
rect 158462 800 158662 856
rect 158830 800 158938 856
rect 159106 800 159306 856
rect 159474 800 159674 856
rect 159842 800 160042 856
rect 160210 800 160410 856
rect 160578 800 160778 856
rect 160946 800 161146 856
rect 161314 800 161514 856
rect 161682 800 161790 856
rect 161958 800 162158 856
rect 162326 800 162526 856
rect 162694 800 162894 856
rect 163062 800 163262 856
rect 163430 800 163630 856
rect 163798 800 163998 856
rect 164166 800 164366 856
rect 164534 800 164734 856
rect 164902 800 165010 856
rect 165178 800 165378 856
rect 165546 800 165746 856
rect 165914 800 166114 856
rect 166282 800 166482 856
rect 166650 800 166850 856
rect 167018 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167862 856
rect 168030 800 168230 856
rect 168398 800 168598 856
rect 168766 800 168966 856
rect 169134 800 169334 856
rect 169502 800 169702 856
rect 169870 800 170070 856
rect 170238 800 170438 856
rect 170606 800 170806 856
rect 170974 800 171082 856
rect 171250 800 171450 856
rect 171618 800 171818 856
rect 171986 800 172186 856
rect 172354 800 172554 856
rect 172722 800 172922 856
rect 173090 800 173290 856
rect 173458 800 173658 856
rect 173826 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175038 856
rect 175206 800 175406 856
rect 175574 800 175774 856
rect 175942 800 176142 856
rect 176310 800 176510 856
rect 176678 800 176878 856
rect 177046 800 177154 856
rect 177322 800 177522 856
rect 177690 800 177890 856
rect 178058 800 178186 856
<< metal3 >>
rect 0 111392 800 111512
rect 179200 107856 180000 107976
rect 0 94256 800 94376
rect 179200 83920 180000 84040
rect 0 77120 800 77240
rect 0 59984 800 60104
rect 179200 59848 180000 59968
rect 0 42848 800 42968
rect 179200 35912 180000 36032
rect 0 25712 800 25832
rect 179200 11976 180000 12096
rect 0 8576 800 8696
<< obsm3 >>
rect 800 111592 179200 117741
rect 880 111312 179200 111592
rect 800 108056 179200 111312
rect 800 107776 179120 108056
rect 800 94456 179200 107776
rect 880 94176 179200 94456
rect 800 84120 179200 94176
rect 800 83840 179120 84120
rect 800 77320 179200 83840
rect 880 77040 179200 77320
rect 800 60184 179200 77040
rect 880 60048 179200 60184
rect 880 59904 179120 60048
rect 800 59768 179120 59904
rect 800 43048 179200 59768
rect 880 42768 179200 43048
rect 800 36112 179200 42768
rect 800 35832 179120 36112
rect 800 25912 179200 35832
rect 880 25632 179200 25912
rect 800 12176 179200 25632
rect 800 11896 179120 12176
rect 800 8776 179200 11896
rect 880 8496 179200 8776
rect 800 2143 179200 8496
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 88195 6155 96288 117469
rect 96768 6155 96909 117469
<< labels >>
rlabel metal2 s 175094 0 175150 800 6 active
port 1 nsew signal input
rlabel metal2 s 168930 119200 168986 120000 6 analog_io[0]
port 2 nsew signal bidirectional
rlabel metal3 s 0 42848 800 42968 6 analog_io[10]
port 3 nsew signal bidirectional
rlabel metal2 s 177946 0 178002 800 6 analog_io[11]
port 4 nsew signal bidirectional
rlabel metal3 s 0 59984 800 60104 6 analog_io[12]
port 5 nsew signal bidirectional
rlabel metal2 s 173346 119200 173402 120000 6 analog_io[13]
port 6 nsew signal bidirectional
rlabel metal2 s 174818 119200 174874 120000 6 analog_io[14]
port 7 nsew signal bidirectional
rlabel metal2 s 178314 0 178370 800 6 analog_io[15]
port 8 nsew signal bidirectional
rlabel metal2 s 176290 119200 176346 120000 6 analog_io[16]
port 9 nsew signal bidirectional
rlabel metal2 s 178682 0 178738 800 6 analog_io[17]
port 10 nsew signal bidirectional
rlabel metal3 s 0 77120 800 77240 6 analog_io[18]
port 11 nsew signal bidirectional
rlabel metal3 s 0 94256 800 94376 6 analog_io[19]
port 12 nsew signal bidirectional
rlabel metal2 s 175462 0 175518 800 6 analog_io[1]
port 13 nsew signal bidirectional
rlabel metal2 s 179050 0 179106 800 6 analog_io[20]
port 14 nsew signal bidirectional
rlabel metal2 s 177762 119200 177818 120000 6 analog_io[21]
port 15 nsew signal bidirectional
rlabel metal3 s 179200 59848 180000 59968 6 analog_io[22]
port 16 nsew signal bidirectional
rlabel metal3 s 0 111392 800 111512 6 analog_io[23]
port 17 nsew signal bidirectional
rlabel metal2 s 179418 0 179474 800 6 analog_io[24]
port 18 nsew signal bidirectional
rlabel metal2 s 179234 119200 179290 120000 6 analog_io[25]
port 19 nsew signal bidirectional
rlabel metal3 s 179200 83920 180000 84040 6 analog_io[26]
port 20 nsew signal bidirectional
rlabel metal2 s 179786 0 179842 800 6 analog_io[27]
port 21 nsew signal bidirectional
rlabel metal3 s 179200 107856 180000 107976 6 analog_io[28]
port 22 nsew signal bidirectional
rlabel metal2 s 176198 0 176254 800 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 170402 119200 170458 120000 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal2 s 171874 119200 171930 120000 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal2 s 176566 0 176622 800 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal2 s 176934 0 176990 800 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal2 s 177210 0 177266 800 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 0 25712 800 25832 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal2 s 177578 0 177634 800 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 31 nsew signal input
rlabel metal2 s 45006 119200 45062 120000 6 io_in[10]
port 32 nsew signal input
rlabel metal2 s 49422 119200 49478 120000 6 io_in[11]
port 33 nsew signal input
rlabel metal2 s 53838 119200 53894 120000 6 io_in[12]
port 34 nsew signal input
rlabel metal2 s 58254 119200 58310 120000 6 io_in[13]
port 35 nsew signal input
rlabel metal2 s 62670 119200 62726 120000 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 67086 119200 67142 120000 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 71502 119200 71558 120000 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 76010 119200 76066 120000 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 80426 119200 80482 120000 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 84842 119200 84898 120000 6 io_in[19]
port 41 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 89258 119200 89314 120000 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 93674 119200 93730 120000 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 98090 119200 98146 120000 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 102506 119200 102562 120000 6 io_in[23]
port 46 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 io_in[24]
port 47 nsew signal input
rlabel metal2 s 111430 119200 111486 120000 6 io_in[25]
port 48 nsew signal input
rlabel metal2 s 115846 119200 115902 120000 6 io_in[26]
port 49 nsew signal input
rlabel metal2 s 120262 119200 120318 120000 6 io_in[27]
port 50 nsew signal input
rlabel metal2 s 124678 119200 124734 120000 6 io_in[28]
port 51 nsew signal input
rlabel metal2 s 129094 119200 129150 120000 6 io_in[29]
port 52 nsew signal input
rlabel metal2 s 9586 119200 9642 120000 6 io_in[2]
port 53 nsew signal input
rlabel metal2 s 133510 119200 133566 120000 6 io_in[30]
port 54 nsew signal input
rlabel metal2 s 137926 119200 137982 120000 6 io_in[31]
port 55 nsew signal input
rlabel metal2 s 142342 119200 142398 120000 6 io_in[32]
port 56 nsew signal input
rlabel metal2 s 146850 119200 146906 120000 6 io_in[33]
port 57 nsew signal input
rlabel metal2 s 151266 119200 151322 120000 6 io_in[34]
port 58 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[35]
port 59 nsew signal input
rlabel metal2 s 160098 119200 160154 120000 6 io_in[36]
port 60 nsew signal input
rlabel metal2 s 164514 119200 164570 120000 6 io_in[37]
port 61 nsew signal input
rlabel metal2 s 14002 119200 14058 120000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 18418 119200 18474 120000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 22834 119200 22890 120000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 27250 119200 27306 120000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 31666 119200 31722 120000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 40590 119200 40646 120000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 46478 119200 46534 120000 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 50894 119200 50950 120000 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 55310 119200 55366 120000 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 59726 119200 59782 120000 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 68558 119200 68614 120000 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 73066 119200 73122 120000 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 77482 119200 77538 120000 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 81898 119200 81954 120000 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 86314 119200 86370 120000 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 90730 119200 90786 120000 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 95146 119200 95202 120000 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 99562 119200 99618 120000 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 103978 119200 104034 120000 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 108394 119200 108450 120000 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 112902 119200 112958 120000 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 117318 119200 117374 120000 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 121734 119200 121790 120000 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 126150 119200 126206 120000 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 130566 119200 130622 120000 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 11058 119200 11114 120000 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 139398 119200 139454 120000 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 143814 119200 143870 120000 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 148322 119200 148378 120000 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 152738 119200 152794 120000 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 161570 119200 161626 120000 6 io_oeb[36]
port 98 nsew signal output
rlabel metal2 s 165986 119200 166042 120000 6 io_oeb[37]
port 99 nsew signal output
rlabel metal2 s 15474 119200 15530 120000 6 io_oeb[3]
port 100 nsew signal output
rlabel metal2 s 19890 119200 19946 120000 6 io_oeb[4]
port 101 nsew signal output
rlabel metal2 s 24306 119200 24362 120000 6 io_oeb[5]
port 102 nsew signal output
rlabel metal2 s 28722 119200 28778 120000 6 io_oeb[6]
port 103 nsew signal output
rlabel metal2 s 33138 119200 33194 120000 6 io_oeb[7]
port 104 nsew signal output
rlabel metal2 s 37646 119200 37702 120000 6 io_oeb[8]
port 105 nsew signal output
rlabel metal2 s 42062 119200 42118 120000 6 io_oeb[9]
port 106 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 107 nsew signal output
rlabel metal2 s 47950 119200 48006 120000 6 io_out[10]
port 108 nsew signal output
rlabel metal2 s 52366 119200 52422 120000 6 io_out[11]
port 109 nsew signal output
rlabel metal2 s 56782 119200 56838 120000 6 io_out[12]
port 110 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 io_out[13]
port 111 nsew signal output
rlabel metal2 s 65614 119200 65670 120000 6 io_out[14]
port 112 nsew signal output
rlabel metal2 s 70030 119200 70086 120000 6 io_out[15]
port 113 nsew signal output
rlabel metal2 s 74538 119200 74594 120000 6 io_out[16]
port 114 nsew signal output
rlabel metal2 s 78954 119200 79010 120000 6 io_out[17]
port 115 nsew signal output
rlabel metal2 s 83370 119200 83426 120000 6 io_out[18]
port 116 nsew signal output
rlabel metal2 s 87786 119200 87842 120000 6 io_out[19]
port 117 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 118 nsew signal output
rlabel metal2 s 92202 119200 92258 120000 6 io_out[20]
port 119 nsew signal output
rlabel metal2 s 96618 119200 96674 120000 6 io_out[21]
port 120 nsew signal output
rlabel metal2 s 101034 119200 101090 120000 6 io_out[22]
port 121 nsew signal output
rlabel metal2 s 105450 119200 105506 120000 6 io_out[23]
port 122 nsew signal output
rlabel metal2 s 109958 119200 110014 120000 6 io_out[24]
port 123 nsew signal output
rlabel metal2 s 114374 119200 114430 120000 6 io_out[25]
port 124 nsew signal output
rlabel metal2 s 118790 119200 118846 120000 6 io_out[26]
port 125 nsew signal output
rlabel metal2 s 123206 119200 123262 120000 6 io_out[27]
port 126 nsew signal output
rlabel metal2 s 127622 119200 127678 120000 6 io_out[28]
port 127 nsew signal output
rlabel metal2 s 132038 119200 132094 120000 6 io_out[29]
port 128 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_out[2]
port 129 nsew signal output
rlabel metal2 s 136454 119200 136510 120000 6 io_out[30]
port 130 nsew signal output
rlabel metal2 s 140870 119200 140926 120000 6 io_out[31]
port 131 nsew signal output
rlabel metal2 s 145378 119200 145434 120000 6 io_out[32]
port 132 nsew signal output
rlabel metal2 s 149794 119200 149850 120000 6 io_out[33]
port 133 nsew signal output
rlabel metal2 s 154210 119200 154266 120000 6 io_out[34]
port 134 nsew signal output
rlabel metal2 s 158626 119200 158682 120000 6 io_out[35]
port 135 nsew signal output
rlabel metal2 s 163042 119200 163098 120000 6 io_out[36]
port 136 nsew signal output
rlabel metal2 s 167458 119200 167514 120000 6 io_out[37]
port 137 nsew signal output
rlabel metal2 s 16946 119200 17002 120000 6 io_out[3]
port 138 nsew signal output
rlabel metal2 s 21362 119200 21418 120000 6 io_out[4]
port 139 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_out[5]
port 140 nsew signal output
rlabel metal2 s 30194 119200 30250 120000 6 io_out[6]
port 141 nsew signal output
rlabel metal2 s 34610 119200 34666 120000 6 io_out[7]
port 142 nsew signal output
rlabel metal2 s 39118 119200 39174 120000 6 io_out[8]
port 143 nsew signal output
rlabel metal2 s 43534 119200 43590 120000 6 io_out[9]
port 144 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_data_out[0]
port 273 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[100]
port 274 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[101]
port 275 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[102]
port 276 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[103]
port 277 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[104]
port 278 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 la_data_out[105]
port 279 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 la_data_out[106]
port 280 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[107]
port 281 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 la_data_out[108]
port 282 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[109]
port 283 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[10]
port 284 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[110]
port 285 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[111]
port 286 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 la_data_out[112]
port 287 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[113]
port 288 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[114]
port 289 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 la_data_out[115]
port 290 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[116]
port 291 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[117]
port 292 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[118]
port 293 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[119]
port 294 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[11]
port 295 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[120]
port 296 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 la_data_out[121]
port 297 nsew signal output
rlabel metal2 s 169022 0 169078 800 6 la_data_out[122]
port 298 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[123]
port 299 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[124]
port 300 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 la_data_out[125]
port 301 nsew signal output
rlabel metal2 s 173346 0 173402 800 6 la_data_out[126]
port 302 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[127]
port 303 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[12]
port 304 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[13]
port 305 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[14]
port 306 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[15]
port 307 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[16]
port 308 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 la_data_out[17]
port 309 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[18]
port 310 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[19]
port 311 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 la_data_out[1]
port 312 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 la_data_out[20]
port 313 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[21]
port 314 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[22]
port 315 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[23]
port 316 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[24]
port 317 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[25]
port 318 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[26]
port 319 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[27]
port 320 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[28]
port 321 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[29]
port 322 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[2]
port 323 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[30]
port 324 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[31]
port 325 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[32]
port 326 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 la_data_out[33]
port 327 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[34]
port 328 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 la_data_out[35]
port 329 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[36]
port 330 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[37]
port 331 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[38]
port 332 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[39]
port 333 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[3]
port 334 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[40]
port 335 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[41]
port 336 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[42]
port 337 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[43]
port 338 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[44]
port 339 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[45]
port 340 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[46]
port 341 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 la_data_out[47]
port 342 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[48]
port 343 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[49]
port 344 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[4]
port 345 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[50]
port 346 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[51]
port 347 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[52]
port 348 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[53]
port 349 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[54]
port 350 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[55]
port 351 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[56]
port 352 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[57]
port 353 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[58]
port 354 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 la_data_out[59]
port 355 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[5]
port 356 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[60]
port 357 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[61]
port 358 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[62]
port 359 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[63]
port 360 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[64]
port 361 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[65]
port 362 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[66]
port 363 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[67]
port 364 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[68]
port 365 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[69]
port 366 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[6]
port 367 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[70]
port 368 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[71]
port 369 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 la_data_out[72]
port 370 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[73]
port 371 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 la_data_out[74]
port 372 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[75]
port 373 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[76]
port 374 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_out[77]
port 375 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_out[78]
port 376 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[79]
port 377 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 la_data_out[7]
port 378 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[80]
port 379 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[81]
port 380 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[82]
port 381 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[83]
port 382 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[84]
port 383 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[85]
port 384 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[86]
port 385 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[87]
port 386 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 la_data_out[88]
port 387 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[89]
port 388 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[8]
port 389 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[90]
port 390 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[91]
port 391 nsew signal output
rlabel metal2 s 136914 0 136970 800 6 la_data_out[92]
port 392 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 la_data_out[93]
port 393 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[94]
port 394 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[95]
port 395 nsew signal output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[96]
port 396 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 la_data_out[97]
port 397 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[98]
port 398 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 la_data_out[99]
port 399 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[9]
port 400 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_oenb[0]
port 401 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[100]
port 402 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[101]
port 403 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[102]
port 404 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[103]
port 405 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 la_oenb[104]
port 406 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[105]
port 407 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_oenb[106]
port 408 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[107]
port 409 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[108]
port 410 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_oenb[109]
port 411 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[10]
port 412 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_oenb[110]
port 413 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 la_oenb[111]
port 414 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[112]
port 415 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[113]
port 416 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[114]
port 417 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_oenb[115]
port 418 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_oenb[116]
port 419 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[117]
port 420 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[118]
port 421 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oenb[119]
port 422 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[11]
port 423 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oenb[120]
port 424 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oenb[121]
port 425 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 la_oenb[122]
port 426 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_oenb[123]
port 427 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_oenb[124]
port 428 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_oenb[125]
port 429 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_oenb[126]
port 430 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_oenb[127]
port 431 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_oenb[12]
port 432 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[13]
port 433 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[14]
port 434 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[15]
port 435 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[16]
port 436 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[17]
port 437 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[18]
port 438 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[19]
port 439 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_oenb[1]
port 440 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_oenb[20]
port 441 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[21]
port 442 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[22]
port 443 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[23]
port 444 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[24]
port 445 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[25]
port 446 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[26]
port 447 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_oenb[27]
port 448 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[28]
port 449 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[29]
port 450 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_oenb[2]
port 451 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[30]
port 452 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[31]
port 453 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[32]
port 454 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_oenb[33]
port 455 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_oenb[34]
port 456 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[35]
port 457 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_oenb[36]
port 458 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_oenb[37]
port 459 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oenb[38]
port 460 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 la_oenb[39]
port 461 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[3]
port 462 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 la_oenb[40]
port 463 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[41]
port 464 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[42]
port 465 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[43]
port 466 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[44]
port 467 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[45]
port 468 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[46]
port 469 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[47]
port 470 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[48]
port 471 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[49]
port 472 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[4]
port 473 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[50]
port 474 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[51]
port 475 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[52]
port 476 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[53]
port 477 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[54]
port 478 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[55]
port 479 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[56]
port 480 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[57]
port 481 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[58]
port 482 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[59]
port 483 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 la_oenb[5]
port 484 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_oenb[60]
port 485 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[61]
port 486 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[62]
port 487 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[63]
port 488 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[64]
port 489 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_oenb[65]
port 490 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[66]
port 491 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[67]
port 492 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[68]
port 493 nsew signal input
rlabel metal2 s 112626 0 112682 800 6 la_oenb[69]
port 494 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[6]
port 495 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[70]
port 496 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[71]
port 497 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_oenb[72]
port 498 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[73]
port 499 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_oenb[74]
port 500 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[75]
port 501 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[76]
port 502 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_oenb[77]
port 503 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[78]
port 504 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[79]
port 505 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[7]
port 506 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[80]
port 507 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[81]
port 508 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_oenb[82]
port 509 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oenb[83]
port 510 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[84]
port 511 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[85]
port 512 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_oenb[86]
port 513 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[87]
port 514 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[88]
port 515 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[89]
port 516 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_oenb[8]
port 517 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[90]
port 518 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[91]
port 519 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[92]
port 520 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[93]
port 521 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[94]
port 522 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[95]
port 523 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[96]
port 524 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[97]
port 525 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[98]
port 526 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[99]
port 527 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[9]
port 528 nsew signal input
rlabel metal3 s 179200 11976 180000 12096 6 user_clock2
port 529 nsew signal input
rlabel metal3 s 179200 35912 180000 36032 6 user_irq[0]
port 530 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 user_irq[1]
port 531 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 user_irq[2]
port 532 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 533 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 534 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 534 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 535 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 537 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[0]
port 538 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[10]
port 539 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[11]
port 540 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[12]
port 541 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[13]
port 542 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[14]
port 543 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[15]
port 544 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[16]
port 545 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[17]
port 546 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[18]
port 547 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_adr_i[19]
port 548 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_adr_i[1]
port 549 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[20]
port 550 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[21]
port 551 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[22]
port 552 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[23]
port 553 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_adr_i[24]
port 554 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_adr_i[25]
port 555 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[26]
port 556 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[27]
port 557 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[28]
port 558 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[29]
port 559 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[2]
port 560 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[30]
port 561 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_adr_i[31]
port 562 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[3]
port 563 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_adr_i[4]
port 564 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[5]
port 565 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[6]
port 566 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[7]
port 567 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[8]
port 568 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[9]
port 569 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_cyc_i
port 570 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[0]
port 571 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[10]
port 572 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[11]
port 573 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[12]
port 574 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[13]
port 575 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[14]
port 576 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_i[15]
port 577 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[16]
port 578 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[17]
port 579 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[18]
port 580 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[19]
port 581 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_i[1]
port 582 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[20]
port 583 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[21]
port 584 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[22]
port 585 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[23]
port 586 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[24]
port 587 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_i[25]
port 588 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[26]
port 589 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[27]
port 590 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[28]
port 591 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[29]
port 592 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_dat_i[2]
port 593 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[30]
port 594 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[31]
port 595 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_i[3]
port 596 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_i[4]
port 597 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[5]
port 598 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[6]
port 599 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[7]
port 600 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[8]
port 601 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[9]
port 602 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_o[0]
port 603 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_o[10]
port 604 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[11]
port 605 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[12]
port 606 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[13]
port 607 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[14]
port 608 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_o[15]
port 609 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[16]
port 610 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[17]
port 611 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[18]
port 612 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[19]
port 613 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[1]
port 614 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[20]
port 615 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[21]
port 616 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[22]
port 617 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_o[23]
port 618 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[24]
port 619 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[25]
port 620 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[26]
port 621 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[27]
port 622 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[28]
port 623 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[29]
port 624 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[2]
port 625 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_o[30]
port 626 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[31]
port 627 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[3]
port 628 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[4]
port 629 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[5]
port 630 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[6]
port 631 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[7]
port 632 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[8]
port 633 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_o[9]
port 634 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_sel_i[0]
port 635 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[1]
port 636 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[2]
port 637 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_sel_i[3]
port 638 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_stb_i
port 639 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_we_i
port 640 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7790302
string GDS_FILE /opt/mpw6/sel_set/openlane/user_proj_example/runs/user_proj_example/results/finishing/macro_la.magic.gds
string GDS_START 294060
<< end >>

