VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1115.570 1421.780 1115.890 1421.840 ;
        RECT 2900.830 1421.780 2901.150 1421.840 ;
        RECT 1115.570 1421.640 2901.150 1421.780 ;
        RECT 1115.570 1421.580 1115.890 1421.640 ;
        RECT 2900.830 1421.580 2901.150 1421.640 ;
      LAYER via ;
        RECT 1115.600 1421.580 1115.860 1421.840 ;
        RECT 2900.860 1421.580 2901.120 1421.840 ;
      LAYER met2 ;
        RECT 2900.850 1426.795 2901.130 1427.165 ;
        RECT 2900.920 1421.870 2901.060 1426.795 ;
        RECT 1115.600 1421.550 1115.860 1421.870 ;
        RECT 2900.860 1421.550 2901.120 1421.870 ;
        RECT 1115.660 424.165 1115.800 1421.550 ;
        RECT 1115.590 423.795 1115.870 424.165 ;
      LAYER via2 ;
        RECT 2900.850 1426.840 2901.130 1427.120 ;
        RECT 1115.590 423.840 1115.870 424.120 ;
      LAYER met3 ;
        RECT 2900.825 1427.130 2901.155 1427.145 ;
        RECT 2917.600 1427.130 2924.800 1427.580 ;
        RECT 2900.825 1426.830 2924.800 1427.130 ;
        RECT 2900.825 1426.815 2901.155 1426.830 ;
        RECT 2917.600 1426.380 2924.800 1426.830 ;
        RECT 1115.565 424.130 1115.895 424.145 ;
        RECT 1098.790 423.830 1115.895 424.130 ;
        RECT 1098.790 421.720 1099.090 423.830 ;
        RECT 1115.565 423.815 1115.895 423.830 ;
        RECT 1096.000 421.120 1100.000 421.720 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 682.960 1117.730 683.020 ;
        RECT 2228.770 682.960 2229.090 683.020 ;
        RECT 1117.410 682.820 2229.090 682.960 ;
        RECT 1117.410 682.760 1117.730 682.820 ;
        RECT 2228.770 682.760 2229.090 682.820 ;
      LAYER via ;
        RECT 1117.440 682.760 1117.700 683.020 ;
        RECT 2228.800 682.760 2229.060 683.020 ;
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
        RECT 2230.700 3512.170 2230.840 3517.600 ;
        RECT 2228.860 3512.030 2230.840 3512.170 ;
        RECT 2228.860 683.050 2229.000 3512.030 ;
        RECT 1117.440 682.730 1117.700 683.050 ;
        RECT 2228.800 682.730 2229.060 683.050 ;
        RECT 1117.500 680.525 1117.640 682.730 ;
        RECT 1117.430 680.155 1117.710 680.525 ;
      LAYER via2 ;
        RECT 1117.430 680.200 1117.710 680.480 ;
      LAYER met3 ;
        RECT 1117.405 680.490 1117.735 680.505 ;
        RECT 1098.790 680.190 1117.735 680.490 ;
        RECT 1098.790 678.760 1099.090 680.190 ;
        RECT 1117.405 680.175 1117.735 680.190 ;
        RECT 1096.000 678.160 1100.000 678.760 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 724.440 1117.730 724.500 ;
        RECT 1904.470 724.440 1904.790 724.500 ;
        RECT 1117.410 724.300 1904.790 724.440 ;
        RECT 1117.410 724.240 1117.730 724.300 ;
        RECT 1904.470 724.240 1904.790 724.300 ;
      LAYER via ;
        RECT 1117.440 724.240 1117.700 724.500 ;
        RECT 1904.500 724.240 1904.760 724.500 ;
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
        RECT 1905.940 3512.170 1906.080 3517.600 ;
        RECT 1904.560 3512.030 1906.080 3512.170 ;
        RECT 1904.560 724.530 1904.700 3512.030 ;
        RECT 1117.440 724.210 1117.700 724.530 ;
        RECT 1904.500 724.210 1904.760 724.530 ;
        RECT 1117.500 722.685 1117.640 724.210 ;
        RECT 1117.430 722.315 1117.710 722.685 ;
      LAYER via2 ;
        RECT 1117.430 722.360 1117.710 722.640 ;
      LAYER met3 ;
        RECT 1117.405 722.650 1117.735 722.665 ;
        RECT 1098.790 722.350 1117.735 722.650 ;
        RECT 1098.790 721.600 1099.090 722.350 ;
        RECT 1117.405 722.335 1117.735 722.350 ;
        RECT 1096.000 721.000 1100.000 721.600 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 191.430 1004.260 191.750 1004.320 ;
        RECT 1580.170 1004.260 1580.490 1004.320 ;
        RECT 191.430 1004.120 1580.490 1004.260 ;
        RECT 191.430 1004.060 191.750 1004.120 ;
        RECT 1580.170 1004.060 1580.490 1004.120 ;
      LAYER via ;
        RECT 191.460 1004.060 191.720 1004.320 ;
        RECT 1580.200 1004.060 1580.460 1004.320 ;
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
        RECT 1581.640 3512.170 1581.780 3517.600 ;
        RECT 1580.260 3512.030 1581.780 3512.170 ;
        RECT 1580.260 1004.350 1580.400 3512.030 ;
        RECT 191.460 1004.030 191.720 1004.350 ;
        RECT 1580.200 1004.030 1580.460 1004.350 ;
        RECT 191.520 702.965 191.660 1004.030 ;
        RECT 191.450 702.595 191.730 702.965 ;
      LAYER via2 ;
        RECT 191.450 702.640 191.730 702.920 ;
      LAYER met3 ;
        RECT 191.425 702.930 191.755 702.945 ;
        RECT 191.425 702.630 201.170 702.930 ;
        RECT 191.425 702.615 191.755 702.630 ;
        RECT 200.870 700.520 201.170 702.630 ;
        RECT 200.000 699.920 204.000 700.520 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 765.580 1117.730 765.640 ;
        RECT 1255.870 765.580 1256.190 765.640 ;
        RECT 1117.410 765.440 1256.190 765.580 ;
        RECT 1117.410 765.380 1117.730 765.440 ;
        RECT 1255.870 765.380 1256.190 765.440 ;
      LAYER via ;
        RECT 1117.440 765.380 1117.700 765.640 ;
        RECT 1255.900 765.380 1256.160 765.640 ;
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
        RECT 1257.340 3512.170 1257.480 3517.600 ;
        RECT 1255.960 3512.030 1257.480 3512.170 ;
        RECT 1255.960 765.670 1256.100 3512.030 ;
        RECT 1117.440 765.525 1117.700 765.670 ;
        RECT 1117.430 765.155 1117.710 765.525 ;
        RECT 1255.900 765.350 1256.160 765.670 ;
      LAYER via2 ;
        RECT 1117.430 765.200 1117.710 765.480 ;
      LAYER met3 ;
        RECT 1117.405 765.490 1117.735 765.505 ;
        RECT 1097.870 765.190 1117.735 765.490 ;
        RECT 1097.870 764.440 1098.170 765.190 ;
        RECT 1117.405 765.175 1117.735 765.190 ;
        RECT 1096.000 763.840 1100.000 764.440 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 2784.500 931.890 2784.560 ;
        RECT 1053.470 2784.500 1053.790 2784.560 ;
        RECT 931.570 2784.360 1053.790 2784.500 ;
        RECT 931.570 2784.300 931.890 2784.360 ;
        RECT 1053.470 2784.300 1053.790 2784.360 ;
        RECT 1053.470 1014.120 1053.790 1014.180 ;
        RECT 1080.150 1014.120 1080.470 1014.180 ;
        RECT 1053.470 1013.980 1080.470 1014.120 ;
        RECT 1053.470 1013.920 1053.790 1013.980 ;
        RECT 1080.150 1013.920 1080.470 1013.980 ;
      LAYER via ;
        RECT 931.600 2784.300 931.860 2784.560 ;
        RECT 1053.500 2784.300 1053.760 2784.560 ;
        RECT 1053.500 1013.920 1053.760 1014.180 ;
        RECT 1080.180 1013.920 1080.440 1014.180 ;
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
        RECT 932.580 3415.570 932.720 3517.600 ;
        RECT 931.660 3415.430 932.720 3415.570 ;
        RECT 931.660 2784.590 931.800 3415.430 ;
        RECT 931.600 2784.270 931.860 2784.590 ;
        RECT 1053.500 2784.270 1053.760 2784.590 ;
        RECT 1053.560 1014.210 1053.700 2784.270 ;
        RECT 1053.500 1013.890 1053.760 1014.210 ;
        RECT 1080.180 1013.890 1080.440 1014.210 ;
        RECT 1080.240 999.330 1080.380 1013.890 ;
        RECT 1081.450 999.330 1081.730 1000.000 ;
        RECT 1080.240 999.190 1081.730 999.330 ;
        RECT 1081.450 996.000 1081.730 999.190 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.270 1005.280 607.590 1005.340 ;
        RECT 1110.970 1005.280 1111.290 1005.340 ;
        RECT 607.270 1005.140 1111.290 1005.280 ;
        RECT 607.270 1005.080 607.590 1005.140 ;
        RECT 1110.970 1005.080 1111.290 1005.140 ;
      LAYER via ;
        RECT 607.300 1005.080 607.560 1005.340 ;
        RECT 1111.000 1005.080 1111.260 1005.340 ;
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
        RECT 608.280 3512.170 608.420 3517.600 ;
        RECT 607.360 3512.030 608.420 3512.170 ;
        RECT 607.360 1005.370 607.500 3512.030 ;
        RECT 607.300 1005.050 607.560 1005.370 ;
        RECT 1111.000 1005.050 1111.260 1005.370 ;
        RECT 1111.060 806.325 1111.200 1005.050 ;
        RECT 1110.990 805.955 1111.270 806.325 ;
      LAYER via2 ;
        RECT 1110.990 806.000 1111.270 806.280 ;
      LAYER met3 ;
        RECT 1096.000 806.680 1100.000 807.280 ;
        RECT 1098.790 806.290 1099.090 806.680 ;
        RECT 1110.965 806.290 1111.295 806.305 ;
        RECT 1098.790 805.990 1111.295 806.290 ;
        RECT 1110.965 805.975 1111.295 805.990 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.970 2784.160 283.290 2784.220 ;
        RECT 1053.010 2784.160 1053.330 2784.220 ;
        RECT 282.970 2784.020 1053.330 2784.160 ;
        RECT 282.970 2783.960 283.290 2784.020 ;
        RECT 1053.010 2783.960 1053.330 2784.020 ;
        RECT 1053.010 1013.780 1053.330 1013.840 ;
        RECT 1087.510 1013.780 1087.830 1013.840 ;
        RECT 1053.010 1013.640 1087.830 1013.780 ;
        RECT 1053.010 1013.580 1053.330 1013.640 ;
        RECT 1087.510 1013.580 1087.830 1013.640 ;
      LAYER via ;
        RECT 283.000 2783.960 283.260 2784.220 ;
        RECT 1053.040 2783.960 1053.300 2784.220 ;
        RECT 1053.040 1013.580 1053.300 1013.840 ;
        RECT 1087.540 1013.580 1087.800 1013.840 ;
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
        RECT 283.980 3415.570 284.120 3517.600 ;
        RECT 283.060 3415.430 284.120 3415.570 ;
        RECT 283.060 2784.250 283.200 3415.430 ;
        RECT 283.000 2783.930 283.260 2784.250 ;
        RECT 1053.040 2783.930 1053.300 2784.250 ;
        RECT 1053.100 1013.870 1053.240 2783.930 ;
        RECT 1053.040 1013.550 1053.300 1013.870 ;
        RECT 1087.540 1013.550 1087.800 1013.870 ;
        RECT 1087.600 999.330 1087.740 1013.550 ;
        RECT 1088.810 999.330 1089.090 1000.000 ;
        RECT 1087.600 999.190 1089.090 999.330 ;
        RECT 1088.810 996.000 1089.090 999.190 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.090 786.660 17.410 786.720 ;
        RECT 190.050 786.660 190.370 786.720 ;
        RECT 17.090 786.520 190.370 786.660 ;
        RECT 17.090 786.460 17.410 786.520 ;
        RECT 190.050 786.460 190.370 786.520 ;
      LAYER via ;
        RECT 17.120 786.460 17.380 786.720 ;
        RECT 190.080 786.460 190.340 786.720 ;
      LAYER met2 ;
        RECT 17.110 3486.515 17.390 3486.885 ;
        RECT 17.180 786.750 17.320 3486.515 ;
        RECT 17.120 786.430 17.380 786.750 ;
        RECT 190.080 786.430 190.340 786.750 ;
        RECT 190.140 785.245 190.280 786.430 ;
        RECT 190.070 784.875 190.350 785.245 ;
      LAYER via2 ;
        RECT 17.110 3486.560 17.390 3486.840 ;
        RECT 190.070 784.920 190.350 785.200 ;
      LAYER met3 ;
        RECT -4.800 3486.850 2.400 3487.300 ;
        RECT 17.085 3486.850 17.415 3486.865 ;
        RECT -4.800 3486.550 17.415 3486.850 ;
        RECT -4.800 3486.100 2.400 3486.550 ;
        RECT 17.085 3486.535 17.415 3486.550 ;
        RECT 200.000 785.600 204.000 786.200 ;
        RECT 190.045 785.210 190.375 785.225 ;
        RECT 200.870 785.210 201.170 785.600 ;
        RECT 190.045 784.910 201.170 785.210 ;
        RECT 190.045 784.895 190.375 784.910 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.410 400.180 1093.690 404.000 ;
        RECT 1093.410 400.000 1093.720 400.180 ;
        RECT 1093.580 393.565 1093.720 400.000 ;
        RECT 1093.510 393.195 1093.790 393.565 ;
      LAYER via2 ;
        RECT 1093.510 393.240 1093.790 393.520 ;
      LAYER met3 ;
        RECT -4.800 3225.730 2.400 3226.180 ;
        RECT 16.830 3225.730 17.210 3225.740 ;
        RECT -4.800 3225.430 17.210 3225.730 ;
        RECT -4.800 3224.980 2.400 3225.430 ;
        RECT 16.830 3225.420 17.210 3225.430 ;
        RECT 16.830 393.530 17.210 393.540 ;
        RECT 1093.485 393.530 1093.815 393.545 ;
        RECT 16.830 393.230 1093.815 393.530 ;
        RECT 16.830 393.220 17.210 393.230 ;
        RECT 1093.485 393.215 1093.815 393.230 ;
      LAYER via3 ;
        RECT 16.860 3225.420 17.180 3225.740 ;
        RECT 16.860 393.220 17.180 393.540 ;
      LAYER met4 ;
        RECT 16.855 3225.415 17.185 3225.745 ;
        RECT 16.870 393.545 17.170 3225.415 ;
        RECT 16.855 393.215 17.185 393.545 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2960.280 16.030 2960.340 ;
        RECT 1097.170 2960.280 1097.490 2960.340 ;
        RECT 15.710 2960.140 1097.490 2960.280 ;
        RECT 15.710 2960.080 16.030 2960.140 ;
        RECT 1097.170 2960.080 1097.490 2960.140 ;
      LAYER via ;
        RECT 15.740 2960.080 16.000 2960.340 ;
        RECT 1097.200 2960.080 1097.460 2960.340 ;
      LAYER met2 ;
        RECT 15.730 2964.955 16.010 2965.325 ;
        RECT 15.800 2960.370 15.940 2964.955 ;
        RECT 15.740 2960.050 16.000 2960.370 ;
        RECT 1097.200 2960.050 1097.460 2960.370 ;
        RECT 1097.260 852.565 1097.400 2960.050 ;
        RECT 1097.190 852.195 1097.470 852.565 ;
      LAYER via2 ;
        RECT 15.730 2965.000 16.010 2965.280 ;
        RECT 1097.190 852.240 1097.470 852.520 ;
      LAYER met3 ;
        RECT -4.800 2965.290 2.400 2965.740 ;
        RECT 15.705 2965.290 16.035 2965.305 ;
        RECT -4.800 2964.990 16.035 2965.290 ;
        RECT -4.800 2964.540 2.400 2964.990 ;
        RECT 15.705 2964.975 16.035 2964.990 ;
        RECT 1097.165 852.530 1097.495 852.545 ;
        RECT 1096.950 852.215 1097.495 852.530 ;
        RECT 1096.950 850.120 1097.250 852.215 ;
        RECT 1096.000 849.520 1100.000 850.120 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1115.110 1690.720 1115.430 1690.780 ;
        RECT 2900.830 1690.720 2901.150 1690.780 ;
        RECT 1115.110 1690.580 2901.150 1690.720 ;
        RECT 1115.110 1690.520 1115.430 1690.580 ;
        RECT 2900.830 1690.520 2901.150 1690.580 ;
      LAYER via ;
        RECT 1115.140 1690.520 1115.400 1690.780 ;
        RECT 2900.860 1690.520 2901.120 1690.780 ;
      LAYER met2 ;
        RECT 2900.850 1692.675 2901.130 1693.045 ;
        RECT 2900.920 1690.810 2901.060 1692.675 ;
        RECT 1115.140 1690.490 1115.400 1690.810 ;
        RECT 2900.860 1690.490 2901.120 1690.810 ;
        RECT 1115.200 509.845 1115.340 1690.490 ;
        RECT 1115.130 509.475 1115.410 509.845 ;
      LAYER via2 ;
        RECT 2900.850 1692.720 2901.130 1693.000 ;
        RECT 1115.130 509.520 1115.410 509.800 ;
      LAYER met3 ;
        RECT 2900.825 1693.010 2901.155 1693.025 ;
        RECT 2917.600 1693.010 2924.800 1693.460 ;
        RECT 2900.825 1692.710 2924.800 1693.010 ;
        RECT 2900.825 1692.695 2901.155 1692.710 ;
        RECT 2917.600 1692.260 2924.800 1692.710 ;
        RECT 1115.105 509.810 1115.435 509.825 ;
        RECT 1098.790 509.510 1115.435 509.810 ;
        RECT 1098.790 507.400 1099.090 509.510 ;
        RECT 1115.105 509.495 1115.435 509.510 ;
        RECT 1096.000 506.800 1100.000 507.400 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.250 400.180 1095.530 404.000 ;
        RECT 1095.250 400.000 1095.560 400.180 ;
        RECT 1095.420 394.245 1095.560 400.000 ;
        RECT 1095.350 393.875 1095.630 394.245 ;
      LAYER via2 ;
        RECT 1095.350 393.920 1095.630 394.200 ;
      LAYER met3 ;
        RECT -4.800 2704.170 2.400 2704.620 ;
        RECT 17.750 2704.170 18.130 2704.180 ;
        RECT -4.800 2703.870 18.130 2704.170 ;
        RECT -4.800 2703.420 2.400 2703.870 ;
        RECT 17.750 2703.860 18.130 2703.870 ;
        RECT 17.750 394.210 18.130 394.220 ;
        RECT 1095.325 394.210 1095.655 394.225 ;
        RECT 17.750 393.910 1095.655 394.210 ;
        RECT 17.750 393.900 18.130 393.910 ;
        RECT 1095.325 393.895 1095.655 393.910 ;
      LAYER via3 ;
        RECT 17.780 2703.860 18.100 2704.180 ;
        RECT 17.780 393.900 18.100 394.220 ;
      LAYER met4 ;
        RECT 17.775 2703.855 18.105 2704.185 ;
        RECT 17.790 394.225 18.090 2703.855 ;
        RECT 17.775 393.895 18.105 394.225 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2442.800 17.870 2442.860 ;
        RECT 1104.070 2442.800 1104.390 2442.860 ;
        RECT 17.550 2442.660 1104.390 2442.800 ;
        RECT 17.550 2442.600 17.870 2442.660 ;
        RECT 1104.070 2442.600 1104.390 2442.660 ;
      LAYER via ;
        RECT 17.580 2442.600 17.840 2442.860 ;
        RECT 1104.100 2442.600 1104.360 2442.860 ;
      LAYER met2 ;
        RECT 17.570 2443.395 17.850 2443.765 ;
        RECT 17.640 2442.890 17.780 2443.395 ;
        RECT 17.580 2442.570 17.840 2442.890 ;
        RECT 1104.100 2442.570 1104.360 2442.890 ;
        RECT 1104.160 895.405 1104.300 2442.570 ;
        RECT 1104.090 895.035 1104.370 895.405 ;
      LAYER via2 ;
        RECT 17.570 2443.440 17.850 2443.720 ;
        RECT 1104.090 895.080 1104.370 895.360 ;
      LAYER met3 ;
        RECT -4.800 2443.730 2.400 2444.180 ;
        RECT 17.545 2443.730 17.875 2443.745 ;
        RECT -4.800 2443.430 17.875 2443.730 ;
        RECT -4.800 2442.980 2.400 2443.430 ;
        RECT 17.545 2443.415 17.875 2443.430 ;
        RECT 1104.065 895.370 1104.395 895.385 ;
        RECT 1098.790 895.070 1104.395 895.370 ;
        RECT 1098.790 892.960 1099.090 895.070 ;
        RECT 1104.065 895.055 1104.395 895.070 ;
        RECT 1096.000 892.360 1100.000 892.960 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2180.660 17.870 2180.720 ;
        RECT 941.690 2180.660 942.010 2180.720 ;
        RECT 17.550 2180.520 942.010 2180.660 ;
        RECT 17.550 2180.460 17.870 2180.520 ;
        RECT 941.690 2180.460 942.010 2180.520 ;
        RECT 941.690 1011.740 942.010 1011.800 ;
        RECT 1094.870 1011.740 1095.190 1011.800 ;
        RECT 941.690 1011.600 1095.190 1011.740 ;
        RECT 941.690 1011.540 942.010 1011.600 ;
        RECT 1094.870 1011.540 1095.190 1011.600 ;
      LAYER via ;
        RECT 17.580 2180.460 17.840 2180.720 ;
        RECT 941.720 2180.460 941.980 2180.720 ;
        RECT 941.720 1011.540 941.980 1011.800 ;
        RECT 1094.900 1011.540 1095.160 1011.800 ;
      LAYER met2 ;
        RECT 17.570 2182.955 17.850 2183.325 ;
        RECT 17.640 2180.750 17.780 2182.955 ;
        RECT 17.580 2180.430 17.840 2180.750 ;
        RECT 941.720 2180.430 941.980 2180.750 ;
        RECT 941.780 1011.830 941.920 2180.430 ;
        RECT 941.720 1011.510 941.980 1011.830 ;
        RECT 1094.900 1011.510 1095.160 1011.830 ;
        RECT 1094.960 999.330 1095.100 1011.510 ;
        RECT 1096.170 999.330 1096.450 1000.000 ;
        RECT 1094.960 999.190 1096.450 999.330 ;
        RECT 1096.170 996.000 1096.450 999.190 ;
      LAYER via2 ;
        RECT 17.570 2183.000 17.850 2183.280 ;
      LAYER met3 ;
        RECT -4.800 2183.290 2.400 2183.740 ;
        RECT 17.545 2183.290 17.875 2183.305 ;
        RECT -4.800 2182.990 17.875 2183.290 ;
        RECT -4.800 2182.540 2.400 2182.990 ;
        RECT 17.545 2182.975 17.875 2182.990 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.790 1918.520 15.110 1918.580 ;
        RECT 1097.630 1918.520 1097.950 1918.580 ;
        RECT 14.790 1918.380 1097.950 1918.520 ;
        RECT 14.790 1918.320 15.110 1918.380 ;
        RECT 1097.630 1918.320 1097.950 1918.380 ;
      LAYER via ;
        RECT 14.820 1918.320 15.080 1918.580 ;
        RECT 1097.660 1918.320 1097.920 1918.580 ;
      LAYER met2 ;
        RECT 14.810 1921.835 15.090 1922.205 ;
        RECT 14.880 1918.610 15.020 1921.835 ;
        RECT 14.820 1918.290 15.080 1918.610 ;
        RECT 1097.660 1918.290 1097.920 1918.610 ;
        RECT 1097.720 938.245 1097.860 1918.290 ;
        RECT 1097.650 937.875 1097.930 938.245 ;
      LAYER via2 ;
        RECT 14.810 1921.880 15.090 1922.160 ;
        RECT 1097.650 937.920 1097.930 938.200 ;
      LAYER met3 ;
        RECT -4.800 1922.170 2.400 1922.620 ;
        RECT 14.785 1922.170 15.115 1922.185 ;
        RECT -4.800 1921.870 15.115 1922.170 ;
        RECT -4.800 1921.420 2.400 1921.870 ;
        RECT 14.785 1921.855 15.115 1921.870 ;
        RECT 1097.625 938.210 1097.955 938.225 ;
        RECT 1097.625 937.895 1098.170 938.210 ;
        RECT 1097.870 935.800 1098.170 937.895 ;
        RECT 1096.000 935.200 1100.000 935.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 890.020 15.570 890.080 ;
        RECT 18.010 890.020 18.330 890.080 ;
        RECT 15.250 889.880 18.330 890.020 ;
        RECT 15.250 889.820 15.570 889.880 ;
        RECT 18.010 889.820 18.330 889.880 ;
        RECT 15.250 876.080 15.570 876.140 ;
        RECT 190.050 876.080 190.370 876.140 ;
        RECT 15.250 875.940 190.370 876.080 ;
        RECT 15.250 875.880 15.570 875.940 ;
        RECT 190.050 875.880 190.370 875.940 ;
      LAYER via ;
        RECT 15.280 889.820 15.540 890.080 ;
        RECT 18.040 889.820 18.300 890.080 ;
        RECT 15.280 875.880 15.540 876.140 ;
        RECT 190.080 875.880 190.340 876.140 ;
      LAYER met2 ;
        RECT 18.030 1661.395 18.310 1661.765 ;
        RECT 18.100 890.110 18.240 1661.395 ;
        RECT 15.280 889.790 15.540 890.110 ;
        RECT 18.040 889.790 18.300 890.110 ;
        RECT 15.340 876.170 15.480 889.790 ;
        RECT 15.280 875.850 15.540 876.170 ;
        RECT 190.080 875.850 190.340 876.170 ;
        RECT 190.140 873.645 190.280 875.850 ;
        RECT 190.070 873.275 190.350 873.645 ;
      LAYER via2 ;
        RECT 18.030 1661.440 18.310 1661.720 ;
        RECT 190.070 873.320 190.350 873.600 ;
      LAYER met3 ;
        RECT -4.800 1661.730 2.400 1662.180 ;
        RECT 18.005 1661.730 18.335 1661.745 ;
        RECT -4.800 1661.430 18.335 1661.730 ;
        RECT -4.800 1660.980 2.400 1661.430 ;
        RECT 18.005 1661.415 18.335 1661.430 ;
        RECT 190.045 873.610 190.375 873.625 ;
        RECT 190.045 873.310 201.170 873.610 ;
        RECT 190.045 873.295 190.375 873.310 ;
        RECT 200.870 871.880 201.170 873.310 ;
        RECT 200.000 871.280 204.000 871.880 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1393.900 17.870 1393.960 ;
        RECT 1104.990 1393.900 1105.310 1393.960 ;
        RECT 17.550 1393.760 1105.310 1393.900 ;
        RECT 17.550 1393.700 17.870 1393.760 ;
        RECT 1104.990 1393.700 1105.310 1393.760 ;
      LAYER via ;
        RECT 17.580 1393.700 17.840 1393.960 ;
        RECT 1105.020 1393.700 1105.280 1393.960 ;
      LAYER met2 ;
        RECT 17.570 1400.275 17.850 1400.645 ;
        RECT 17.640 1393.990 17.780 1400.275 ;
        RECT 17.580 1393.670 17.840 1393.990 ;
        RECT 1105.020 1393.670 1105.280 1393.990 ;
        RECT 1105.080 979.725 1105.220 1393.670 ;
        RECT 1105.010 979.355 1105.290 979.725 ;
      LAYER via2 ;
        RECT 17.570 1400.320 17.850 1400.600 ;
        RECT 1105.010 979.400 1105.290 979.680 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.545 1400.610 17.875 1400.625 ;
        RECT -4.800 1400.310 17.875 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.545 1400.295 17.875 1400.310 ;
        RECT 1104.985 979.690 1105.315 979.705 ;
        RECT 1098.790 979.390 1105.315 979.690 ;
        RECT 1098.790 978.640 1099.090 979.390 ;
        RECT 1104.985 979.375 1105.315 979.390 ;
        RECT 1096.000 978.040 1100.000 978.640 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1138.900 17.870 1138.960 ;
        RECT 1098.090 1138.900 1098.410 1138.960 ;
        RECT 17.550 1138.760 1098.410 1138.900 ;
        RECT 17.550 1138.700 17.870 1138.760 ;
        RECT 1098.090 1138.700 1098.410 1138.760 ;
      LAYER via ;
        RECT 17.580 1138.700 17.840 1138.960 ;
        RECT 1098.120 1138.700 1098.380 1138.960 ;
      LAYER met2 ;
        RECT 17.570 1139.835 17.850 1140.205 ;
        RECT 17.640 1138.990 17.780 1139.835 ;
        RECT 17.580 1138.670 17.840 1138.990 ;
        RECT 1098.120 1138.670 1098.380 1138.990 ;
        RECT 1097.090 403.650 1097.370 404.000 ;
        RECT 1098.180 403.650 1098.320 1138.670 ;
        RECT 1097.090 403.510 1098.320 403.650 ;
        RECT 1097.090 400.000 1097.370 403.510 ;
      LAYER via2 ;
        RECT 17.570 1139.880 17.850 1140.160 ;
      LAYER met3 ;
        RECT -4.800 1140.170 2.400 1140.620 ;
        RECT 17.545 1140.170 17.875 1140.185 ;
        RECT -4.800 1139.870 17.875 1140.170 ;
        RECT -4.800 1139.420 2.400 1139.870 ;
        RECT 17.545 1139.855 17.875 1139.870 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.010 883.220 18.330 883.280 ;
        RECT 189.590 883.220 189.910 883.280 ;
        RECT 18.010 883.080 189.910 883.220 ;
        RECT 18.010 883.020 18.330 883.080 ;
        RECT 189.590 883.020 189.910 883.080 ;
      LAYER via ;
        RECT 18.040 883.020 18.300 883.280 ;
        RECT 189.620 883.020 189.880 883.280 ;
      LAYER met2 ;
        RECT 189.610 954.195 189.890 954.565 ;
        RECT 189.680 883.310 189.820 954.195 ;
        RECT 18.040 882.990 18.300 883.310 ;
        RECT 189.620 882.990 189.880 883.310 ;
        RECT 18.100 879.765 18.240 882.990 ;
        RECT 18.030 879.395 18.310 879.765 ;
      LAYER via2 ;
        RECT 189.610 954.240 189.890 954.520 ;
        RECT 18.030 879.440 18.310 879.720 ;
      LAYER met3 ;
        RECT 200.000 956.960 204.000 957.560 ;
        RECT 189.585 954.530 189.915 954.545 ;
        RECT 200.870 954.530 201.170 956.960 ;
        RECT 189.585 954.230 201.170 954.530 ;
        RECT 189.585 954.215 189.915 954.230 ;
        RECT -4.800 879.730 2.400 880.180 ;
        RECT 18.005 879.730 18.335 879.745 ;
        RECT -4.800 879.430 18.335 879.730 ;
        RECT -4.800 878.980 2.400 879.430 ;
        RECT 18.005 879.415 18.335 879.430 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1099.010 394.300 1099.330 394.360 ;
        RECT 1000.430 394.160 1099.330 394.300 ;
        RECT 17.090 393.620 17.410 393.680 ;
        RECT 1000.430 393.620 1000.570 394.160 ;
        RECT 1099.010 394.100 1099.330 394.160 ;
        RECT 17.090 393.480 1000.570 393.620 ;
        RECT 17.090 393.420 17.410 393.480 ;
      LAYER via ;
        RECT 17.120 393.420 17.380 393.680 ;
        RECT 1099.040 394.100 1099.300 394.360 ;
      LAYER met2 ;
        RECT 17.110 618.275 17.390 618.645 ;
        RECT 17.180 393.710 17.320 618.275 ;
        RECT 1098.930 400.180 1099.210 404.000 ;
        RECT 1098.930 400.000 1099.240 400.180 ;
        RECT 1099.100 394.390 1099.240 400.000 ;
        RECT 1099.040 394.070 1099.300 394.390 ;
        RECT 17.120 393.390 17.380 393.710 ;
      LAYER via2 ;
        RECT 17.110 618.320 17.390 618.600 ;
      LAYER met3 ;
        RECT -4.800 618.610 2.400 619.060 ;
        RECT 17.085 618.610 17.415 618.625 ;
        RECT -4.800 618.310 17.415 618.610 ;
        RECT -4.800 617.860 2.400 618.310 ;
        RECT 17.085 618.295 17.415 618.310 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.650 1952.860 1114.970 1952.920 ;
        RECT 2900.830 1952.860 2901.150 1952.920 ;
        RECT 1114.650 1952.720 2901.150 1952.860 ;
        RECT 1114.650 1952.660 1114.970 1952.720 ;
        RECT 2900.830 1952.660 2901.150 1952.720 ;
      LAYER via ;
        RECT 1114.680 1952.660 1114.940 1952.920 ;
        RECT 2900.860 1952.660 2901.120 1952.920 ;
      LAYER met2 ;
        RECT 2900.850 1958.555 2901.130 1958.925 ;
        RECT 2900.920 1952.950 2901.060 1958.555 ;
        RECT 1114.680 1952.630 1114.940 1952.950 ;
        RECT 2900.860 1952.630 2901.120 1952.950 ;
        RECT 1114.740 552.005 1114.880 1952.630 ;
        RECT 1114.670 551.635 1114.950 552.005 ;
      LAYER via2 ;
        RECT 2900.850 1958.600 2901.130 1958.880 ;
        RECT 1114.670 551.680 1114.950 551.960 ;
      LAYER met3 ;
        RECT 2900.825 1958.890 2901.155 1958.905 ;
        RECT 2917.600 1958.890 2924.800 1959.340 ;
        RECT 2900.825 1958.590 2924.800 1958.890 ;
        RECT 2900.825 1958.575 2901.155 1958.590 ;
        RECT 2917.600 1958.140 2924.800 1958.590 ;
        RECT 1114.645 551.970 1114.975 551.985 ;
        RECT 1098.790 551.670 1114.975 551.970 ;
        RECT 1098.790 550.240 1099.090 551.670 ;
        RECT 1114.645 551.655 1114.975 551.670 ;
        RECT 1096.000 549.640 1100.000 550.240 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1062.670 2222.140 1062.990 2222.200 ;
        RECT 2900.830 2222.140 2901.150 2222.200 ;
        RECT 1062.670 2222.000 2901.150 2222.140 ;
        RECT 1062.670 2221.940 1062.990 2222.000 ;
        RECT 2900.830 2221.940 2901.150 2222.000 ;
      LAYER via ;
        RECT 1062.700 2221.940 1062.960 2222.200 ;
        RECT 2900.860 2221.940 2901.120 2222.200 ;
      LAYER met2 ;
        RECT 2900.850 2223.755 2901.130 2224.125 ;
        RECT 2900.920 2222.230 2901.060 2223.755 ;
        RECT 1062.700 2221.910 1062.960 2222.230 ;
        RECT 2900.860 2221.910 2901.120 2222.230 ;
        RECT 1062.760 1048.870 1062.900 2221.910 ;
        RECT 1062.760 1048.730 1065.200 1048.870 ;
        RECT 1065.060 999.330 1065.200 1048.730 ;
        RECT 1066.730 999.330 1067.010 1000.000 ;
        RECT 1065.060 999.190 1067.010 999.330 ;
        RECT 1066.730 996.000 1067.010 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2223.800 2901.130 2224.080 ;
      LAYER met3 ;
        RECT 2900.825 2224.090 2901.155 2224.105 ;
        RECT 2917.600 2224.090 2924.800 2224.540 ;
        RECT 2900.825 2223.790 2924.800 2224.090 ;
        RECT 2900.825 2223.775 2901.155 2223.790 ;
        RECT 2917.600 2223.340 2924.800 2223.790 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.190 2484.280 1114.510 2484.340 ;
        RECT 2900.830 2484.280 2901.150 2484.340 ;
        RECT 1114.190 2484.140 2901.150 2484.280 ;
        RECT 1114.190 2484.080 1114.510 2484.140 ;
        RECT 2900.830 2484.080 2901.150 2484.140 ;
      LAYER via ;
        RECT 1114.220 2484.080 1114.480 2484.340 ;
        RECT 2900.860 2484.080 2901.120 2484.340 ;
      LAYER met2 ;
        RECT 2900.850 2489.635 2901.130 2490.005 ;
        RECT 2900.920 2484.370 2901.060 2489.635 ;
        RECT 1114.220 2484.050 1114.480 2484.370 ;
        RECT 2900.860 2484.050 2901.120 2484.370 ;
        RECT 1114.280 592.125 1114.420 2484.050 ;
        RECT 1114.210 591.755 1114.490 592.125 ;
      LAYER via2 ;
        RECT 2900.850 2489.680 2901.130 2489.960 ;
        RECT 1114.210 591.800 1114.490 592.080 ;
      LAYER met3 ;
        RECT 2900.825 2489.970 2901.155 2489.985 ;
        RECT 2917.600 2489.970 2924.800 2490.420 ;
        RECT 2900.825 2489.670 2924.800 2489.970 ;
        RECT 2900.825 2489.655 2901.155 2489.670 ;
        RECT 2917.600 2489.220 2924.800 2489.670 ;
        RECT 1096.000 592.480 1100.000 593.080 ;
        RECT 1098.790 592.090 1099.090 592.480 ;
        RECT 1114.185 592.090 1114.515 592.105 ;
        RECT 1098.790 591.790 1114.515 592.090 ;
        RECT 1114.185 591.775 1114.515 591.790 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.350 2753.220 192.670 2753.280 ;
        RECT 2900.830 2753.220 2901.150 2753.280 ;
        RECT 192.350 2753.080 2901.150 2753.220 ;
        RECT 192.350 2753.020 192.670 2753.080 ;
        RECT 2900.830 2753.020 2901.150 2753.080 ;
      LAYER via ;
        RECT 192.380 2753.020 192.640 2753.280 ;
        RECT 2900.860 2753.020 2901.120 2753.280 ;
      LAYER met2 ;
        RECT 2900.850 2755.515 2901.130 2755.885 ;
        RECT 2900.920 2753.310 2901.060 2755.515 ;
        RECT 192.380 2752.990 192.640 2753.310 ;
        RECT 2900.860 2752.990 2901.120 2753.310 ;
        RECT 192.440 445.925 192.580 2752.990 ;
        RECT 192.370 445.555 192.650 445.925 ;
      LAYER via2 ;
        RECT 2900.850 2755.560 2901.130 2755.840 ;
        RECT 192.370 445.600 192.650 445.880 ;
      LAYER met3 ;
        RECT 2900.825 2755.850 2901.155 2755.865 ;
        RECT 2917.600 2755.850 2924.800 2756.300 ;
        RECT 2900.825 2755.550 2924.800 2755.850 ;
        RECT 2900.825 2755.535 2901.155 2755.550 ;
        RECT 2917.600 2755.100 2924.800 2755.550 ;
        RECT 192.345 445.890 192.675 445.905 ;
        RECT 192.345 445.590 201.170 445.890 ;
        RECT 192.345 445.575 192.675 445.590 ;
        RECT 200.870 443.480 201.170 445.590 ;
        RECT 200.000 442.880 204.000 443.480 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.570 3015.700 1069.890 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1069.570 3015.560 2901.150 3015.700 ;
        RECT 1069.570 3015.500 1069.890 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1069.600 3015.500 1069.860 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1069.600 3015.470 1069.860 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1069.660 1048.870 1069.800 3015.470 ;
        RECT 1069.660 1048.730 1072.560 1048.870 ;
        RECT 1072.420 999.330 1072.560 1048.730 ;
        RECT 1074.090 999.330 1074.370 1000.000 ;
        RECT 1072.420 999.190 1074.370 999.330 ;
        RECT 1074.090 996.000 1074.370 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 192.810 3284.640 193.130 3284.700 ;
        RECT 2900.830 3284.640 2901.150 3284.700 ;
        RECT 192.810 3284.500 2901.150 3284.640 ;
        RECT 192.810 3284.440 193.130 3284.500 ;
        RECT 2900.830 3284.440 2901.150 3284.500 ;
      LAYER via ;
        RECT 192.840 3284.440 193.100 3284.700 ;
        RECT 2900.860 3284.440 2901.120 3284.700 ;
      LAYER met2 ;
        RECT 2900.850 3286.595 2901.130 3286.965 ;
        RECT 2900.920 3284.730 2901.060 3286.595 ;
        RECT 192.840 3284.410 193.100 3284.730 ;
        RECT 2900.860 3284.410 2901.120 3284.730 ;
        RECT 192.900 530.925 193.040 3284.410 ;
        RECT 192.830 530.555 193.110 530.925 ;
      LAYER via2 ;
        RECT 2900.850 3286.640 2901.130 3286.920 ;
        RECT 192.830 530.600 193.110 530.880 ;
      LAYER met3 ;
        RECT 2900.825 3286.930 2901.155 3286.945 ;
        RECT 2917.600 3286.930 2924.800 3287.380 ;
        RECT 2900.825 3286.630 2924.800 3286.930 ;
        RECT 2900.825 3286.615 2901.155 3286.630 ;
        RECT 2917.600 3286.180 2924.800 3286.630 ;
        RECT 192.805 530.890 193.135 530.905 ;
        RECT 192.805 530.590 201.170 530.890 ;
        RECT 192.805 530.575 193.135 530.590 ;
        RECT 200.870 529.160 201.170 530.590 ;
        RECT 200.000 528.560 204.000 529.160 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 191.890 1003.920 192.210 1003.980 ;
        RECT 2877.370 1003.920 2877.690 1003.980 ;
        RECT 191.890 1003.780 2877.690 1003.920 ;
        RECT 191.890 1003.720 192.210 1003.780 ;
        RECT 2877.370 1003.720 2877.690 1003.780 ;
      LAYER via ;
        RECT 191.920 1003.720 192.180 1003.980 ;
        RECT 2877.400 1003.720 2877.660 1003.980 ;
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
        RECT 2879.300 3512.170 2879.440 3517.600 ;
        RECT 2877.460 3512.030 2879.440 3512.170 ;
        RECT 2877.460 1004.010 2877.600 3512.030 ;
        RECT 191.920 1003.690 192.180 1004.010 ;
        RECT 2877.400 1003.690 2877.660 1004.010 ;
        RECT 191.980 617.285 192.120 1003.690 ;
        RECT 191.910 616.915 192.190 617.285 ;
      LAYER via2 ;
        RECT 191.910 616.960 192.190 617.240 ;
      LAYER met3 ;
        RECT 191.885 617.250 192.215 617.265 ;
        RECT 191.885 616.950 201.170 617.250 ;
        RECT 191.885 616.935 192.215 616.950 ;
        RECT 200.870 614.840 201.170 616.950 ;
        RECT 200.000 614.240 204.000 614.840 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.410 641.480 1117.730 641.540 ;
        RECT 2553.070 641.480 2553.390 641.540 ;
        RECT 1117.410 641.340 2553.390 641.480 ;
        RECT 1117.410 641.280 1117.730 641.340 ;
        RECT 2553.070 641.280 2553.390 641.340 ;
      LAYER via ;
        RECT 1117.440 641.280 1117.700 641.540 ;
        RECT 2553.100 641.280 2553.360 641.540 ;
      LAYER met2 ;
        RECT 2553.160 3517.910 2554.220 3518.050 ;
        RECT 2553.160 641.570 2553.300 3517.910 ;
        RECT 2554.080 3517.370 2554.220 3517.910 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
        RECT 2555.000 3517.370 2555.140 3517.600 ;
        RECT 2554.080 3517.230 2555.140 3517.370 ;
        RECT 1117.440 641.250 1117.700 641.570 ;
        RECT 2553.100 641.250 2553.360 641.570 ;
        RECT 1117.500 638.365 1117.640 641.250 ;
        RECT 1117.430 637.995 1117.710 638.365 ;
      LAYER via2 ;
        RECT 1117.430 638.040 1117.710 638.320 ;
      LAYER met3 ;
        RECT 1117.405 638.330 1117.735 638.345 ;
        RECT 1098.790 638.030 1117.735 638.330 ;
        RECT 1098.790 635.920 1099.090 638.030 ;
        RECT 1117.405 638.015 1117.735 638.030 ;
        RECT 1096.000 635.320 1100.000 635.920 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 201.550 327.800 201.870 328.060 ;
        RECT 201.640 327.040 201.780 327.800 ;
        RECT 201.550 326.780 201.870 327.040 ;
      LAYER via ;
        RECT 201.580 327.800 201.840 328.060 ;
        RECT 201.580 326.780 201.840 327.040 ;
      LAYER met2 ;
        RECT 203.770 996.610 204.050 1000.000 ;
        RECT 201.640 996.470 204.050 996.610 ;
        RECT 201.640 420.970 201.780 996.470 ;
        RECT 203.770 996.000 204.050 996.470 ;
        RECT 200.260 420.830 201.780 420.970 ;
        RECT 200.260 396.850 200.400 420.830 ;
        RECT 200.260 396.710 201.780 396.850 ;
        RECT 201.640 328.090 201.780 396.710 ;
        RECT 201.580 327.770 201.840 328.090 ;
        RECT 201.580 326.750 201.840 327.070 ;
        RECT 201.640 107.285 201.780 326.750 ;
        RECT 201.570 106.915 201.850 107.285 ;
        RECT 2901.770 106.915 2902.050 107.285 ;
        RECT 2901.840 33.165 2901.980 106.915 ;
        RECT 2901.770 32.795 2902.050 33.165 ;
      LAYER via2 ;
        RECT 201.570 106.960 201.850 107.240 ;
        RECT 2901.770 106.960 2902.050 107.240 ;
        RECT 2901.770 32.840 2902.050 33.120 ;
      LAYER met3 ;
        RECT 201.545 107.250 201.875 107.265 ;
        RECT 2901.745 107.250 2902.075 107.265 ;
        RECT 201.545 106.950 2902.075 107.250 ;
        RECT 201.545 106.935 201.875 106.950 ;
        RECT 2901.745 106.935 2902.075 106.950 ;
        RECT 2901.745 33.130 2902.075 33.145 ;
        RECT 2917.600 33.130 2924.800 33.580 ;
        RECT 2901.745 32.830 2924.800 33.130 ;
        RECT 2901.745 32.815 2902.075 32.830 ;
        RECT 2917.600 32.380 2924.800 32.830 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 2284.020 421.290 2284.080 ;
        RECT 2900.830 2284.020 2901.150 2284.080 ;
        RECT 420.970 2283.880 2901.150 2284.020 ;
        RECT 420.970 2283.820 421.290 2283.880 ;
        RECT 2900.830 2283.820 2901.150 2283.880 ;
      LAYER via ;
        RECT 421.000 2283.820 421.260 2284.080 ;
        RECT 2900.860 2283.820 2901.120 2284.080 ;
      LAYER met2 ;
        RECT 2900.850 2290.395 2901.130 2290.765 ;
        RECT 2900.920 2284.110 2901.060 2290.395 ;
        RECT 421.000 2283.790 421.260 2284.110 ;
        RECT 2900.860 2283.790 2901.120 2284.110 ;
        RECT 421.060 1048.870 421.200 2283.790 ;
        RECT 421.060 1048.730 424.880 1048.870 ;
        RECT 424.740 999.330 424.880 1048.730 ;
        RECT 426.870 999.330 427.150 1000.000 ;
        RECT 424.740 999.190 427.150 999.330 ;
        RECT 426.870 996.000 427.150 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2290.440 2901.130 2290.720 ;
      LAYER met3 ;
        RECT 2900.825 2290.730 2901.155 2290.745 ;
        RECT 2917.600 2290.730 2924.800 2291.180 ;
        RECT 2900.825 2290.430 2924.800 2290.730 ;
        RECT 2900.825 2290.415 2901.155 2290.430 ;
        RECT 2917.600 2289.980 2924.800 2290.430 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 2553.300 448.890 2553.360 ;
        RECT 2900.830 2553.300 2901.150 2553.360 ;
        RECT 448.570 2553.160 2901.150 2553.300 ;
        RECT 448.570 2553.100 448.890 2553.160 ;
        RECT 2900.830 2553.100 2901.150 2553.160 ;
      LAYER via ;
        RECT 448.600 2553.100 448.860 2553.360 ;
        RECT 2900.860 2553.100 2901.120 2553.360 ;
      LAYER met2 ;
        RECT 2900.850 2556.275 2901.130 2556.645 ;
        RECT 2900.920 2553.390 2901.060 2556.275 ;
        RECT 448.600 2553.070 448.860 2553.390 ;
        RECT 2900.860 2553.070 2901.120 2553.390 ;
        RECT 448.660 999.330 448.800 2553.070 ;
        RECT 448.950 999.330 449.230 1000.000 ;
        RECT 448.660 999.190 449.230 999.330 ;
        RECT 448.950 996.000 449.230 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2556.320 2901.130 2556.600 ;
      LAYER met3 ;
        RECT 2900.825 2556.610 2901.155 2556.625 ;
        RECT 2917.600 2556.610 2924.800 2557.060 ;
        RECT 2900.825 2556.310 2924.800 2556.610 ;
        RECT 2900.825 2556.295 2901.155 2556.310 ;
        RECT 2917.600 2555.860 2924.800 2556.310 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 2815.440 469.590 2815.500 ;
        RECT 2898.990 2815.440 2899.310 2815.500 ;
        RECT 469.270 2815.300 2899.310 2815.440 ;
        RECT 469.270 2815.240 469.590 2815.300 ;
        RECT 2898.990 2815.240 2899.310 2815.300 ;
      LAYER via ;
        RECT 469.300 2815.240 469.560 2815.500 ;
        RECT 2899.020 2815.240 2899.280 2815.500 ;
      LAYER met2 ;
        RECT 2899.010 2821.475 2899.290 2821.845 ;
        RECT 2899.080 2815.530 2899.220 2821.475 ;
        RECT 469.300 2815.210 469.560 2815.530 ;
        RECT 2899.020 2815.210 2899.280 2815.530 ;
        RECT 469.360 1048.870 469.500 2815.210 ;
        RECT 469.360 1048.730 469.960 1048.870 ;
        RECT 469.820 999.330 469.960 1048.730 ;
        RECT 471.490 999.330 471.770 1000.000 ;
        RECT 469.820 999.190 471.770 999.330 ;
        RECT 471.490 996.000 471.770 999.190 ;
      LAYER via2 ;
        RECT 2899.010 2821.520 2899.290 2821.800 ;
      LAYER met3 ;
        RECT 2898.985 2821.810 2899.315 2821.825 ;
        RECT 2917.600 2821.810 2924.800 2822.260 ;
        RECT 2898.985 2821.510 2924.800 2821.810 ;
        RECT 2898.985 2821.495 2899.315 2821.510 ;
        RECT 2917.600 2821.060 2924.800 2821.510 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 3084.380 490.290 3084.440 ;
        RECT 2900.830 3084.380 2901.150 3084.440 ;
        RECT 489.970 3084.240 2901.150 3084.380 ;
        RECT 489.970 3084.180 490.290 3084.240 ;
        RECT 2900.830 3084.180 2901.150 3084.240 ;
      LAYER via ;
        RECT 490.000 3084.180 490.260 3084.440 ;
        RECT 2900.860 3084.180 2901.120 3084.440 ;
      LAYER met2 ;
        RECT 2900.850 3087.355 2901.130 3087.725 ;
        RECT 2900.920 3084.470 2901.060 3087.355 ;
        RECT 490.000 3084.150 490.260 3084.470 ;
        RECT 2900.860 3084.150 2901.120 3084.470 ;
        RECT 490.060 1048.870 490.200 3084.150 ;
        RECT 490.060 1048.730 492.040 1048.870 ;
        RECT 491.900 999.330 492.040 1048.730 ;
        RECT 493.570 999.330 493.850 1000.000 ;
        RECT 491.900 999.190 493.850 999.330 ;
        RECT 493.570 996.000 493.850 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3087.400 2901.130 3087.680 ;
      LAYER met3 ;
        RECT 2900.825 3087.690 2901.155 3087.705 ;
        RECT 2917.600 3087.690 2924.800 3088.140 ;
        RECT 2900.825 3087.390 2924.800 3087.690 ;
        RECT 2900.825 3087.375 2901.155 3087.390 ;
        RECT 2917.600 3086.940 2924.800 3087.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 3353.660 510.990 3353.720 ;
        RECT 2900.830 3353.660 2901.150 3353.720 ;
        RECT 510.670 3353.520 2901.150 3353.660 ;
        RECT 510.670 3353.460 510.990 3353.520 ;
        RECT 2900.830 3353.460 2901.150 3353.520 ;
      LAYER via ;
        RECT 510.700 3353.460 510.960 3353.720 ;
        RECT 2900.860 3353.460 2901.120 3353.720 ;
      LAYER met2 ;
        RECT 510.700 3353.430 510.960 3353.750 ;
        RECT 2900.860 3353.605 2901.120 3353.750 ;
        RECT 510.760 1048.870 510.900 3353.430 ;
        RECT 2900.850 3353.235 2901.130 3353.605 ;
        RECT 510.760 1048.730 514.120 1048.870 ;
        RECT 513.980 999.330 514.120 1048.730 ;
        RECT 516.110 999.330 516.390 1000.000 ;
        RECT 513.980 999.190 516.390 999.330 ;
        RECT 516.110 996.000 516.390 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3353.280 2901.130 3353.560 ;
      LAYER met3 ;
        RECT 2900.825 3353.570 2901.155 3353.585 ;
        RECT 2917.600 3353.570 2924.800 3354.020 ;
        RECT 2900.825 3353.270 2924.800 3353.570 ;
        RECT 2900.825 3353.255 2901.155 3353.270 ;
        RECT 2917.600 3352.820 2924.800 3353.270 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 1017.860 539.050 1017.920 ;
        RECT 2794.570 1017.860 2794.890 1017.920 ;
        RECT 538.730 1017.720 2794.890 1017.860 ;
        RECT 538.730 1017.660 539.050 1017.720 ;
        RECT 2794.570 1017.660 2794.890 1017.720 ;
      LAYER via ;
        RECT 538.760 1017.660 539.020 1017.920 ;
        RECT 2794.600 1017.660 2794.860 1017.920 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3512.170 2798.480 3517.600 ;
        RECT 2794.660 3512.030 2798.480 3512.170 ;
        RECT 2794.660 1017.950 2794.800 3512.030 ;
        RECT 538.760 1017.630 539.020 1017.950 ;
        RECT 2794.600 1017.630 2794.860 1017.950 ;
        RECT 538.190 999.330 538.470 1000.000 ;
        RECT 538.820 999.330 538.960 1017.630 ;
        RECT 538.190 999.190 538.960 999.330 ;
        RECT 538.190 996.000 538.470 999.190 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 1018.200 559.290 1018.260 ;
        RECT 2470.270 1018.200 2470.590 1018.260 ;
        RECT 558.970 1018.060 2470.590 1018.200 ;
        RECT 558.970 1018.000 559.290 1018.060 ;
        RECT 2470.270 1018.000 2470.590 1018.060 ;
      LAYER via ;
        RECT 559.000 1018.000 559.260 1018.260 ;
        RECT 2470.300 1018.000 2470.560 1018.260 ;
      LAYER met2 ;
        RECT 2470.360 3517.910 2473.260 3518.050 ;
        RECT 2470.360 1018.290 2470.500 3517.910 ;
        RECT 2473.120 3517.370 2473.260 3517.910 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2473.120 3517.230 2474.180 3517.370 ;
        RECT 559.000 1017.970 559.260 1018.290 ;
        RECT 2470.300 1017.970 2470.560 1018.290 ;
        RECT 559.060 999.330 559.200 1017.970 ;
        RECT 560.730 999.330 561.010 1000.000 ;
        RECT 559.060 999.190 561.010 999.330 ;
        RECT 560.730 996.000 561.010 999.190 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.050 1018.540 581.370 1018.600 ;
        RECT 2145.970 1018.540 2146.290 1018.600 ;
        RECT 581.050 1018.400 2146.290 1018.540 ;
        RECT 581.050 1018.340 581.370 1018.400 ;
        RECT 2145.970 1018.340 2146.290 1018.400 ;
      LAYER via ;
        RECT 581.080 1018.340 581.340 1018.600 ;
        RECT 2146.000 1018.340 2146.260 1018.600 ;
      LAYER met2 ;
        RECT 2146.060 3517.910 2148.500 3518.050 ;
        RECT 2146.060 1018.630 2146.200 3517.910 ;
        RECT 2148.360 3517.370 2148.500 3517.910 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2148.360 3517.230 2149.420 3517.370 ;
        RECT 581.080 1018.310 581.340 1018.630 ;
        RECT 2146.000 1018.310 2146.260 1018.630 ;
        RECT 581.140 999.330 581.280 1018.310 ;
        RECT 582.810 999.330 583.090 1000.000 ;
        RECT 581.140 999.190 583.090 999.330 ;
        RECT 582.810 996.000 583.090 999.190 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 603.130 1018.880 603.450 1018.940 ;
        RECT 1821.670 1018.880 1821.990 1018.940 ;
        RECT 603.130 1018.740 1821.990 1018.880 ;
        RECT 603.130 1018.680 603.450 1018.740 ;
        RECT 1821.670 1018.680 1821.990 1018.740 ;
      LAYER via ;
        RECT 603.160 1018.680 603.420 1018.940 ;
        RECT 1821.700 1018.680 1821.960 1018.940 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3512.170 1825.120 3517.600 ;
        RECT 1821.760 3512.030 1825.120 3512.170 ;
        RECT 1821.760 1018.970 1821.900 3512.030 ;
        RECT 603.160 1018.650 603.420 1018.970 ;
        RECT 1821.700 1018.650 1821.960 1018.970 ;
        RECT 603.220 999.330 603.360 1018.650 ;
        RECT 605.350 999.330 605.630 1000.000 ;
        RECT 603.220 999.190 605.630 999.330 ;
        RECT 605.350 996.000 605.630 999.190 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1052.090 3504.620 1052.410 3504.680 ;
        RECT 1500.590 3504.620 1500.910 3504.680 ;
        RECT 1052.090 3504.480 1500.910 3504.620 ;
        RECT 1052.090 3504.420 1052.410 3504.480 ;
        RECT 1500.590 3504.420 1500.910 3504.480 ;
        RECT 625.210 1021.260 625.530 1021.320 ;
        RECT 1052.090 1021.260 1052.410 1021.320 ;
        RECT 625.210 1021.120 1052.410 1021.260 ;
        RECT 625.210 1021.060 625.530 1021.120 ;
        RECT 1052.090 1021.060 1052.410 1021.120 ;
      LAYER via ;
        RECT 1052.120 3504.420 1052.380 3504.680 ;
        RECT 1500.620 3504.420 1500.880 3504.680 ;
        RECT 625.240 1021.060 625.500 1021.320 ;
        RECT 1052.120 1021.060 1052.380 1021.320 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3504.710 1500.820 3517.600 ;
        RECT 1052.120 3504.390 1052.380 3504.710 ;
        RECT 1500.620 3504.390 1500.880 3504.710 ;
        RECT 1052.180 1021.350 1052.320 3504.390 ;
        RECT 625.240 1021.030 625.500 1021.350 ;
        RECT 1052.120 1021.030 1052.380 1021.350 ;
        RECT 625.300 999.330 625.440 1021.030 ;
        RECT 627.430 999.330 627.710 1000.000 ;
        RECT 625.300 999.190 627.710 999.330 ;
        RECT 627.430 996.000 627.710 999.190 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 227.770 997.260 228.090 997.520 ;
        RECT 227.860 995.420 228.000 997.260 ;
        RECT 227.860 995.280 276.070 995.420 ;
        RECT 275.930 994.060 276.070 995.280 ;
        RECT 2902.210 994.060 2902.530 994.120 ;
        RECT 275.930 993.920 2902.530 994.060 ;
        RECT 2902.210 993.860 2902.530 993.920 ;
      LAYER via ;
        RECT 227.800 997.260 228.060 997.520 ;
        RECT 2902.240 993.860 2902.500 994.120 ;
      LAYER met2 ;
        RECT 225.850 997.290 226.130 1000.000 ;
        RECT 227.800 997.290 228.060 997.550 ;
        RECT 225.850 997.230 228.060 997.290 ;
        RECT 225.850 997.150 228.000 997.230 ;
        RECT 225.850 996.000 226.130 997.150 ;
        RECT 2902.240 993.830 2902.500 994.150 ;
        RECT 2902.300 231.725 2902.440 993.830 ;
        RECT 2902.230 231.355 2902.510 231.725 ;
      LAYER via2 ;
        RECT 2902.230 231.400 2902.510 231.680 ;
      LAYER met3 ;
        RECT 2902.205 231.690 2902.535 231.705 ;
        RECT 2917.600 231.690 2924.800 232.140 ;
        RECT 2902.205 231.390 2924.800 231.690 ;
        RECT 2902.205 231.375 2902.535 231.390 ;
        RECT 2917.600 230.940 2924.800 231.390 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1052.550 3500.880 1052.870 3500.940 ;
        RECT 1175.830 3500.880 1176.150 3500.940 ;
        RECT 1052.550 3500.740 1176.150 3500.880 ;
        RECT 1052.550 3500.680 1052.870 3500.740 ;
        RECT 1175.830 3500.680 1176.150 3500.740 ;
        RECT 648.670 1017.520 648.990 1017.580 ;
        RECT 1052.550 1017.520 1052.870 1017.580 ;
        RECT 648.670 1017.380 1052.870 1017.520 ;
        RECT 648.670 1017.320 648.990 1017.380 ;
        RECT 1052.550 1017.320 1052.870 1017.380 ;
      LAYER via ;
        RECT 1052.580 3500.680 1052.840 3500.940 ;
        RECT 1175.860 3500.680 1176.120 3500.940 ;
        RECT 648.700 1017.320 648.960 1017.580 ;
        RECT 1052.580 1017.320 1052.840 1017.580 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3500.970 1176.060 3517.600 ;
        RECT 1052.580 3500.650 1052.840 3500.970 ;
        RECT 1175.860 3500.650 1176.120 3500.970 ;
        RECT 1052.640 1017.610 1052.780 3500.650 ;
        RECT 648.700 1017.290 648.960 1017.610 ;
        RECT 1052.580 1017.290 1052.840 1017.610 ;
        RECT 648.760 999.330 648.900 1017.290 ;
        RECT 649.970 999.330 650.250 1000.000 ;
        RECT 648.760 999.190 650.250 999.330 ;
        RECT 649.970 996.000 650.250 999.190 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.370 3501.220 669.690 3501.280 ;
        RECT 851.530 3501.220 851.850 3501.280 ;
        RECT 669.370 3501.080 851.850 3501.220 ;
        RECT 669.370 3501.020 669.690 3501.080 ;
        RECT 851.530 3501.020 851.850 3501.080 ;
      LAYER via ;
        RECT 669.400 3501.020 669.660 3501.280 ;
        RECT 851.560 3501.020 851.820 3501.280 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.310 851.760 3517.600 ;
        RECT 669.400 3500.990 669.660 3501.310 ;
        RECT 851.560 3500.990 851.820 3501.310 ;
        RECT 669.460 1048.870 669.600 3500.990 ;
        RECT 669.460 1048.730 670.520 1048.870 ;
        RECT 670.380 999.330 670.520 1048.730 ;
        RECT 672.050 999.330 672.330 1000.000 ;
        RECT 670.380 999.190 672.330 999.330 ;
        RECT 672.050 996.000 672.330 999.190 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.230 3500.880 527.550 3500.940 ;
        RECT 690.070 3500.880 690.390 3500.940 ;
        RECT 527.230 3500.740 690.390 3500.880 ;
        RECT 527.230 3500.680 527.550 3500.740 ;
        RECT 690.070 3500.680 690.390 3500.740 ;
      LAYER via ;
        RECT 527.260 3500.680 527.520 3500.940 ;
        RECT 690.100 3500.680 690.360 3500.940 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3500.970 527.460 3517.600 ;
        RECT 527.260 3500.650 527.520 3500.970 ;
        RECT 690.100 3500.650 690.360 3500.970 ;
        RECT 690.160 1048.870 690.300 3500.650 ;
        RECT 690.160 1048.730 692.600 1048.870 ;
        RECT 692.460 999.330 692.600 1048.730 ;
        RECT 694.590 999.330 694.870 1000.000 ;
        RECT 692.460 999.190 694.870 999.330 ;
        RECT 694.590 996.000 694.870 999.190 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 202.470 3503.260 202.790 3503.320 ;
        RECT 224.090 3503.260 224.410 3503.320 ;
        RECT 202.470 3503.120 224.410 3503.260 ;
        RECT 202.470 3503.060 202.790 3503.120 ;
        RECT 224.090 3503.060 224.410 3503.120 ;
        RECT 224.090 1020.580 224.410 1020.640 ;
        RECT 714.450 1020.580 714.770 1020.640 ;
        RECT 224.090 1020.440 714.770 1020.580 ;
        RECT 224.090 1020.380 224.410 1020.440 ;
        RECT 714.450 1020.380 714.770 1020.440 ;
      LAYER via ;
        RECT 202.500 3503.060 202.760 3503.320 ;
        RECT 224.120 3503.060 224.380 3503.320 ;
        RECT 224.120 1020.380 224.380 1020.640 ;
        RECT 714.480 1020.380 714.740 1020.640 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3503.350 202.700 3517.600 ;
        RECT 202.500 3503.030 202.760 3503.350 ;
        RECT 224.120 3503.030 224.380 3503.350 ;
        RECT 224.180 1020.670 224.320 3503.030 ;
        RECT 224.120 1020.350 224.380 1020.670 ;
        RECT 714.480 1020.350 714.740 1020.670 ;
        RECT 714.540 999.330 714.680 1020.350 ;
        RECT 716.670 999.330 716.950 1000.000 ;
        RECT 714.540 999.190 716.950 999.330 ;
        RECT 716.670 996.000 716.950 999.190 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 3415.880 16.030 3415.940 ;
        RECT 224.550 3415.880 224.870 3415.940 ;
        RECT 15.710 3415.740 224.870 3415.880 ;
        RECT 15.710 3415.680 16.030 3415.740 ;
        RECT 224.550 3415.680 224.870 3415.740 ;
        RECT 224.550 1020.240 224.870 1020.300 ;
        RECT 738.370 1020.240 738.690 1020.300 ;
        RECT 224.550 1020.100 738.690 1020.240 ;
        RECT 224.550 1020.040 224.870 1020.100 ;
        RECT 738.370 1020.040 738.690 1020.100 ;
      LAYER via ;
        RECT 15.740 3415.680 16.000 3415.940 ;
        RECT 224.580 3415.680 224.840 3415.940 ;
        RECT 224.580 1020.040 224.840 1020.300 ;
        RECT 738.400 1020.040 738.660 1020.300 ;
      LAYER met2 ;
        RECT 15.730 3421.235 16.010 3421.605 ;
        RECT 15.800 3415.970 15.940 3421.235 ;
        RECT 15.740 3415.650 16.000 3415.970 ;
        RECT 224.580 3415.650 224.840 3415.970 ;
        RECT 224.640 1020.330 224.780 3415.650 ;
        RECT 224.580 1020.010 224.840 1020.330 ;
        RECT 738.400 1020.010 738.660 1020.330 ;
        RECT 738.460 999.330 738.600 1020.010 ;
        RECT 739.210 999.330 739.490 1000.000 ;
        RECT 738.460 999.190 739.490 999.330 ;
        RECT 739.210 996.000 739.490 999.190 ;
      LAYER via2 ;
        RECT 15.730 3421.280 16.010 3421.560 ;
      LAYER met3 ;
        RECT -4.800 3421.570 2.400 3422.020 ;
        RECT 15.705 3421.570 16.035 3421.585 ;
        RECT -4.800 3421.270 16.035 3421.570 ;
        RECT -4.800 3420.820 2.400 3421.270 ;
        RECT 15.705 3421.255 16.035 3421.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3160.540 17.870 3160.600 ;
        RECT 225.010 3160.540 225.330 3160.600 ;
        RECT 17.550 3160.400 225.330 3160.540 ;
        RECT 17.550 3160.340 17.870 3160.400 ;
        RECT 225.010 3160.340 225.330 3160.400 ;
        RECT 225.010 1019.560 225.330 1019.620 ;
        RECT 759.530 1019.560 759.850 1019.620 ;
        RECT 225.010 1019.420 759.850 1019.560 ;
        RECT 225.010 1019.360 225.330 1019.420 ;
        RECT 759.530 1019.360 759.850 1019.420 ;
      LAYER via ;
        RECT 17.580 3160.340 17.840 3160.600 ;
        RECT 225.040 3160.340 225.300 3160.600 ;
        RECT 225.040 1019.360 225.300 1019.620 ;
        RECT 759.560 1019.360 759.820 1019.620 ;
      LAYER met2 ;
        RECT 17.580 3160.485 17.840 3160.630 ;
        RECT 17.570 3160.115 17.850 3160.485 ;
        RECT 225.040 3160.310 225.300 3160.630 ;
        RECT 225.100 1019.650 225.240 3160.310 ;
        RECT 225.040 1019.330 225.300 1019.650 ;
        RECT 759.560 1019.330 759.820 1019.650 ;
        RECT 759.620 999.330 759.760 1019.330 ;
        RECT 761.750 999.330 762.030 1000.000 ;
        RECT 759.620 999.190 762.030 999.330 ;
        RECT 761.750 996.000 762.030 999.190 ;
      LAYER via2 ;
        RECT 17.570 3160.160 17.850 3160.440 ;
      LAYER met3 ;
        RECT -4.800 3160.450 2.400 3160.900 ;
        RECT 17.545 3160.450 17.875 3160.465 ;
        RECT -4.800 3160.150 17.875 3160.450 ;
        RECT -4.800 3159.700 2.400 3160.150 ;
        RECT 17.545 3160.135 17.875 3160.150 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2898.400 16.950 2898.460 ;
        RECT 225.470 2898.400 225.790 2898.460 ;
        RECT 16.630 2898.260 225.790 2898.400 ;
        RECT 16.630 2898.200 16.950 2898.260 ;
        RECT 225.470 2898.200 225.790 2898.260 ;
        RECT 225.470 1019.220 225.790 1019.280 ;
        RECT 781.610 1019.220 781.930 1019.280 ;
        RECT 225.470 1019.080 781.930 1019.220 ;
        RECT 225.470 1019.020 225.790 1019.080 ;
        RECT 781.610 1019.020 781.930 1019.080 ;
      LAYER via ;
        RECT 16.660 2898.200 16.920 2898.460 ;
        RECT 225.500 2898.200 225.760 2898.460 ;
        RECT 225.500 1019.020 225.760 1019.280 ;
        RECT 781.640 1019.020 781.900 1019.280 ;
      LAYER met2 ;
        RECT 16.650 2899.675 16.930 2900.045 ;
        RECT 16.720 2898.490 16.860 2899.675 ;
        RECT 16.660 2898.170 16.920 2898.490 ;
        RECT 225.500 2898.170 225.760 2898.490 ;
        RECT 225.560 1019.310 225.700 2898.170 ;
        RECT 225.500 1018.990 225.760 1019.310 ;
        RECT 781.640 1018.990 781.900 1019.310 ;
        RECT 781.700 999.330 781.840 1018.990 ;
        RECT 783.830 999.330 784.110 1000.000 ;
        RECT 781.700 999.190 784.110 999.330 ;
        RECT 783.830 996.000 784.110 999.190 ;
      LAYER via2 ;
        RECT 16.650 2899.720 16.930 2900.000 ;
      LAYER met3 ;
        RECT -4.800 2900.010 2.400 2900.460 ;
        RECT 16.625 2900.010 16.955 2900.025 ;
        RECT -4.800 2899.710 16.955 2900.010 ;
        RECT -4.800 2899.260 2.400 2899.710 ;
        RECT 16.625 2899.695 16.955 2899.710 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.790 2635.920 15.110 2635.980 ;
        RECT 800.470 2635.920 800.790 2635.980 ;
        RECT 14.790 2635.780 800.790 2635.920 ;
        RECT 14.790 2635.720 15.110 2635.780 ;
        RECT 800.470 2635.720 800.790 2635.780 ;
      LAYER via ;
        RECT 14.820 2635.720 15.080 2635.980 ;
        RECT 800.500 2635.720 800.760 2635.980 ;
      LAYER met2 ;
        RECT 14.810 2639.235 15.090 2639.605 ;
        RECT 14.880 2636.010 15.020 2639.235 ;
        RECT 14.820 2635.690 15.080 2636.010 ;
        RECT 800.500 2635.690 800.760 2636.010 ;
        RECT 800.560 1048.870 800.700 2635.690 ;
        RECT 800.560 1048.730 804.840 1048.870 ;
        RECT 804.700 999.330 804.840 1048.730 ;
        RECT 806.370 999.330 806.650 1000.000 ;
        RECT 804.700 999.190 806.650 999.330 ;
        RECT 806.370 996.000 806.650 999.190 ;
      LAYER via2 ;
        RECT 14.810 2639.280 15.090 2639.560 ;
      LAYER met3 ;
        RECT -4.800 2639.570 2.400 2640.020 ;
        RECT 14.785 2639.570 15.115 2639.585 ;
        RECT -4.800 2639.270 15.115 2639.570 ;
        RECT -4.800 2638.820 2.400 2639.270 ;
        RECT 14.785 2639.255 15.115 2639.270 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2373.780 15.570 2373.840 ;
        RECT 828.070 2373.780 828.390 2373.840 ;
        RECT 15.250 2373.640 828.390 2373.780 ;
        RECT 15.250 2373.580 15.570 2373.640 ;
        RECT 828.070 2373.580 828.390 2373.640 ;
      LAYER via ;
        RECT 15.280 2373.580 15.540 2373.840 ;
        RECT 828.100 2373.580 828.360 2373.840 ;
      LAYER met2 ;
        RECT 15.270 2378.115 15.550 2378.485 ;
        RECT 15.340 2373.870 15.480 2378.115 ;
        RECT 15.280 2373.550 15.540 2373.870 ;
        RECT 828.100 2373.550 828.360 2373.870 ;
        RECT 828.160 999.330 828.300 2373.550 ;
        RECT 828.450 999.330 828.730 1000.000 ;
        RECT 828.160 999.190 828.730 999.330 ;
        RECT 828.450 996.000 828.730 999.190 ;
      LAYER via2 ;
        RECT 15.270 2378.160 15.550 2378.440 ;
      LAYER met3 ;
        RECT -4.800 2378.450 2.400 2378.900 ;
        RECT 15.245 2378.450 15.575 2378.465 ;
        RECT -4.800 2378.150 15.575 2378.450 ;
        RECT -4.800 2377.700 2.400 2378.150 ;
        RECT 15.245 2378.135 15.575 2378.150 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2111.640 17.870 2111.700 ;
        RECT 848.770 2111.640 849.090 2111.700 ;
        RECT 17.550 2111.500 849.090 2111.640 ;
        RECT 17.550 2111.440 17.870 2111.500 ;
        RECT 848.770 2111.440 849.090 2111.500 ;
      LAYER via ;
        RECT 17.580 2111.440 17.840 2111.700 ;
        RECT 848.800 2111.440 849.060 2111.700 ;
      LAYER met2 ;
        RECT 17.570 2117.675 17.850 2118.045 ;
        RECT 17.640 2111.730 17.780 2117.675 ;
        RECT 17.580 2111.410 17.840 2111.730 ;
        RECT 848.800 2111.410 849.060 2111.730 ;
        RECT 848.860 999.330 849.000 2111.410 ;
        RECT 850.990 999.330 851.270 1000.000 ;
        RECT 848.860 999.190 851.270 999.330 ;
        RECT 850.990 996.000 851.270 999.190 ;
      LAYER via2 ;
        RECT 17.570 2117.720 17.850 2118.000 ;
      LAYER met3 ;
        RECT -4.800 2118.010 2.400 2118.460 ;
        RECT 17.545 2118.010 17.875 2118.025 ;
        RECT -4.800 2117.710 17.875 2118.010 ;
        RECT -4.800 2117.260 2.400 2117.710 ;
        RECT 17.545 2117.695 17.875 2117.710 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 249.850 1001.540 250.170 1001.600 ;
        RECT 2903.590 1001.540 2903.910 1001.600 ;
        RECT 249.850 1001.400 2903.910 1001.540 ;
        RECT 249.850 1001.340 250.170 1001.400 ;
        RECT 2903.590 1001.340 2903.910 1001.400 ;
      LAYER via ;
        RECT 249.880 1001.340 250.140 1001.600 ;
        RECT 2903.620 1001.340 2903.880 1001.600 ;
      LAYER met2 ;
        RECT 249.880 1001.310 250.140 1001.630 ;
        RECT 2903.620 1001.310 2903.880 1001.630 ;
        RECT 248.390 999.330 248.670 1000.000 ;
        RECT 249.940 999.330 250.080 1001.310 ;
        RECT 248.390 999.190 250.080 999.330 ;
        RECT 248.390 996.000 248.670 999.190 ;
        RECT 2903.680 430.965 2903.820 1001.310 ;
        RECT 2903.610 430.595 2903.890 430.965 ;
      LAYER via2 ;
        RECT 2903.610 430.640 2903.890 430.920 ;
      LAYER met3 ;
        RECT 2903.585 430.930 2903.915 430.945 ;
        RECT 2917.600 430.930 2924.800 431.380 ;
        RECT 2903.585 430.630 2924.800 430.930 ;
        RECT 2903.585 430.615 2903.915 430.630 ;
        RECT 2917.600 430.180 2924.800 430.630 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1856.300 17.870 1856.360 ;
        RECT 869.470 1856.300 869.790 1856.360 ;
        RECT 17.550 1856.160 869.790 1856.300 ;
        RECT 17.550 1856.100 17.870 1856.160 ;
        RECT 869.470 1856.100 869.790 1856.160 ;
      LAYER via ;
        RECT 17.580 1856.100 17.840 1856.360 ;
        RECT 869.500 1856.100 869.760 1856.360 ;
      LAYER met2 ;
        RECT 17.570 1856.555 17.850 1856.925 ;
        RECT 17.640 1856.390 17.780 1856.555 ;
        RECT 17.580 1856.070 17.840 1856.390 ;
        RECT 869.500 1856.070 869.760 1856.390 ;
        RECT 869.560 1048.870 869.700 1856.070 ;
        RECT 869.560 1048.730 871.080 1048.870 ;
        RECT 870.940 999.330 871.080 1048.730 ;
        RECT 873.070 999.330 873.350 1000.000 ;
        RECT 870.940 999.190 873.350 999.330 ;
        RECT 873.070 996.000 873.350 999.190 ;
      LAYER via2 ;
        RECT 17.570 1856.600 17.850 1856.880 ;
      LAYER met3 ;
        RECT -4.800 1856.890 2.400 1857.340 ;
        RECT 17.545 1856.890 17.875 1856.905 ;
        RECT -4.800 1856.590 17.875 1856.890 ;
        RECT -4.800 1856.140 2.400 1856.590 ;
        RECT 17.545 1856.575 17.875 1856.590 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1594.160 16.950 1594.220 ;
        RECT 890.170 1594.160 890.490 1594.220 ;
        RECT 16.630 1594.020 890.490 1594.160 ;
        RECT 16.630 1593.960 16.950 1594.020 ;
        RECT 890.170 1593.960 890.490 1594.020 ;
      LAYER via ;
        RECT 16.660 1593.960 16.920 1594.220 ;
        RECT 890.200 1593.960 890.460 1594.220 ;
      LAYER met2 ;
        RECT 16.650 1596.115 16.930 1596.485 ;
        RECT 16.720 1594.250 16.860 1596.115 ;
        RECT 16.660 1593.930 16.920 1594.250 ;
        RECT 890.200 1593.930 890.460 1594.250 ;
        RECT 890.260 1048.870 890.400 1593.930 ;
        RECT 890.260 1048.730 894.080 1048.870 ;
        RECT 893.940 999.330 894.080 1048.730 ;
        RECT 895.610 999.330 895.890 1000.000 ;
        RECT 893.940 999.190 895.890 999.330 ;
        RECT 895.610 996.000 895.890 999.190 ;
      LAYER via2 ;
        RECT 16.650 1596.160 16.930 1596.440 ;
      LAYER met3 ;
        RECT -4.800 1596.450 2.400 1596.900 ;
        RECT 16.625 1596.450 16.955 1596.465 ;
        RECT -4.800 1596.150 16.955 1596.450 ;
        RECT -4.800 1595.700 2.400 1596.150 ;
        RECT 16.625 1596.135 16.955 1596.150 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1332.020 17.870 1332.080 ;
        RECT 917.770 1332.020 918.090 1332.080 ;
        RECT 17.550 1331.880 918.090 1332.020 ;
        RECT 17.550 1331.820 17.870 1331.880 ;
        RECT 917.770 1331.820 918.090 1331.880 ;
      LAYER via ;
        RECT 17.580 1331.820 17.840 1332.080 ;
        RECT 917.800 1331.820 918.060 1332.080 ;
      LAYER met2 ;
        RECT 17.570 1335.675 17.850 1336.045 ;
        RECT 17.640 1332.110 17.780 1335.675 ;
        RECT 17.580 1331.790 17.840 1332.110 ;
        RECT 917.800 1331.790 918.060 1332.110 ;
        RECT 917.860 1048.870 918.000 1331.790 ;
        RECT 917.860 1048.730 918.460 1048.870 ;
        RECT 917.690 999.330 917.970 1000.000 ;
        RECT 918.320 999.330 918.460 1048.730 ;
        RECT 917.690 999.190 918.460 999.330 ;
        RECT 917.690 996.000 917.970 999.190 ;
      LAYER via2 ;
        RECT 17.570 1335.720 17.850 1336.000 ;
      LAYER met3 ;
        RECT -4.800 1336.010 2.400 1336.460 ;
        RECT 17.545 1336.010 17.875 1336.025 ;
        RECT -4.800 1335.710 17.875 1336.010 ;
        RECT -4.800 1335.260 2.400 1335.710 ;
        RECT 17.545 1335.695 17.875 1335.710 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1069.880 17.870 1069.940 ;
        RECT 927.890 1069.880 928.210 1069.940 ;
        RECT 17.550 1069.740 928.210 1069.880 ;
        RECT 17.550 1069.680 17.870 1069.740 ;
        RECT 927.890 1069.680 928.210 1069.740 ;
        RECT 927.890 1014.120 928.210 1014.180 ;
        RECT 938.470 1014.120 938.790 1014.180 ;
        RECT 927.890 1013.980 938.790 1014.120 ;
        RECT 927.890 1013.920 928.210 1013.980 ;
        RECT 938.470 1013.920 938.790 1013.980 ;
      LAYER via ;
        RECT 17.580 1069.680 17.840 1069.940 ;
        RECT 927.920 1069.680 928.180 1069.940 ;
        RECT 927.920 1013.920 928.180 1014.180 ;
        RECT 938.500 1013.920 938.760 1014.180 ;
      LAYER met2 ;
        RECT 17.570 1074.555 17.850 1074.925 ;
        RECT 17.640 1069.970 17.780 1074.555 ;
        RECT 17.580 1069.650 17.840 1069.970 ;
        RECT 927.920 1069.650 928.180 1069.970 ;
        RECT 927.980 1014.210 928.120 1069.650 ;
        RECT 927.920 1013.890 928.180 1014.210 ;
        RECT 938.500 1013.890 938.760 1014.210 ;
        RECT 938.560 999.330 938.700 1013.890 ;
        RECT 940.230 999.330 940.510 1000.000 ;
        RECT 938.560 999.190 940.510 999.330 ;
        RECT 940.230 996.000 940.510 999.190 ;
      LAYER via2 ;
        RECT 17.570 1074.600 17.850 1074.880 ;
      LAYER met3 ;
        RECT -4.800 1074.890 2.400 1075.340 ;
        RECT 17.545 1074.890 17.875 1074.905 ;
        RECT -4.800 1074.590 17.875 1074.890 ;
        RECT -4.800 1074.140 2.400 1074.590 ;
        RECT 17.545 1074.575 17.875 1074.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 927.890 1012.080 928.210 1012.140 ;
        RECT 960.550 1012.080 960.870 1012.140 ;
        RECT 927.890 1011.940 960.870 1012.080 ;
        RECT 927.890 1011.880 928.210 1011.940 ;
        RECT 960.550 1011.880 960.870 1011.940 ;
        RECT 15.710 1008.680 16.030 1008.740 ;
        RECT 927.890 1008.680 928.210 1008.740 ;
        RECT 15.710 1008.540 928.210 1008.680 ;
        RECT 15.710 1008.480 16.030 1008.540 ;
        RECT 927.890 1008.480 928.210 1008.540 ;
      LAYER via ;
        RECT 927.920 1011.880 928.180 1012.140 ;
        RECT 960.580 1011.880 960.840 1012.140 ;
        RECT 15.740 1008.480 16.000 1008.740 ;
        RECT 927.920 1008.480 928.180 1008.740 ;
      LAYER met2 ;
        RECT 927.920 1011.850 928.180 1012.170 ;
        RECT 960.580 1011.850 960.840 1012.170 ;
        RECT 927.980 1008.770 928.120 1011.850 ;
        RECT 15.740 1008.450 16.000 1008.770 ;
        RECT 927.920 1008.450 928.180 1008.770 ;
        RECT 15.800 814.485 15.940 1008.450 ;
        RECT 960.640 999.330 960.780 1011.850 ;
        RECT 962.310 999.330 962.590 1000.000 ;
        RECT 960.640 999.190 962.590 999.330 ;
        RECT 962.310 996.000 962.590 999.190 ;
        RECT 15.730 814.115 16.010 814.485 ;
      LAYER via2 ;
        RECT 15.730 814.160 16.010 814.440 ;
      LAYER met3 ;
        RECT -4.800 814.450 2.400 814.900 ;
        RECT 15.705 814.450 16.035 814.465 ;
        RECT -4.800 814.150 16.035 814.450 ;
        RECT -4.800 813.700 2.400 814.150 ;
        RECT 15.705 814.135 16.035 814.150 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1008.340 16.950 1008.400 ;
        RECT 983.550 1008.340 983.870 1008.400 ;
        RECT 16.630 1008.200 983.870 1008.340 ;
        RECT 16.630 1008.140 16.950 1008.200 ;
        RECT 983.550 1008.140 983.870 1008.200 ;
      LAYER via ;
        RECT 16.660 1008.140 16.920 1008.400 ;
        RECT 983.580 1008.140 983.840 1008.400 ;
      LAYER met2 ;
        RECT 16.660 1008.110 16.920 1008.430 ;
        RECT 983.580 1008.110 983.840 1008.430 ;
        RECT 16.720 553.365 16.860 1008.110 ;
        RECT 983.640 999.330 983.780 1008.110 ;
        RECT 984.850 999.330 985.130 1000.000 ;
        RECT 983.640 999.190 985.130 999.330 ;
        RECT 984.850 996.000 985.130 999.190 ;
        RECT 16.650 552.995 16.930 553.365 ;
      LAYER via2 ;
        RECT 16.650 553.040 16.930 553.320 ;
      LAYER met3 ;
        RECT -4.800 553.330 2.400 553.780 ;
        RECT 16.625 553.330 16.955 553.345 ;
        RECT -4.800 553.030 16.955 553.330 ;
        RECT -4.800 552.580 2.400 553.030 ;
        RECT 16.625 553.015 16.955 553.030 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 217.650 998.140 217.970 998.200 ;
        RECT 228.690 998.140 229.010 998.200 ;
        RECT 217.650 998.000 229.010 998.140 ;
        RECT 217.650 997.940 217.970 998.000 ;
        RECT 228.690 997.940 229.010 998.000 ;
        RECT 217.650 997.460 217.970 997.520 ;
        RECT 213.830 997.320 217.970 997.460 ;
        RECT 19.390 994.740 19.710 994.800 ;
        RECT 19.390 994.600 131.170 994.740 ;
        RECT 19.390 994.540 19.710 994.600 ;
        RECT 131.030 994.060 131.170 994.600 ;
        RECT 131.030 993.920 179.470 994.060 ;
        RECT 179.330 993.380 179.470 993.920 ;
        RECT 179.330 993.240 186.370 993.380 ;
        RECT 186.230 992.360 186.370 993.240 ;
        RECT 213.830 992.360 213.970 997.320 ;
        RECT 217.650 997.260 217.970 997.320 ;
        RECT 228.690 997.260 229.010 997.520 ;
        RECT 280.670 997.460 280.990 997.520 ;
        RECT 265.580 997.320 280.990 997.460 ;
        RECT 228.780 996.440 228.920 997.260 ;
        RECT 265.580 996.440 265.720 997.320 ;
        RECT 280.670 997.260 280.990 997.320 ;
        RECT 281.590 997.460 281.910 997.520 ;
        RECT 1005.630 997.460 1005.950 997.520 ;
        RECT 281.590 997.320 303.670 997.460 ;
        RECT 281.590 997.260 281.910 997.320 ;
        RECT 228.780 996.300 265.720 996.440 ;
        RECT 303.530 996.440 303.670 997.320 ;
        RECT 1000.430 997.320 1005.950 997.460 ;
        RECT 303.530 996.300 309.880 996.440 ;
        RECT 309.740 994.740 309.880 996.300 ;
        RECT 1000.430 994.740 1000.570 997.320 ;
        RECT 1005.630 997.260 1005.950 997.320 ;
        RECT 309.740 994.600 1000.570 994.740 ;
        RECT 186.230 992.220 213.970 992.360 ;
      LAYER via ;
        RECT 217.680 997.940 217.940 998.200 ;
        RECT 228.720 997.940 228.980 998.200 ;
        RECT 19.420 994.540 19.680 994.800 ;
        RECT 217.680 997.260 217.940 997.520 ;
        RECT 228.720 997.260 228.980 997.520 ;
        RECT 280.700 997.260 280.960 997.520 ;
        RECT 281.620 997.260 281.880 997.520 ;
        RECT 1005.660 997.260 1005.920 997.520 ;
      LAYER met2 ;
        RECT 280.760 998.510 281.820 998.650 ;
        RECT 217.680 997.910 217.940 998.230 ;
        RECT 228.720 997.910 228.980 998.230 ;
        RECT 217.740 997.550 217.880 997.910 ;
        RECT 228.780 997.550 228.920 997.910 ;
        RECT 280.760 997.550 280.900 998.510 ;
        RECT 281.680 997.550 281.820 998.510 ;
        RECT 217.680 997.230 217.940 997.550 ;
        RECT 228.720 997.230 228.980 997.550 ;
        RECT 280.700 997.230 280.960 997.550 ;
        RECT 281.620 997.230 281.880 997.550 ;
        RECT 1005.660 997.290 1005.920 997.550 ;
        RECT 1006.930 997.290 1007.210 1000.000 ;
        RECT 1005.660 997.230 1007.210 997.290 ;
        RECT 1005.720 997.150 1007.210 997.230 ;
        RECT 1006.930 996.000 1007.210 997.150 ;
        RECT 19.420 994.510 19.680 994.830 ;
        RECT 19.480 358.205 19.620 994.510 ;
        RECT 19.410 357.835 19.690 358.205 ;
      LAYER via2 ;
        RECT 19.410 357.880 19.690 358.160 ;
      LAYER met3 ;
        RECT -4.800 358.170 2.400 358.620 ;
        RECT 19.385 358.170 19.715 358.185 ;
        RECT -4.800 357.870 19.715 358.170 ;
        RECT -4.800 357.420 2.400 357.870 ;
        RECT 19.385 357.855 19.715 357.870 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1002.900 17.870 1002.960 ;
        RECT 1028.170 1002.900 1028.490 1002.960 ;
        RECT 17.550 1002.760 1028.490 1002.900 ;
        RECT 17.550 1002.700 17.870 1002.760 ;
        RECT 1028.170 1002.700 1028.490 1002.760 ;
      LAYER via ;
        RECT 17.580 1002.700 17.840 1002.960 ;
        RECT 1028.200 1002.700 1028.460 1002.960 ;
      LAYER met2 ;
        RECT 17.580 1002.670 17.840 1002.990 ;
        RECT 1028.200 1002.670 1028.460 1002.990 ;
        RECT 17.640 162.365 17.780 1002.670 ;
        RECT 1028.260 999.330 1028.400 1002.670 ;
        RECT 1029.470 999.330 1029.750 1000.000 ;
        RECT 1028.260 999.190 1029.750 999.330 ;
        RECT 1029.470 996.000 1029.750 999.190 ;
        RECT 17.570 161.995 17.850 162.365 ;
      LAYER via2 ;
        RECT 17.570 162.040 17.850 162.320 ;
      LAYER met3 ;
        RECT -4.800 162.330 2.400 162.780 ;
        RECT 17.545 162.330 17.875 162.345 ;
        RECT -4.800 162.030 17.875 162.330 ;
        RECT -4.800 161.580 2.400 162.030 ;
        RECT 17.545 162.015 17.875 162.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 271.930 1009.700 272.250 1009.760 ;
        RECT 1100.850 1009.700 1101.170 1009.760 ;
        RECT 271.930 1009.560 1101.170 1009.700 ;
        RECT 271.930 1009.500 272.250 1009.560 ;
        RECT 1100.850 1009.500 1101.170 1009.560 ;
        RECT 1100.850 634.680 1101.170 634.740 ;
        RECT 2899.910 634.680 2900.230 634.740 ;
        RECT 1100.850 634.540 2900.230 634.680 ;
        RECT 1100.850 634.480 1101.170 634.540 ;
        RECT 2899.910 634.480 2900.230 634.540 ;
      LAYER via ;
        RECT 271.960 1009.500 272.220 1009.760 ;
        RECT 1100.880 1009.500 1101.140 1009.760 ;
        RECT 1100.880 634.480 1101.140 634.740 ;
        RECT 2899.940 634.480 2900.200 634.740 ;
      LAYER met2 ;
        RECT 271.960 1009.470 272.220 1009.790 ;
        RECT 1100.880 1009.470 1101.140 1009.790 ;
        RECT 270.470 999.330 270.750 1000.000 ;
        RECT 272.020 999.330 272.160 1009.470 ;
        RECT 270.470 999.190 272.160 999.330 ;
        RECT 270.470 996.000 270.750 999.190 ;
        RECT 1100.940 634.770 1101.080 1009.470 ;
        RECT 1100.880 634.450 1101.140 634.770 ;
        RECT 2899.940 634.450 2900.200 634.770 ;
        RECT 2900.000 630.205 2900.140 634.450 ;
        RECT 2899.930 629.835 2900.210 630.205 ;
      LAYER via2 ;
        RECT 2899.930 629.880 2900.210 630.160 ;
      LAYER met3 ;
        RECT 2899.905 630.170 2900.235 630.185 ;
        RECT 2917.600 630.170 2924.800 630.620 ;
        RECT 2899.905 629.870 2924.800 630.170 ;
        RECT 2899.905 629.855 2900.235 629.870 ;
        RECT 2917.600 629.420 2924.800 629.870 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.930 1010.720 295.250 1010.780 ;
        RECT 1102.230 1010.720 1102.550 1010.780 ;
        RECT 294.930 1010.580 1102.550 1010.720 ;
        RECT 294.930 1010.520 295.250 1010.580 ;
        RECT 1102.230 1010.520 1102.550 1010.580 ;
        RECT 1102.230 834.940 1102.550 835.000 ;
        RECT 2900.830 834.940 2901.150 835.000 ;
        RECT 1102.230 834.800 2901.150 834.940 ;
        RECT 1102.230 834.740 1102.550 834.800 ;
        RECT 2900.830 834.740 2901.150 834.800 ;
      LAYER via ;
        RECT 294.960 1010.520 295.220 1010.780 ;
        RECT 1102.260 1010.520 1102.520 1010.780 ;
        RECT 1102.260 834.740 1102.520 835.000 ;
        RECT 2900.860 834.740 2901.120 835.000 ;
      LAYER met2 ;
        RECT 294.960 1010.490 295.220 1010.810 ;
        RECT 1102.260 1010.490 1102.520 1010.810 ;
        RECT 293.010 999.330 293.290 1000.000 ;
        RECT 295.020 999.330 295.160 1010.490 ;
        RECT 293.010 999.190 295.160 999.330 ;
        RECT 293.010 996.000 293.290 999.190 ;
        RECT 1102.320 835.030 1102.460 1010.490 ;
        RECT 1102.260 834.710 1102.520 835.030 ;
        RECT 2900.860 834.710 2901.120 835.030 ;
        RECT 2900.920 829.445 2901.060 834.710 ;
        RECT 2900.850 829.075 2901.130 829.445 ;
      LAYER via2 ;
        RECT 2900.850 829.120 2901.130 829.400 ;
      LAYER met3 ;
        RECT 2900.825 829.410 2901.155 829.425 ;
        RECT 2917.600 829.410 2924.800 829.860 ;
        RECT 2900.825 829.110 2924.800 829.410 ;
        RECT 2900.825 829.095 2901.155 829.110 ;
        RECT 2917.600 828.660 2924.800 829.110 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 313.330 1028.400 313.650 1028.460 ;
        RECT 2900.830 1028.400 2901.150 1028.460 ;
        RECT 313.330 1028.260 2901.150 1028.400 ;
        RECT 313.330 1028.200 313.650 1028.260 ;
        RECT 2900.830 1028.200 2901.150 1028.260 ;
      LAYER via ;
        RECT 313.360 1028.200 313.620 1028.460 ;
        RECT 2900.860 1028.200 2901.120 1028.460 ;
      LAYER met2 ;
        RECT 313.360 1028.170 313.620 1028.490 ;
        RECT 2900.850 1028.315 2901.130 1028.685 ;
        RECT 2900.860 1028.170 2901.120 1028.315 ;
        RECT 313.420 999.330 313.560 1028.170 ;
        RECT 315.090 999.330 315.370 1000.000 ;
        RECT 313.420 999.190 315.370 999.330 ;
        RECT 315.090 996.000 315.370 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1028.360 2901.130 1028.640 ;
      LAYER met3 ;
        RECT 2900.825 1028.650 2901.155 1028.665 ;
        RECT 2917.600 1028.650 2924.800 1029.100 ;
        RECT 2900.825 1028.350 2924.800 1028.650 ;
        RECT 2900.825 1028.335 2901.155 1028.350 ;
        RECT 2917.600 1027.900 2924.800 1028.350 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 1221.520 331.590 1221.580 ;
        RECT 2898.990 1221.520 2899.310 1221.580 ;
        RECT 331.270 1221.380 2899.310 1221.520 ;
        RECT 331.270 1221.320 331.590 1221.380 ;
        RECT 2898.990 1221.320 2899.310 1221.380 ;
      LAYER via ;
        RECT 331.300 1221.320 331.560 1221.580 ;
        RECT 2899.020 1221.320 2899.280 1221.580 ;
      LAYER met2 ;
        RECT 2899.010 1227.555 2899.290 1227.925 ;
        RECT 2899.080 1221.610 2899.220 1227.555 ;
        RECT 331.300 1221.290 331.560 1221.610 ;
        RECT 2899.020 1221.290 2899.280 1221.610 ;
        RECT 331.360 1048.870 331.500 1221.290 ;
        RECT 331.360 1048.730 335.640 1048.870 ;
        RECT 335.500 999.330 335.640 1048.730 ;
        RECT 337.630 999.330 337.910 1000.000 ;
        RECT 335.500 999.190 337.910 999.330 ;
        RECT 337.630 996.000 337.910 999.190 ;
      LAYER via2 ;
        RECT 2899.010 1227.600 2899.290 1227.880 ;
      LAYER met3 ;
        RECT 2898.985 1227.890 2899.315 1227.905 ;
        RECT 2917.600 1227.890 2924.800 1228.340 ;
        RECT 2898.985 1227.590 2924.800 1227.890 ;
        RECT 2898.985 1227.575 2899.315 1227.590 ;
        RECT 2917.600 1227.140 2924.800 1227.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.330 1490.800 359.650 1490.860 ;
        RECT 2900.830 1490.800 2901.150 1490.860 ;
        RECT 359.330 1490.660 2901.150 1490.800 ;
        RECT 359.330 1490.600 359.650 1490.660 ;
        RECT 2900.830 1490.600 2901.150 1490.660 ;
      LAYER via ;
        RECT 359.360 1490.600 359.620 1490.860 ;
        RECT 2900.860 1490.600 2901.120 1490.860 ;
      LAYER met2 ;
        RECT 2900.850 1493.435 2901.130 1493.805 ;
        RECT 2900.920 1490.890 2901.060 1493.435 ;
        RECT 359.360 1490.570 359.620 1490.890 ;
        RECT 2900.860 1490.570 2901.120 1490.890 ;
        RECT 359.420 999.330 359.560 1490.570 ;
        RECT 359.710 999.330 359.990 1000.000 ;
        RECT 359.420 999.190 359.990 999.330 ;
        RECT 359.710 996.000 359.990 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1493.480 2901.130 1493.760 ;
      LAYER met3 ;
        RECT 2900.825 1493.770 2901.155 1493.785 ;
        RECT 2917.600 1493.770 2924.800 1494.220 ;
        RECT 2900.825 1493.470 2924.800 1493.770 ;
        RECT 2900.825 1493.455 2901.155 1493.470 ;
        RECT 2917.600 1493.020 2924.800 1493.470 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 379.570 1759.740 379.890 1759.800 ;
        RECT 2900.830 1759.740 2901.150 1759.800 ;
        RECT 379.570 1759.600 2901.150 1759.740 ;
        RECT 379.570 1759.540 379.890 1759.600 ;
        RECT 2900.830 1759.540 2901.150 1759.600 ;
      LAYER via ;
        RECT 379.600 1759.540 379.860 1759.800 ;
        RECT 2900.860 1759.540 2901.120 1759.800 ;
      LAYER met2 ;
        RECT 379.600 1759.510 379.860 1759.830 ;
        RECT 2900.860 1759.685 2901.120 1759.830 ;
        RECT 379.660 1048.870 379.800 1759.510 ;
        RECT 2900.850 1759.315 2901.130 1759.685 ;
        RECT 379.660 1048.730 380.720 1048.870 ;
        RECT 380.580 999.330 380.720 1048.730 ;
        RECT 382.250 999.330 382.530 1000.000 ;
        RECT 380.580 999.190 382.530 999.330 ;
        RECT 382.250 996.000 382.530 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1759.360 2901.130 1759.640 ;
      LAYER met3 ;
        RECT 2900.825 1759.650 2901.155 1759.665 ;
        RECT 2917.600 1759.650 2924.800 1760.100 ;
        RECT 2900.825 1759.350 2924.800 1759.650 ;
        RECT 2900.825 1759.335 2901.155 1759.350 ;
        RECT 2917.600 1758.900 2924.800 1759.350 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 2021.880 400.590 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 400.270 2021.740 2901.150 2021.880 ;
        RECT 400.270 2021.680 400.590 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 400.300 2021.680 400.560 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2024.515 2901.130 2024.885 ;
        RECT 2900.920 2021.970 2901.060 2024.515 ;
        RECT 400.300 2021.650 400.560 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 400.360 1048.870 400.500 2021.650 ;
        RECT 400.360 1048.730 402.800 1048.870 ;
        RECT 402.660 999.330 402.800 1048.730 ;
        RECT 404.330 999.330 404.610 1000.000 ;
        RECT 402.660 999.190 404.610 999.330 ;
        RECT 404.330 996.000 404.610 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2024.560 2901.130 2024.840 ;
      LAYER met3 ;
        RECT 2900.825 2024.850 2901.155 2024.865 ;
        RECT 2917.600 2024.850 2924.800 2025.300 ;
        RECT 2900.825 2024.550 2924.800 2024.850 ;
        RECT 2900.825 2024.535 2901.155 2024.550 ;
        RECT 2917.600 2024.100 2924.800 2024.550 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 213.050 1000.860 213.370 1000.920 ;
        RECT 2901.750 1000.860 2902.070 1000.920 ;
        RECT 213.050 1000.720 2902.070 1000.860 ;
        RECT 213.050 1000.660 213.370 1000.720 ;
        RECT 2901.750 1000.660 2902.070 1000.720 ;
      LAYER via ;
        RECT 213.080 1000.660 213.340 1000.920 ;
        RECT 2901.780 1000.660 2902.040 1000.920 ;
      LAYER met2 ;
        RECT 213.080 1000.630 213.340 1000.950 ;
        RECT 2901.780 1000.630 2902.040 1000.950 ;
        RECT 211.130 999.330 211.410 1000.000 ;
        RECT 213.140 999.330 213.280 1000.630 ;
        RECT 211.130 999.190 213.280 999.330 ;
        RECT 211.130 996.000 211.410 999.190 ;
        RECT 2901.840 165.765 2901.980 1000.630 ;
        RECT 2901.770 165.395 2902.050 165.765 ;
      LAYER via2 ;
        RECT 2901.770 165.440 2902.050 165.720 ;
      LAYER met3 ;
        RECT 2901.745 165.730 2902.075 165.745 ;
        RECT 2917.600 165.730 2924.800 166.180 ;
        RECT 2901.745 165.430 2924.800 165.730 ;
        RECT 2901.745 165.415 2902.075 165.430 ;
        RECT 2917.600 164.980 2924.800 165.430 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 2422.060 428.190 2422.120 ;
        RECT 2900.830 2422.060 2901.150 2422.120 ;
        RECT 427.870 2421.920 2901.150 2422.060 ;
        RECT 427.870 2421.860 428.190 2421.920 ;
        RECT 2900.830 2421.860 2901.150 2421.920 ;
      LAYER via ;
        RECT 427.900 2421.860 428.160 2422.120 ;
        RECT 2900.860 2421.860 2901.120 2422.120 ;
      LAYER met2 ;
        RECT 2900.850 2422.995 2901.130 2423.365 ;
        RECT 2900.920 2422.150 2901.060 2422.995 ;
        RECT 427.900 2421.830 428.160 2422.150 ;
        RECT 2900.860 2421.830 2901.120 2422.150 ;
        RECT 427.960 1048.870 428.100 2421.830 ;
        RECT 427.960 1048.730 432.240 1048.870 ;
        RECT 432.100 999.330 432.240 1048.730 ;
        RECT 434.230 999.330 434.510 1000.000 ;
        RECT 432.100 999.190 434.510 999.330 ;
        RECT 434.230 996.000 434.510 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2423.040 2901.130 2423.320 ;
      LAYER met3 ;
        RECT 2900.825 2423.330 2901.155 2423.345 ;
        RECT 2917.600 2423.330 2924.800 2423.780 ;
        RECT 2900.825 2423.030 2924.800 2423.330 ;
        RECT 2900.825 2423.015 2901.155 2423.030 ;
        RECT 2917.600 2422.580 2924.800 2423.030 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 2684.200 455.790 2684.260 ;
        RECT 2900.830 2684.200 2901.150 2684.260 ;
        RECT 455.470 2684.060 2901.150 2684.200 ;
        RECT 455.470 2684.000 455.790 2684.060 ;
        RECT 2900.830 2684.000 2901.150 2684.060 ;
      LAYER via ;
        RECT 455.500 2684.000 455.760 2684.260 ;
        RECT 2900.860 2684.000 2901.120 2684.260 ;
      LAYER met2 ;
        RECT 2900.850 2688.875 2901.130 2689.245 ;
        RECT 2900.920 2684.290 2901.060 2688.875 ;
        RECT 455.500 2683.970 455.760 2684.290 ;
        RECT 2900.860 2683.970 2901.120 2684.290 ;
        RECT 455.560 999.330 455.700 2683.970 ;
        RECT 456.310 999.330 456.590 1000.000 ;
        RECT 455.560 999.190 456.590 999.330 ;
        RECT 456.310 996.000 456.590 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2688.920 2901.130 2689.200 ;
      LAYER met3 ;
        RECT 2900.825 2689.210 2901.155 2689.225 ;
        RECT 2917.600 2689.210 2924.800 2689.660 ;
        RECT 2900.825 2688.910 2924.800 2689.210 ;
        RECT 2900.825 2688.895 2901.155 2688.910 ;
        RECT 2917.600 2688.460 2924.800 2688.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 2953.480 476.490 2953.540 ;
        RECT 2898.990 2953.480 2899.310 2953.540 ;
        RECT 476.170 2953.340 2899.310 2953.480 ;
        RECT 476.170 2953.280 476.490 2953.340 ;
        RECT 2898.990 2953.280 2899.310 2953.340 ;
      LAYER via ;
        RECT 476.200 2953.280 476.460 2953.540 ;
        RECT 2899.020 2953.280 2899.280 2953.540 ;
      LAYER met2 ;
        RECT 2899.010 2954.755 2899.290 2955.125 ;
        RECT 2899.080 2953.570 2899.220 2954.755 ;
        RECT 476.200 2953.250 476.460 2953.570 ;
        RECT 2899.020 2953.250 2899.280 2953.570 ;
        RECT 476.260 1048.870 476.400 2953.250 ;
        RECT 476.260 1048.730 477.320 1048.870 ;
        RECT 477.180 999.330 477.320 1048.730 ;
        RECT 478.850 999.330 479.130 1000.000 ;
        RECT 477.180 999.190 479.130 999.330 ;
        RECT 478.850 996.000 479.130 999.190 ;
      LAYER via2 ;
        RECT 2899.010 2954.800 2899.290 2955.080 ;
      LAYER met3 ;
        RECT 2898.985 2955.090 2899.315 2955.105 ;
        RECT 2917.600 2955.090 2924.800 2955.540 ;
        RECT 2898.985 2954.790 2924.800 2955.090 ;
        RECT 2898.985 2954.775 2899.315 2954.790 ;
        RECT 2917.600 2954.340 2924.800 2954.790 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 3215.620 497.190 3215.680 ;
        RECT 2900.830 3215.620 2901.150 3215.680 ;
        RECT 496.870 3215.480 2901.150 3215.620 ;
        RECT 496.870 3215.420 497.190 3215.480 ;
        RECT 2900.830 3215.420 2901.150 3215.480 ;
      LAYER via ;
        RECT 496.900 3215.420 497.160 3215.680 ;
        RECT 2900.860 3215.420 2901.120 3215.680 ;
      LAYER met2 ;
        RECT 2900.850 3219.955 2901.130 3220.325 ;
        RECT 2900.920 3215.710 2901.060 3219.955 ;
        RECT 496.900 3215.390 497.160 3215.710 ;
        RECT 2900.860 3215.390 2901.120 3215.710 ;
        RECT 496.960 1048.870 497.100 3215.390 ;
        RECT 496.960 1048.730 499.400 1048.870 ;
        RECT 499.260 999.330 499.400 1048.730 ;
        RECT 500.930 999.330 501.210 1000.000 ;
        RECT 499.260 999.190 501.210 999.330 ;
        RECT 500.930 996.000 501.210 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3220.000 2901.130 3220.280 ;
      LAYER met3 ;
        RECT 2900.825 3220.290 2901.155 3220.305 ;
        RECT 2917.600 3220.290 2924.800 3220.740 ;
        RECT 2900.825 3219.990 2924.800 3220.290 ;
        RECT 2900.825 3219.975 2901.155 3219.990 ;
        RECT 2917.600 3219.540 2924.800 3219.990 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 3484.900 517.890 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 517.570 3484.760 2901.150 3484.900 ;
        RECT 517.570 3484.700 517.890 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 517.600 3484.700 517.860 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3485.835 2901.130 3486.205 ;
        RECT 2900.920 3484.990 2901.060 3485.835 ;
        RECT 517.600 3484.670 517.860 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 517.660 1048.870 517.800 3484.670 ;
        RECT 517.660 1048.730 521.480 1048.870 ;
        RECT 521.340 999.330 521.480 1048.730 ;
        RECT 523.470 999.330 523.750 1000.000 ;
        RECT 521.340 999.190 523.750 999.330 ;
        RECT 523.470 996.000 523.750 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3485.880 2901.130 3486.160 ;
      LAYER met3 ;
        RECT 2900.825 3486.170 2901.155 3486.185 ;
        RECT 2917.600 3486.170 2924.800 3486.620 ;
        RECT 2900.825 3485.870 2924.800 3486.170 ;
        RECT 2900.825 3485.855 2901.155 3485.870 ;
        RECT 2917.600 3485.420 2924.800 3485.870 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1003.790 3502.580 1004.110 3502.640 ;
        RECT 2635.870 3502.580 2636.190 3502.640 ;
        RECT 1003.790 3502.440 2636.190 3502.580 ;
        RECT 1003.790 3502.380 1004.110 3502.440 ;
        RECT 2635.870 3502.380 2636.190 3502.440 ;
        RECT 545.170 1020.920 545.490 1020.980 ;
        RECT 1003.790 1020.920 1004.110 1020.980 ;
        RECT 545.170 1020.780 1004.110 1020.920 ;
        RECT 545.170 1020.720 545.490 1020.780 ;
        RECT 1003.790 1020.720 1004.110 1020.780 ;
      LAYER via ;
        RECT 1003.820 3502.380 1004.080 3502.640 ;
        RECT 2635.900 3502.380 2636.160 3502.640 ;
        RECT 545.200 1020.720 545.460 1020.980 ;
        RECT 1003.820 1020.720 1004.080 1020.980 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.670 2636.100 3517.600 ;
        RECT 1003.820 3502.350 1004.080 3502.670 ;
        RECT 2635.900 3502.350 2636.160 3502.670 ;
        RECT 1003.880 1021.010 1004.020 3502.350 ;
        RECT 545.200 1020.690 545.460 1021.010 ;
        RECT 1003.820 1020.690 1004.080 1021.010 ;
        RECT 545.260 999.330 545.400 1020.690 ;
        RECT 545.550 999.330 545.830 1000.000 ;
        RECT 545.260 999.190 545.830 999.330 ;
        RECT 545.550 996.000 545.830 999.190 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 3502.240 566.190 3502.300 ;
        RECT 2311.570 3502.240 2311.890 3502.300 ;
        RECT 565.870 3502.100 2311.890 3502.240 ;
        RECT 565.870 3502.040 566.190 3502.100 ;
        RECT 2311.570 3502.040 2311.890 3502.100 ;
      LAYER via ;
        RECT 565.900 3502.040 566.160 3502.300 ;
        RECT 2311.600 3502.040 2311.860 3502.300 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3502.330 2311.800 3517.600 ;
        RECT 565.900 3502.010 566.160 3502.330 ;
        RECT 2311.600 3502.010 2311.860 3502.330 ;
        RECT 565.960 1048.870 566.100 3502.010 ;
        RECT 565.960 1048.730 566.560 1048.870 ;
        RECT 566.420 999.330 566.560 1048.730 ;
        RECT 568.090 999.330 568.370 1000.000 ;
        RECT 566.420 999.190 568.370 999.330 ;
        RECT 568.090 996.000 568.370 999.190 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 3503.260 586.890 3503.320 ;
        RECT 1987.270 3503.260 1987.590 3503.320 ;
        RECT 586.570 3503.120 1987.590 3503.260 ;
        RECT 586.570 3503.060 586.890 3503.120 ;
        RECT 1987.270 3503.060 1987.590 3503.120 ;
      LAYER via ;
        RECT 586.600 3503.060 586.860 3503.320 ;
        RECT 1987.300 3503.060 1987.560 3503.320 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3503.350 1987.500 3517.600 ;
        RECT 586.600 3503.030 586.860 3503.350 ;
        RECT 1987.300 3503.030 1987.560 3503.350 ;
        RECT 586.660 1048.870 586.800 3503.030 ;
        RECT 586.660 1048.730 588.640 1048.870 ;
        RECT 588.500 999.330 588.640 1048.730 ;
        RECT 590.630 999.330 590.910 1000.000 ;
        RECT 588.500 999.190 590.910 999.330 ;
        RECT 590.630 996.000 590.910 999.190 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 3503.940 608.050 3504.000 ;
        RECT 1662.510 3503.940 1662.830 3504.000 ;
        RECT 607.730 3503.800 1662.830 3503.940 ;
        RECT 607.730 3503.740 608.050 3503.800 ;
        RECT 1662.510 3503.740 1662.830 3503.800 ;
      LAYER via ;
        RECT 607.760 3503.740 608.020 3504.000 ;
        RECT 1662.540 3503.740 1662.800 3504.000 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3504.030 1662.740 3517.600 ;
        RECT 607.760 3503.710 608.020 3504.030 ;
        RECT 1662.540 3503.710 1662.800 3504.030 ;
        RECT 607.820 1048.870 607.960 3503.710 ;
        RECT 607.820 1048.730 610.720 1048.870 ;
        RECT 610.580 999.330 610.720 1048.730 ;
        RECT 612.710 999.330 612.990 1000.000 ;
        RECT 610.580 999.190 612.990 999.330 ;
        RECT 612.710 996.000 612.990 999.190 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1004.710 3501.220 1005.030 3501.280 ;
        RECT 1338.210 3501.220 1338.530 3501.280 ;
        RECT 1004.710 3501.080 1338.530 3501.220 ;
        RECT 1004.710 3501.020 1005.030 3501.080 ;
        RECT 1338.210 3501.020 1338.530 3501.080 ;
        RECT 634.870 1017.180 635.190 1017.240 ;
        RECT 1004.710 1017.180 1005.030 1017.240 ;
        RECT 634.870 1017.040 1005.030 1017.180 ;
        RECT 634.870 1016.980 635.190 1017.040 ;
        RECT 1004.710 1016.980 1005.030 1017.040 ;
      LAYER via ;
        RECT 1004.740 3501.020 1005.000 3501.280 ;
        RECT 1338.240 3501.020 1338.500 3501.280 ;
        RECT 634.900 1016.980 635.160 1017.240 ;
        RECT 1004.740 1016.980 1005.000 1017.240 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3501.310 1338.440 3517.600 ;
        RECT 1004.740 3500.990 1005.000 3501.310 ;
        RECT 1338.240 3500.990 1338.500 3501.310 ;
        RECT 1004.800 1017.270 1004.940 3500.990 ;
        RECT 634.900 1016.950 635.160 1017.270 ;
        RECT 1004.740 1016.950 1005.000 1017.270 ;
        RECT 634.960 999.330 635.100 1016.950 ;
        RECT 635.250 999.330 635.530 1000.000 ;
        RECT 634.960 999.190 635.530 999.330 ;
        RECT 635.250 996.000 635.530 999.190 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.210 1001.200 234.530 1001.260 ;
        RECT 2903.130 1001.200 2903.450 1001.260 ;
        RECT 234.210 1001.060 2903.450 1001.200 ;
        RECT 234.210 1001.000 234.530 1001.060 ;
        RECT 2903.130 1001.000 2903.450 1001.060 ;
      LAYER via ;
        RECT 234.240 1001.000 234.500 1001.260 ;
        RECT 2903.160 1001.000 2903.420 1001.260 ;
      LAYER met2 ;
        RECT 234.240 1000.970 234.500 1001.290 ;
        RECT 2903.160 1000.970 2903.420 1001.290 ;
        RECT 233.210 999.330 233.490 1000.000 ;
        RECT 234.300 999.330 234.440 1000.970 ;
        RECT 233.210 999.190 234.440 999.330 ;
        RECT 233.210 996.000 233.490 999.190 ;
        RECT 2903.220 365.005 2903.360 1000.970 ;
        RECT 2903.150 364.635 2903.430 365.005 ;
      LAYER via2 ;
        RECT 2903.150 364.680 2903.430 364.960 ;
      LAYER met3 ;
        RECT 2903.125 364.970 2903.455 364.985 ;
        RECT 2917.600 364.970 2924.800 365.420 ;
        RECT 2903.125 364.670 2924.800 364.970 ;
        RECT 2903.125 364.655 2903.455 364.670 ;
        RECT 2917.600 364.220 2924.800 364.670 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1004.250 3498.500 1004.570 3498.560 ;
        RECT 1013.910 3498.500 1014.230 3498.560 ;
        RECT 1004.250 3498.360 1014.230 3498.500 ;
        RECT 1004.250 3498.300 1004.570 3498.360 ;
        RECT 1013.910 3498.300 1014.230 3498.360 ;
        RECT 655.570 1016.840 655.890 1016.900 ;
        RECT 1004.250 1016.840 1004.570 1016.900 ;
        RECT 655.570 1016.700 1004.570 1016.840 ;
        RECT 655.570 1016.640 655.890 1016.700 ;
        RECT 1004.250 1016.640 1004.570 1016.700 ;
      LAYER via ;
        RECT 1004.280 3498.300 1004.540 3498.560 ;
        RECT 1013.940 3498.300 1014.200 3498.560 ;
        RECT 655.600 1016.640 655.860 1016.900 ;
        RECT 1004.280 1016.640 1004.540 1016.900 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3498.590 1014.140 3517.600 ;
        RECT 1004.280 3498.270 1004.540 3498.590 ;
        RECT 1013.940 3498.270 1014.200 3498.590 ;
        RECT 1004.340 1016.930 1004.480 3498.270 ;
        RECT 655.600 1016.610 655.860 1016.930 ;
        RECT 1004.280 1016.610 1004.540 1016.930 ;
        RECT 655.660 999.330 655.800 1016.610 ;
        RECT 657.330 999.330 657.610 1000.000 ;
        RECT 655.660 999.190 657.610 999.330 ;
        RECT 657.330 996.000 657.610 999.190 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.260 3517.910 688.460 3518.050 ;
        RECT 683.260 1014.370 683.400 3517.910 ;
        RECT 688.320 3517.370 688.460 3517.910 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3517.370 689.380 3517.600 ;
        RECT 688.320 3517.230 689.380 3517.370 ;
        RECT 681.880 1014.230 683.400 1014.370 ;
        RECT 679.870 999.330 680.150 1000.000 ;
        RECT 681.880 999.330 682.020 1014.230 ;
        RECT 679.870 999.190 682.020 999.330 ;
        RECT 679.870 996.000 680.150 999.190 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 358.870 3515.160 359.190 3515.220 ;
        RECT 364.850 3515.160 365.170 3515.220 ;
        RECT 358.870 3515.020 365.170 3515.160 ;
        RECT 358.870 3514.960 359.190 3515.020 ;
        RECT 364.850 3514.960 365.170 3515.020 ;
        RECT 358.870 1011.740 359.190 1011.800 ;
        RECT 699.730 1011.740 700.050 1011.800 ;
        RECT 358.870 1011.600 700.050 1011.740 ;
        RECT 358.870 1011.540 359.190 1011.600 ;
        RECT 699.730 1011.540 700.050 1011.600 ;
      LAYER via ;
        RECT 358.900 3514.960 359.160 3515.220 ;
        RECT 364.880 3514.960 365.140 3515.220 ;
        RECT 358.900 1011.540 359.160 1011.800 ;
        RECT 699.760 1011.540 700.020 1011.800 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3515.250 365.080 3517.600 ;
        RECT 358.900 3514.930 359.160 3515.250 ;
        RECT 364.880 3514.930 365.140 3515.250 ;
        RECT 358.960 1011.830 359.100 3514.930 ;
        RECT 358.900 1011.510 359.160 1011.830 ;
        RECT 699.760 1011.510 700.020 1011.830 ;
        RECT 699.820 999.330 699.960 1011.510 ;
        RECT 701.950 999.330 702.230 1000.000 ;
        RECT 699.820 999.190 702.230 999.330 ;
        RECT 701.950 996.000 702.230 999.190 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 210.290 3501.560 210.610 3501.620 ;
        RECT 40.550 3501.420 210.610 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 210.290 3501.360 210.610 3501.420 ;
        RECT 210.290 1019.900 210.610 1019.960 ;
        RECT 725.030 1019.900 725.350 1019.960 ;
        RECT 210.290 1019.760 725.350 1019.900 ;
        RECT 210.290 1019.700 210.610 1019.760 ;
        RECT 725.030 1019.700 725.350 1019.760 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 210.320 3501.360 210.580 3501.620 ;
        RECT 210.320 1019.700 210.580 1019.960 ;
        RECT 725.060 1019.700 725.320 1019.960 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.650 40.780 3517.600 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 210.320 3501.330 210.580 3501.650 ;
        RECT 210.380 1019.990 210.520 3501.330 ;
        RECT 210.320 1019.670 210.580 1019.990 ;
        RECT 725.060 1019.670 725.320 1019.990 ;
        RECT 724.490 999.330 724.770 1000.000 ;
        RECT 725.120 999.330 725.260 1019.670 ;
        RECT 724.490 999.190 725.260 999.330 ;
        RECT 724.490 996.000 724.770 999.190 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3284.980 17.870 3285.040 ;
        RECT 745.270 3284.980 745.590 3285.040 ;
        RECT 17.550 3284.840 745.590 3284.980 ;
        RECT 17.550 3284.780 17.870 3284.840 ;
        RECT 745.270 3284.780 745.590 3284.840 ;
      LAYER via ;
        RECT 17.580 3284.780 17.840 3285.040 ;
        RECT 745.300 3284.780 745.560 3285.040 ;
      LAYER met2 ;
        RECT 17.570 3290.675 17.850 3291.045 ;
        RECT 17.640 3285.070 17.780 3290.675 ;
        RECT 17.580 3284.750 17.840 3285.070 ;
        RECT 745.300 3284.750 745.560 3285.070 ;
        RECT 745.360 999.330 745.500 3284.750 ;
        RECT 746.570 999.330 746.850 1000.000 ;
        RECT 745.360 999.190 746.850 999.330 ;
        RECT 746.570 996.000 746.850 999.190 ;
      LAYER via2 ;
        RECT 17.570 3290.720 17.850 3291.000 ;
      LAYER met3 ;
        RECT -4.800 3291.010 2.400 3291.460 ;
        RECT 17.545 3291.010 17.875 3291.025 ;
        RECT -4.800 3290.710 17.875 3291.010 ;
        RECT -4.800 3290.260 2.400 3290.710 ;
        RECT 17.545 3290.695 17.875 3290.710 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3029.300 17.870 3029.360 ;
        RECT 765.970 3029.300 766.290 3029.360 ;
        RECT 17.550 3029.160 766.290 3029.300 ;
        RECT 17.550 3029.100 17.870 3029.160 ;
        RECT 765.970 3029.100 766.290 3029.160 ;
      LAYER via ;
        RECT 17.580 3029.100 17.840 3029.360 ;
        RECT 766.000 3029.100 766.260 3029.360 ;
      LAYER met2 ;
        RECT 17.570 3030.235 17.850 3030.605 ;
        RECT 17.640 3029.390 17.780 3030.235 ;
        RECT 17.580 3029.070 17.840 3029.390 ;
        RECT 766.000 3029.070 766.260 3029.390 ;
        RECT 766.060 1048.870 766.200 3029.070 ;
        RECT 766.060 1048.730 767.120 1048.870 ;
        RECT 766.980 999.330 767.120 1048.730 ;
        RECT 769.110 999.330 769.390 1000.000 ;
        RECT 766.980 999.190 769.390 999.330 ;
        RECT 769.110 996.000 769.390 999.190 ;
      LAYER via2 ;
        RECT 17.570 3030.280 17.850 3030.560 ;
      LAYER met3 ;
        RECT -4.800 3030.570 2.400 3031.020 ;
        RECT 17.545 3030.570 17.875 3030.585 ;
        RECT -4.800 3030.270 17.875 3030.570 ;
        RECT -4.800 3029.820 2.400 3030.270 ;
        RECT 17.545 3030.255 17.875 3030.270 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 2767.160 16.950 2767.220 ;
        RECT 786.670 2767.160 786.990 2767.220 ;
        RECT 16.630 2767.020 786.990 2767.160 ;
        RECT 16.630 2766.960 16.950 2767.020 ;
        RECT 786.670 2766.960 786.990 2767.020 ;
      LAYER via ;
        RECT 16.660 2766.960 16.920 2767.220 ;
        RECT 786.700 2766.960 786.960 2767.220 ;
      LAYER met2 ;
        RECT 16.650 2769.115 16.930 2769.485 ;
        RECT 16.720 2767.250 16.860 2769.115 ;
        RECT 16.660 2766.930 16.920 2767.250 ;
        RECT 786.700 2766.930 786.960 2767.250 ;
        RECT 786.760 1048.870 786.900 2766.930 ;
        RECT 786.760 1048.730 789.200 1048.870 ;
        RECT 789.060 999.330 789.200 1048.730 ;
        RECT 791.190 999.330 791.470 1000.000 ;
        RECT 789.060 999.190 791.470 999.330 ;
        RECT 791.190 996.000 791.470 999.190 ;
      LAYER via2 ;
        RECT 16.650 2769.160 16.930 2769.440 ;
      LAYER met3 ;
        RECT -4.800 2769.450 2.400 2769.900 ;
        RECT 16.625 2769.450 16.955 2769.465 ;
        RECT -4.800 2769.150 16.955 2769.450 ;
        RECT -4.800 2768.700 2.400 2769.150 ;
        RECT 16.625 2769.135 16.955 2769.150 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 2505.020 15.570 2505.080 ;
        RECT 807.370 2505.020 807.690 2505.080 ;
        RECT 15.250 2504.880 807.690 2505.020 ;
        RECT 15.250 2504.820 15.570 2504.880 ;
        RECT 807.370 2504.820 807.690 2504.880 ;
      LAYER via ;
        RECT 15.280 2504.820 15.540 2505.080 ;
        RECT 807.400 2504.820 807.660 2505.080 ;
      LAYER met2 ;
        RECT 15.270 2508.675 15.550 2509.045 ;
        RECT 15.340 2505.110 15.480 2508.675 ;
        RECT 15.280 2504.790 15.540 2505.110 ;
        RECT 807.400 2504.790 807.660 2505.110 ;
        RECT 807.460 1048.870 807.600 2504.790 ;
        RECT 807.460 1048.730 812.200 1048.870 ;
        RECT 812.060 999.330 812.200 1048.730 ;
        RECT 813.730 999.330 814.010 1000.000 ;
        RECT 812.060 999.190 814.010 999.330 ;
        RECT 813.730 996.000 814.010 999.190 ;
      LAYER via2 ;
        RECT 15.270 2508.720 15.550 2509.000 ;
      LAYER met3 ;
        RECT -4.800 2509.010 2.400 2509.460 ;
        RECT 15.245 2509.010 15.575 2509.025 ;
        RECT -4.800 2508.710 15.575 2509.010 ;
        RECT -4.800 2508.260 2.400 2508.710 ;
        RECT 15.245 2508.695 15.575 2508.710 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 2242.880 16.030 2242.940 ;
        RECT 834.970 2242.880 835.290 2242.940 ;
        RECT 15.710 2242.740 835.290 2242.880 ;
        RECT 15.710 2242.680 16.030 2242.740 ;
        RECT 834.970 2242.680 835.290 2242.740 ;
      LAYER via ;
        RECT 15.740 2242.680 16.000 2242.940 ;
        RECT 835.000 2242.680 835.260 2242.940 ;
      LAYER met2 ;
        RECT 15.730 2247.555 16.010 2247.925 ;
        RECT 15.800 2242.970 15.940 2247.555 ;
        RECT 15.740 2242.650 16.000 2242.970 ;
        RECT 835.000 2242.650 835.260 2242.970 ;
        RECT 835.060 999.330 835.200 2242.650 ;
        RECT 835.810 999.330 836.090 1000.000 ;
        RECT 835.060 999.190 836.090 999.330 ;
        RECT 835.810 996.000 836.090 999.190 ;
      LAYER via2 ;
        RECT 15.730 2247.600 16.010 2247.880 ;
      LAYER met3 ;
        RECT -4.800 2247.890 2.400 2248.340 ;
        RECT 15.705 2247.890 16.035 2247.905 ;
        RECT -4.800 2247.590 16.035 2247.890 ;
        RECT -4.800 2247.140 2.400 2247.590 ;
        RECT 15.705 2247.575 16.035 2247.590 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1987.540 17.870 1987.600 ;
        RECT 855.670 1987.540 855.990 1987.600 ;
        RECT 17.550 1987.400 855.990 1987.540 ;
        RECT 17.550 1987.340 17.870 1987.400 ;
        RECT 855.670 1987.340 855.990 1987.400 ;
      LAYER via ;
        RECT 17.580 1987.340 17.840 1987.600 ;
        RECT 855.700 1987.340 855.960 1987.600 ;
      LAYER met2 ;
        RECT 17.580 1987.485 17.840 1987.630 ;
        RECT 17.570 1987.115 17.850 1987.485 ;
        RECT 855.700 1987.310 855.960 1987.630 ;
        RECT 855.760 1048.870 855.900 1987.310 ;
        RECT 855.760 1048.730 856.360 1048.870 ;
        RECT 856.220 999.330 856.360 1048.730 ;
        RECT 858.350 999.330 858.630 1000.000 ;
        RECT 856.220 999.190 858.630 999.330 ;
        RECT 858.350 996.000 858.630 999.190 ;
      LAYER via2 ;
        RECT 17.570 1987.160 17.850 1987.440 ;
      LAYER met3 ;
        RECT -4.800 1987.450 2.400 1987.900 ;
        RECT 17.545 1987.450 17.875 1987.465 ;
        RECT -4.800 1987.150 17.875 1987.450 ;
        RECT -4.800 1986.700 2.400 1987.150 ;
        RECT 17.545 1987.135 17.875 1987.150 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 257.210 1001.880 257.530 1001.940 ;
        RECT 2904.050 1001.880 2904.370 1001.940 ;
        RECT 257.210 1001.740 2904.370 1001.880 ;
        RECT 257.210 1001.680 257.530 1001.740 ;
        RECT 2904.050 1001.680 2904.370 1001.740 ;
      LAYER via ;
        RECT 257.240 1001.680 257.500 1001.940 ;
        RECT 2904.080 1001.680 2904.340 1001.940 ;
      LAYER met2 ;
        RECT 257.240 1001.650 257.500 1001.970 ;
        RECT 2904.080 1001.650 2904.340 1001.970 ;
        RECT 255.750 999.330 256.030 1000.000 ;
        RECT 257.300 999.330 257.440 1001.650 ;
        RECT 255.750 999.190 257.440 999.330 ;
        RECT 255.750 996.000 256.030 999.190 ;
        RECT 2904.140 564.245 2904.280 1001.650 ;
        RECT 2904.070 563.875 2904.350 564.245 ;
      LAYER via2 ;
        RECT 2904.070 563.920 2904.350 564.200 ;
      LAYER met3 ;
        RECT 2904.045 564.210 2904.375 564.225 ;
        RECT 2917.600 564.210 2924.800 564.660 ;
        RECT 2904.045 563.910 2924.800 564.210 ;
        RECT 2904.045 563.895 2904.375 563.910 ;
        RECT 2917.600 563.460 2924.800 563.910 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1725.400 16.950 1725.460 ;
        RECT 876.370 1725.400 876.690 1725.460 ;
        RECT 16.630 1725.260 876.690 1725.400 ;
        RECT 16.630 1725.200 16.950 1725.260 ;
        RECT 876.370 1725.200 876.690 1725.260 ;
      LAYER via ;
        RECT 16.660 1725.200 16.920 1725.460 ;
        RECT 876.400 1725.200 876.660 1725.460 ;
      LAYER met2 ;
        RECT 16.650 1726.675 16.930 1727.045 ;
        RECT 16.720 1725.490 16.860 1726.675 ;
        RECT 16.660 1725.170 16.920 1725.490 ;
        RECT 876.400 1725.170 876.660 1725.490 ;
        RECT 876.460 1048.870 876.600 1725.170 ;
        RECT 876.460 1048.730 878.440 1048.870 ;
        RECT 878.300 999.330 878.440 1048.730 ;
        RECT 880.430 999.330 880.710 1000.000 ;
        RECT 878.300 999.190 880.710 999.330 ;
        RECT 880.430 996.000 880.710 999.190 ;
      LAYER via2 ;
        RECT 16.650 1726.720 16.930 1727.000 ;
      LAYER met3 ;
        RECT -4.800 1727.010 2.400 1727.460 ;
        RECT 16.625 1727.010 16.955 1727.025 ;
        RECT -4.800 1726.710 16.955 1727.010 ;
        RECT -4.800 1726.260 2.400 1726.710 ;
        RECT 16.625 1726.695 16.955 1726.710 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 1462.920 16.950 1462.980 ;
        RECT 700.190 1462.920 700.510 1462.980 ;
        RECT 16.630 1462.780 700.510 1462.920 ;
        RECT 16.630 1462.720 16.950 1462.780 ;
        RECT 700.190 1462.720 700.510 1462.780 ;
        RECT 700.190 1011.740 700.510 1011.800 ;
        RECT 899.830 1011.740 900.150 1011.800 ;
        RECT 700.190 1011.600 900.150 1011.740 ;
        RECT 700.190 1011.540 700.510 1011.600 ;
        RECT 899.830 1011.540 900.150 1011.600 ;
      LAYER via ;
        RECT 16.660 1462.720 16.920 1462.980 ;
        RECT 700.220 1462.720 700.480 1462.980 ;
        RECT 700.220 1011.540 700.480 1011.800 ;
        RECT 899.860 1011.540 900.120 1011.800 ;
      LAYER met2 ;
        RECT 16.650 1465.555 16.930 1465.925 ;
        RECT 16.720 1463.010 16.860 1465.555 ;
        RECT 16.660 1462.690 16.920 1463.010 ;
        RECT 700.220 1462.690 700.480 1463.010 ;
        RECT 700.280 1011.830 700.420 1462.690 ;
        RECT 700.220 1011.510 700.480 1011.830 ;
        RECT 899.860 1011.510 900.120 1011.830 ;
        RECT 899.920 1000.570 900.060 1011.510 ;
        RECT 899.920 1000.430 901.440 1000.570 ;
        RECT 901.300 999.330 901.440 1000.430 ;
        RECT 902.970 999.330 903.250 1000.000 ;
        RECT 901.300 999.190 903.250 999.330 ;
        RECT 902.970 996.000 903.250 999.190 ;
      LAYER via2 ;
        RECT 16.650 1465.600 16.930 1465.880 ;
      LAYER met3 ;
        RECT -4.800 1465.890 2.400 1466.340 ;
        RECT 16.625 1465.890 16.955 1465.905 ;
        RECT -4.800 1465.590 16.955 1465.890 ;
        RECT -4.800 1465.140 2.400 1465.590 ;
        RECT 16.625 1465.575 16.955 1465.590 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1200.780 15.570 1200.840 ;
        RECT 769.190 1200.780 769.510 1200.840 ;
        RECT 15.250 1200.640 769.510 1200.780 ;
        RECT 15.250 1200.580 15.570 1200.640 ;
        RECT 769.190 1200.580 769.510 1200.640 ;
        RECT 769.190 1012.080 769.510 1012.140 ;
        RECT 924.670 1012.080 924.990 1012.140 ;
        RECT 769.190 1011.940 924.990 1012.080 ;
        RECT 769.190 1011.880 769.510 1011.940 ;
        RECT 924.670 1011.880 924.990 1011.940 ;
      LAYER via ;
        RECT 15.280 1200.580 15.540 1200.840 ;
        RECT 769.220 1200.580 769.480 1200.840 ;
        RECT 769.220 1011.880 769.480 1012.140 ;
        RECT 924.700 1011.880 924.960 1012.140 ;
      LAYER met2 ;
        RECT 15.270 1205.115 15.550 1205.485 ;
        RECT 15.340 1200.870 15.480 1205.115 ;
        RECT 15.280 1200.550 15.540 1200.870 ;
        RECT 769.220 1200.550 769.480 1200.870 ;
        RECT 769.280 1012.170 769.420 1200.550 ;
        RECT 769.220 1011.850 769.480 1012.170 ;
        RECT 924.700 1011.850 924.960 1012.170 ;
        RECT 924.760 999.330 924.900 1011.850 ;
        RECT 925.050 999.330 925.330 1000.000 ;
        RECT 924.760 999.190 925.330 999.330 ;
        RECT 925.050 996.000 925.330 999.190 ;
      LAYER via2 ;
        RECT 15.270 1205.160 15.550 1205.440 ;
      LAYER met3 ;
        RECT -4.800 1205.450 2.400 1205.900 ;
        RECT 15.245 1205.450 15.575 1205.465 ;
        RECT -4.800 1205.150 15.575 1205.450 ;
        RECT -4.800 1204.700 2.400 1205.150 ;
        RECT 15.245 1205.135 15.575 1205.150 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.250 1004.940 15.570 1005.000 ;
        RECT 945.830 1004.940 946.150 1005.000 ;
        RECT 15.250 1004.800 946.150 1004.940 ;
        RECT 15.250 1004.740 15.570 1004.800 ;
        RECT 945.830 1004.740 946.150 1004.800 ;
      LAYER via ;
        RECT 15.280 1004.740 15.540 1005.000 ;
        RECT 945.860 1004.740 946.120 1005.000 ;
      LAYER met2 ;
        RECT 15.280 1004.710 15.540 1005.030 ;
        RECT 945.860 1004.710 946.120 1005.030 ;
        RECT 15.340 944.365 15.480 1004.710 ;
        RECT 945.920 999.330 946.060 1004.710 ;
        RECT 947.590 999.330 947.870 1000.000 ;
        RECT 945.920 999.190 947.870 999.330 ;
        RECT 947.590 996.000 947.870 999.190 ;
        RECT 15.270 943.995 15.550 944.365 ;
      LAYER via2 ;
        RECT 15.270 944.040 15.550 944.320 ;
      LAYER met3 ;
        RECT -4.800 944.330 2.400 944.780 ;
        RECT 15.245 944.330 15.575 944.345 ;
        RECT -4.800 944.030 15.575 944.330 ;
        RECT -4.800 943.580 2.400 944.030 ;
        RECT 15.245 944.015 15.575 944.030 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 1004.600 16.490 1004.660 ;
        RECT 967.910 1004.600 968.230 1004.660 ;
        RECT 16.170 1004.460 968.230 1004.600 ;
        RECT 16.170 1004.400 16.490 1004.460 ;
        RECT 967.910 1004.400 968.230 1004.460 ;
      LAYER via ;
        RECT 16.200 1004.400 16.460 1004.660 ;
        RECT 967.940 1004.400 968.200 1004.660 ;
      LAYER met2 ;
        RECT 16.200 1004.370 16.460 1004.690 ;
        RECT 967.940 1004.370 968.200 1004.690 ;
        RECT 16.260 683.925 16.400 1004.370 ;
        RECT 968.000 999.330 968.140 1004.370 ;
        RECT 969.670 999.330 969.950 1000.000 ;
        RECT 968.000 999.190 969.950 999.330 ;
        RECT 969.670 996.000 969.950 999.190 ;
        RECT 16.190 683.555 16.470 683.925 ;
      LAYER via2 ;
        RECT 16.190 683.600 16.470 683.880 ;
      LAYER met3 ;
        RECT -4.800 683.890 2.400 684.340 ;
        RECT 16.165 683.890 16.495 683.905 ;
        RECT -4.800 683.590 16.495 683.890 ;
        RECT -4.800 683.140 2.400 683.590 ;
        RECT 16.165 683.575 16.495 683.590 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 19.850 1003.580 20.170 1003.640 ;
        RECT 990.910 1003.580 991.230 1003.640 ;
        RECT 19.850 1003.440 991.230 1003.580 ;
        RECT 19.850 1003.380 20.170 1003.440 ;
        RECT 990.910 1003.380 991.230 1003.440 ;
      LAYER via ;
        RECT 19.880 1003.380 20.140 1003.640 ;
        RECT 990.940 1003.380 991.200 1003.640 ;
      LAYER met2 ;
        RECT 19.880 1003.350 20.140 1003.670 ;
        RECT 990.940 1003.350 991.200 1003.670 ;
        RECT 19.940 423.485 20.080 1003.350 ;
        RECT 991.000 999.330 991.140 1003.350 ;
        RECT 992.210 999.330 992.490 1000.000 ;
        RECT 991.000 999.190 992.490 999.330 ;
        RECT 992.210 996.000 992.490 999.190 ;
        RECT 19.870 423.115 20.150 423.485 ;
      LAYER via2 ;
        RECT 19.870 423.160 20.150 423.440 ;
      LAYER met3 ;
        RECT -4.800 423.450 2.400 423.900 ;
        RECT 19.845 423.450 20.175 423.465 ;
        RECT -4.800 423.150 20.175 423.450 ;
        RECT -4.800 422.700 2.400 423.150 ;
        RECT 19.845 423.135 20.175 423.150 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.470 1003.240 18.790 1003.300 ;
        RECT 1014.830 1003.240 1015.150 1003.300 ;
        RECT 18.470 1003.100 1015.150 1003.240 ;
        RECT 18.470 1003.040 18.790 1003.100 ;
        RECT 1014.830 1003.040 1015.150 1003.100 ;
      LAYER via ;
        RECT 18.500 1003.040 18.760 1003.300 ;
        RECT 1014.860 1003.040 1015.120 1003.300 ;
      LAYER met2 ;
        RECT 18.500 1003.010 18.760 1003.330 ;
        RECT 1014.860 1003.010 1015.120 1003.330 ;
        RECT 18.560 227.645 18.700 1003.010 ;
        RECT 1014.290 999.330 1014.570 1000.000 ;
        RECT 1014.920 999.330 1015.060 1003.010 ;
        RECT 1014.290 999.190 1015.060 999.330 ;
        RECT 1014.290 996.000 1014.570 999.190 ;
        RECT 18.490 227.275 18.770 227.645 ;
      LAYER via2 ;
        RECT 18.490 227.320 18.770 227.600 ;
      LAYER met3 ;
        RECT -4.800 227.610 2.400 228.060 ;
        RECT 18.465 227.610 18.795 227.625 ;
        RECT -4.800 227.310 18.795 227.610 ;
        RECT -4.800 226.860 2.400 227.310 ;
        RECT 18.465 227.295 18.795 227.310 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 23.990 1002.560 24.310 1002.620 ;
        RECT 1035.070 1002.560 1035.390 1002.620 ;
        RECT 23.990 1002.420 1035.390 1002.560 ;
        RECT 23.990 1002.360 24.310 1002.420 ;
        RECT 1035.070 1002.360 1035.390 1002.420 ;
        RECT 13.870 32.540 14.190 32.600 ;
        RECT 23.990 32.540 24.310 32.600 ;
        RECT 13.870 32.400 24.310 32.540 ;
        RECT 13.870 32.340 14.190 32.400 ;
        RECT 23.990 32.340 24.310 32.400 ;
      LAYER via ;
        RECT 24.020 1002.360 24.280 1002.620 ;
        RECT 1035.100 1002.360 1035.360 1002.620 ;
        RECT 13.900 32.340 14.160 32.600 ;
        RECT 24.020 32.340 24.280 32.600 ;
      LAYER met2 ;
        RECT 24.020 1002.330 24.280 1002.650 ;
        RECT 1035.100 1002.330 1035.360 1002.650 ;
        RECT 24.080 32.630 24.220 1002.330 ;
        RECT 1035.160 999.330 1035.300 1002.330 ;
        RECT 1036.830 999.330 1037.110 1000.000 ;
        RECT 1035.160 999.190 1037.110 999.330 ;
        RECT 1036.830 996.000 1037.110 999.190 ;
        RECT 13.900 32.485 14.160 32.630 ;
        RECT 13.890 32.115 14.170 32.485 ;
        RECT 24.020 32.310 24.280 32.630 ;
      LAYER via2 ;
        RECT 13.890 32.160 14.170 32.440 ;
      LAYER met3 ;
        RECT -4.800 32.450 2.400 32.900 ;
        RECT 13.865 32.450 14.195 32.465 ;
        RECT -4.800 32.150 14.195 32.450 ;
        RECT -4.800 31.700 2.400 32.150 ;
        RECT 13.865 32.135 14.195 32.150 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 279.290 1010.040 279.610 1010.100 ;
        RECT 1101.770 1010.040 1102.090 1010.100 ;
        RECT 279.290 1009.900 1102.090 1010.040 ;
        RECT 279.290 1009.840 279.610 1009.900 ;
        RECT 1101.770 1009.840 1102.090 1009.900 ;
        RECT 1101.770 765.920 1102.090 765.980 ;
        RECT 2898.990 765.920 2899.310 765.980 ;
        RECT 1101.770 765.780 2899.310 765.920 ;
        RECT 1101.770 765.720 1102.090 765.780 ;
        RECT 2898.990 765.720 2899.310 765.780 ;
      LAYER via ;
        RECT 279.320 1009.840 279.580 1010.100 ;
        RECT 1101.800 1009.840 1102.060 1010.100 ;
        RECT 1101.800 765.720 1102.060 765.980 ;
        RECT 2899.020 765.720 2899.280 765.980 ;
      LAYER met2 ;
        RECT 279.320 1009.810 279.580 1010.130 ;
        RECT 1101.800 1009.810 1102.060 1010.130 ;
        RECT 277.830 999.330 278.110 1000.000 ;
        RECT 279.380 999.330 279.520 1009.810 ;
        RECT 277.830 999.190 279.520 999.330 ;
        RECT 277.830 996.000 278.110 999.190 ;
        RECT 1101.860 766.010 1102.000 1009.810 ;
        RECT 1101.800 765.690 1102.060 766.010 ;
        RECT 2899.020 765.690 2899.280 766.010 ;
        RECT 2899.080 763.485 2899.220 765.690 ;
        RECT 2899.010 763.115 2899.290 763.485 ;
      LAYER via2 ;
        RECT 2899.010 763.160 2899.290 763.440 ;
      LAYER met3 ;
        RECT 2898.985 763.450 2899.315 763.465 ;
        RECT 2917.600 763.450 2924.800 763.900 ;
        RECT 2898.985 763.150 2924.800 763.450 ;
        RECT 2898.985 763.135 2899.315 763.150 ;
        RECT 2917.600 762.700 2924.800 763.150 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.830 1011.060 302.150 1011.120 ;
        RECT 1103.150 1011.060 1103.470 1011.120 ;
        RECT 301.830 1010.920 1103.470 1011.060 ;
        RECT 301.830 1010.860 302.150 1010.920 ;
        RECT 1103.150 1010.860 1103.470 1010.920 ;
        RECT 1103.150 965.840 1103.470 965.900 ;
        RECT 2900.830 965.840 2901.150 965.900 ;
        RECT 1103.150 965.700 2901.150 965.840 ;
        RECT 1103.150 965.640 1103.470 965.700 ;
        RECT 2900.830 965.640 2901.150 965.700 ;
      LAYER via ;
        RECT 301.860 1010.860 302.120 1011.120 ;
        RECT 1103.180 1010.860 1103.440 1011.120 ;
        RECT 1103.180 965.640 1103.440 965.900 ;
        RECT 2900.860 965.640 2901.120 965.900 ;
      LAYER met2 ;
        RECT 301.860 1010.830 302.120 1011.150 ;
        RECT 1103.180 1010.830 1103.440 1011.150 ;
        RECT 300.370 999.330 300.650 1000.000 ;
        RECT 301.920 999.330 302.060 1010.830 ;
        RECT 300.370 999.190 302.060 999.330 ;
        RECT 300.370 996.000 300.650 999.190 ;
        RECT 1103.240 965.930 1103.380 1010.830 ;
        RECT 1103.180 965.610 1103.440 965.930 ;
        RECT 2900.860 965.610 2901.120 965.930 ;
        RECT 2900.920 962.725 2901.060 965.610 ;
        RECT 2900.850 962.355 2901.130 962.725 ;
      LAYER via2 ;
        RECT 2900.850 962.400 2901.130 962.680 ;
      LAYER met3 ;
        RECT 2900.825 962.690 2901.155 962.705 ;
        RECT 2917.600 962.690 2924.800 963.140 ;
        RECT 2900.825 962.390 2924.800 962.690 ;
        RECT 2900.825 962.375 2901.155 962.390 ;
        RECT 2917.600 961.940 2924.800 962.390 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.470 1159.300 317.790 1159.360 ;
        RECT 2900.830 1159.300 2901.150 1159.360 ;
        RECT 317.470 1159.160 2901.150 1159.300 ;
        RECT 317.470 1159.100 317.790 1159.160 ;
        RECT 2900.830 1159.100 2901.150 1159.160 ;
      LAYER via ;
        RECT 317.500 1159.100 317.760 1159.360 ;
        RECT 2900.860 1159.100 2901.120 1159.360 ;
      LAYER met2 ;
        RECT 2900.850 1161.595 2901.130 1161.965 ;
        RECT 2900.920 1159.390 2901.060 1161.595 ;
        RECT 317.500 1159.070 317.760 1159.390 ;
        RECT 2900.860 1159.070 2901.120 1159.390 ;
        RECT 317.560 1048.870 317.700 1159.070 ;
        RECT 317.560 1048.730 320.920 1048.870 ;
        RECT 320.780 999.330 320.920 1048.730 ;
        RECT 322.450 999.330 322.730 1000.000 ;
        RECT 320.780 999.190 322.730 999.330 ;
        RECT 322.450 996.000 322.730 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1161.640 2901.130 1161.920 ;
      LAYER met3 ;
        RECT 2900.825 1161.930 2901.155 1161.945 ;
        RECT 2917.600 1161.930 2924.800 1162.380 ;
        RECT 2900.825 1161.630 2924.800 1161.930 ;
        RECT 2900.825 1161.615 2901.155 1161.630 ;
        RECT 2917.600 1161.180 2924.800 1161.630 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 1359.560 345.390 1359.620 ;
        RECT 2898.990 1359.560 2899.310 1359.620 ;
        RECT 345.070 1359.420 2899.310 1359.560 ;
        RECT 345.070 1359.360 345.390 1359.420 ;
        RECT 2898.990 1359.360 2899.310 1359.420 ;
      LAYER via ;
        RECT 345.100 1359.360 345.360 1359.620 ;
        RECT 2899.020 1359.360 2899.280 1359.620 ;
      LAYER met2 ;
        RECT 2899.010 1360.835 2899.290 1361.205 ;
        RECT 2899.080 1359.650 2899.220 1360.835 ;
        RECT 345.100 1359.330 345.360 1359.650 ;
        RECT 2899.020 1359.330 2899.280 1359.650 ;
        RECT 345.160 1048.870 345.300 1359.330 ;
        RECT 345.160 1048.730 345.760 1048.870 ;
        RECT 344.990 999.330 345.270 1000.000 ;
        RECT 345.620 999.330 345.760 1048.730 ;
        RECT 344.990 999.190 345.760 999.330 ;
        RECT 344.990 996.000 345.270 999.190 ;
      LAYER via2 ;
        RECT 2899.010 1360.880 2899.290 1361.160 ;
      LAYER met3 ;
        RECT 2898.985 1361.170 2899.315 1361.185 ;
        RECT 2917.600 1361.170 2924.800 1361.620 ;
        RECT 2898.985 1360.870 2924.800 1361.170 ;
        RECT 2898.985 1360.855 2899.315 1360.870 ;
        RECT 2917.600 1360.420 2924.800 1360.870 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 1621.700 366.090 1621.760 ;
        RECT 2900.830 1621.700 2901.150 1621.760 ;
        RECT 365.770 1621.560 2901.150 1621.700 ;
        RECT 365.770 1621.500 366.090 1621.560 ;
        RECT 2900.830 1621.500 2901.150 1621.560 ;
      LAYER via ;
        RECT 365.800 1621.500 366.060 1621.760 ;
        RECT 2900.860 1621.500 2901.120 1621.760 ;
      LAYER met2 ;
        RECT 2900.850 1626.035 2901.130 1626.405 ;
        RECT 2900.920 1621.790 2901.060 1626.035 ;
        RECT 365.800 1621.470 366.060 1621.790 ;
        RECT 2900.860 1621.470 2901.120 1621.790 ;
        RECT 365.860 999.330 366.000 1621.470 ;
        RECT 367.070 999.330 367.350 1000.000 ;
        RECT 365.860 999.190 367.350 999.330 ;
        RECT 367.070 996.000 367.350 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1626.080 2901.130 1626.360 ;
      LAYER met3 ;
        RECT 2900.825 1626.370 2901.155 1626.385 ;
        RECT 2917.600 1626.370 2924.800 1626.820 ;
        RECT 2900.825 1626.070 2924.800 1626.370 ;
        RECT 2900.825 1626.055 2901.155 1626.070 ;
        RECT 2917.600 1625.620 2924.800 1626.070 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.470 1890.980 386.790 1891.040 ;
        RECT 2900.830 1890.980 2901.150 1891.040 ;
        RECT 386.470 1890.840 2901.150 1890.980 ;
        RECT 386.470 1890.780 386.790 1890.840 ;
        RECT 2900.830 1890.780 2901.150 1890.840 ;
      LAYER via ;
        RECT 386.500 1890.780 386.760 1891.040 ;
        RECT 2900.860 1890.780 2901.120 1891.040 ;
      LAYER met2 ;
        RECT 2900.850 1891.915 2901.130 1892.285 ;
        RECT 2900.920 1891.070 2901.060 1891.915 ;
        RECT 386.500 1890.750 386.760 1891.070 ;
        RECT 2900.860 1890.750 2901.120 1891.070 ;
        RECT 386.560 1048.870 386.700 1890.750 ;
        RECT 386.560 1048.730 388.080 1048.870 ;
        RECT 387.940 999.330 388.080 1048.730 ;
        RECT 389.610 999.330 389.890 1000.000 ;
        RECT 387.940 999.190 389.890 999.330 ;
        RECT 389.610 996.000 389.890 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1891.960 2901.130 1892.240 ;
      LAYER met3 ;
        RECT 2900.825 1892.250 2901.155 1892.265 ;
        RECT 2917.600 1892.250 2924.800 1892.700 ;
        RECT 2900.825 1891.950 2924.800 1892.250 ;
        RECT 2900.825 1891.935 2901.155 1891.950 ;
        RECT 2917.600 1891.500 2924.800 1891.950 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 2153.120 407.490 2153.180 ;
        RECT 2900.830 2153.120 2901.150 2153.180 ;
        RECT 407.170 2152.980 2901.150 2153.120 ;
        RECT 407.170 2152.920 407.490 2152.980 ;
        RECT 2900.830 2152.920 2901.150 2152.980 ;
      LAYER via ;
        RECT 407.200 2152.920 407.460 2153.180 ;
        RECT 2900.860 2152.920 2901.120 2153.180 ;
      LAYER met2 ;
        RECT 2900.850 2157.795 2901.130 2158.165 ;
        RECT 2900.920 2153.210 2901.060 2157.795 ;
        RECT 407.200 2152.890 407.460 2153.210 ;
        RECT 2900.860 2152.890 2901.120 2153.210 ;
        RECT 407.260 1048.870 407.400 2152.890 ;
        RECT 407.260 1048.730 410.160 1048.870 ;
        RECT 410.020 999.330 410.160 1048.730 ;
        RECT 411.690 999.330 411.970 1000.000 ;
        RECT 410.020 999.190 411.970 999.330 ;
        RECT 411.690 996.000 411.970 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2157.840 2901.130 2158.120 ;
      LAYER met3 ;
        RECT 2900.825 2158.130 2901.155 2158.145 ;
        RECT 2917.600 2158.130 2924.800 2158.580 ;
        RECT 2900.825 2157.830 2924.800 2158.130 ;
        RECT 2900.825 2157.815 2901.155 2157.830 ;
        RECT 2917.600 2157.380 2924.800 2157.830 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 220.410 997.260 220.730 997.520 ;
        RECT 220.500 992.360 220.640 997.260 ;
        RECT 2901.290 993.720 2901.610 993.780 ;
        RECT 289.730 993.580 2901.610 993.720 ;
        RECT 289.730 992.700 289.870 993.580 ;
        RECT 2901.290 993.520 2901.610 993.580 ;
        RECT 275.930 992.560 289.870 992.700 ;
        RECT 275.930 992.360 276.070 992.560 ;
        RECT 220.500 992.220 276.070 992.360 ;
      LAYER via ;
        RECT 220.440 997.260 220.700 997.520 ;
        RECT 2901.320 993.520 2901.580 993.780 ;
      LAYER met2 ;
        RECT 218.490 997.290 218.770 1000.000 ;
        RECT 220.440 997.290 220.700 997.550 ;
        RECT 218.490 997.230 220.700 997.290 ;
        RECT 218.490 997.150 220.640 997.230 ;
        RECT 218.490 996.000 218.770 997.150 ;
        RECT 2901.320 993.490 2901.580 993.810 ;
        RECT 2901.380 99.125 2901.520 993.490 ;
        RECT 2901.310 98.755 2901.590 99.125 ;
      LAYER via2 ;
        RECT 2901.310 98.800 2901.590 99.080 ;
      LAYER met3 ;
        RECT 2901.285 99.090 2901.615 99.105 ;
        RECT 2917.600 99.090 2924.800 99.540 ;
        RECT 2901.285 98.790 2924.800 99.090 ;
        RECT 2901.285 98.775 2901.615 98.790 ;
        RECT 2917.600 98.340 2924.800 98.790 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 2353.040 441.990 2353.100 ;
        RECT 2899.910 2353.040 2900.230 2353.100 ;
        RECT 441.670 2352.900 2900.230 2353.040 ;
        RECT 441.670 2352.840 441.990 2352.900 ;
        RECT 2899.910 2352.840 2900.230 2352.900 ;
      LAYER via ;
        RECT 441.700 2352.840 441.960 2353.100 ;
        RECT 2899.940 2352.840 2900.200 2353.100 ;
      LAYER met2 ;
        RECT 2899.930 2357.035 2900.210 2357.405 ;
        RECT 2900.000 2353.130 2900.140 2357.035 ;
        RECT 441.700 2352.810 441.960 2353.130 ;
        RECT 2899.940 2352.810 2900.200 2353.130 ;
        RECT 441.760 1048.870 441.900 2352.810 ;
        RECT 441.760 1048.730 442.360 1048.870 ;
        RECT 441.590 999.330 441.870 1000.000 ;
        RECT 442.220 999.330 442.360 1048.730 ;
        RECT 441.590 999.190 442.360 999.330 ;
        RECT 441.590 996.000 441.870 999.190 ;
      LAYER via2 ;
        RECT 2899.930 2357.080 2900.210 2357.360 ;
      LAYER met3 ;
        RECT 2899.905 2357.370 2900.235 2357.385 ;
        RECT 2917.600 2357.370 2924.800 2357.820 ;
        RECT 2899.905 2357.070 2924.800 2357.370 ;
        RECT 2899.905 2357.055 2900.235 2357.070 ;
        RECT 2917.600 2356.620 2924.800 2357.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 2622.320 462.690 2622.380 ;
        RECT 2900.830 2622.320 2901.150 2622.380 ;
        RECT 462.370 2622.180 2901.150 2622.320 ;
        RECT 462.370 2622.120 462.690 2622.180 ;
        RECT 2900.830 2622.120 2901.150 2622.180 ;
      LAYER via ;
        RECT 462.400 2622.120 462.660 2622.380 ;
        RECT 2900.860 2622.120 2901.120 2622.380 ;
      LAYER met2 ;
        RECT 462.400 2622.090 462.660 2622.410 ;
        RECT 2900.850 2622.235 2901.130 2622.605 ;
        RECT 2900.860 2622.090 2901.120 2622.235 ;
        RECT 462.460 999.330 462.600 2622.090 ;
        RECT 464.130 999.330 464.410 1000.000 ;
        RECT 462.460 999.190 464.410 999.330 ;
        RECT 464.130 996.000 464.410 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2622.280 2901.130 2622.560 ;
      LAYER met3 ;
        RECT 2900.825 2622.570 2901.155 2622.585 ;
        RECT 2917.600 2622.570 2924.800 2623.020 ;
        RECT 2900.825 2622.270 2924.800 2622.570 ;
        RECT 2900.825 2622.255 2901.155 2622.270 ;
        RECT 2917.600 2621.820 2924.800 2622.270 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 2884.460 483.390 2884.520 ;
        RECT 2900.830 2884.460 2901.150 2884.520 ;
        RECT 483.070 2884.320 2901.150 2884.460 ;
        RECT 483.070 2884.260 483.390 2884.320 ;
        RECT 2900.830 2884.260 2901.150 2884.320 ;
      LAYER via ;
        RECT 483.100 2884.260 483.360 2884.520 ;
        RECT 2900.860 2884.260 2901.120 2884.520 ;
      LAYER met2 ;
        RECT 2900.850 2888.115 2901.130 2888.485 ;
        RECT 2900.920 2884.550 2901.060 2888.115 ;
        RECT 483.100 2884.230 483.360 2884.550 ;
        RECT 2900.860 2884.230 2901.120 2884.550 ;
        RECT 483.160 1048.870 483.300 2884.230 ;
        RECT 483.160 1048.730 484.680 1048.870 ;
        RECT 484.540 999.330 484.680 1048.730 ;
        RECT 486.210 999.330 486.490 1000.000 ;
        RECT 484.540 999.190 486.490 999.330 ;
        RECT 486.210 996.000 486.490 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2888.160 2901.130 2888.440 ;
      LAYER met3 ;
        RECT 2900.825 2888.450 2901.155 2888.465 ;
        RECT 2917.600 2888.450 2924.800 2888.900 ;
        RECT 2900.825 2888.150 2924.800 2888.450 ;
        RECT 2900.825 2888.135 2901.155 2888.150 ;
        RECT 2917.600 2887.700 2924.800 2888.150 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 3153.400 504.090 3153.460 ;
        RECT 2900.830 3153.400 2901.150 3153.460 ;
        RECT 503.770 3153.260 2901.150 3153.400 ;
        RECT 503.770 3153.200 504.090 3153.260 ;
        RECT 2900.830 3153.200 2901.150 3153.260 ;
      LAYER via ;
        RECT 503.800 3153.200 504.060 3153.460 ;
        RECT 2900.860 3153.200 2901.120 3153.460 ;
      LAYER met2 ;
        RECT 2900.850 3153.995 2901.130 3154.365 ;
        RECT 2900.920 3153.490 2901.060 3153.995 ;
        RECT 503.800 3153.170 504.060 3153.490 ;
        RECT 2900.860 3153.170 2901.120 3153.490 ;
        RECT 503.860 1048.870 504.000 3153.170 ;
        RECT 503.860 1048.730 506.760 1048.870 ;
        RECT 506.620 999.330 506.760 1048.730 ;
        RECT 508.750 999.330 509.030 1000.000 ;
        RECT 506.620 999.190 509.030 999.330 ;
        RECT 508.750 996.000 509.030 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3154.040 2901.130 3154.320 ;
      LAYER met3 ;
        RECT 2900.825 3154.330 2901.155 3154.345 ;
        RECT 2917.600 3154.330 2924.800 3154.780 ;
        RECT 2900.825 3154.030 2924.800 3154.330 ;
        RECT 2900.825 3154.015 2901.155 3154.030 ;
        RECT 2917.600 3153.580 2924.800 3154.030 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 3415.880 524.790 3415.940 ;
        RECT 2900.830 3415.880 2901.150 3415.940 ;
        RECT 524.470 3415.740 2901.150 3415.880 ;
        RECT 524.470 3415.680 524.790 3415.740 ;
        RECT 2900.830 3415.680 2901.150 3415.740 ;
      LAYER via ;
        RECT 524.500 3415.680 524.760 3415.940 ;
        RECT 2900.860 3415.680 2901.120 3415.940 ;
      LAYER met2 ;
        RECT 2900.850 3419.195 2901.130 3419.565 ;
        RECT 2900.920 3415.970 2901.060 3419.195 ;
        RECT 524.500 3415.650 524.760 3415.970 ;
        RECT 2900.860 3415.650 2901.120 3415.970 ;
        RECT 524.560 1048.870 524.700 3415.650 ;
        RECT 524.560 1048.730 528.840 1048.870 ;
        RECT 528.700 999.330 528.840 1048.730 ;
        RECT 530.830 999.330 531.110 1000.000 ;
        RECT 528.700 999.190 531.110 999.330 ;
        RECT 530.830 996.000 531.110 999.190 ;
      LAYER via2 ;
        RECT 2900.850 3419.240 2901.130 3419.520 ;
      LAYER met3 ;
        RECT 2900.825 3419.530 2901.155 3419.545 ;
        RECT 2917.600 3419.530 2924.800 3419.980 ;
        RECT 2900.825 3419.230 2924.800 3419.530 ;
        RECT 2900.825 3419.215 2901.155 3419.230 ;
        RECT 2917.600 3418.780 2924.800 3419.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 3501.560 552.390 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 552.070 3501.420 2717.610 3501.560 ;
        RECT 552.070 3501.360 552.390 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
      LAYER via ;
        RECT 552.100 3501.360 552.360 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 552.100 3501.330 552.360 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 552.160 999.330 552.300 3501.330 ;
        RECT 553.370 999.330 553.650 1000.000 ;
        RECT 552.160 999.190 553.650 999.330 ;
        RECT 553.370 996.000 553.650 999.190 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 3501.900 573.090 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 572.770 3501.760 2392.850 3501.900 ;
        RECT 572.770 3501.700 573.090 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 572.800 3501.700 573.060 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 572.800 3501.670 573.060 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 572.860 1048.870 573.000 3501.670 ;
        RECT 572.860 1048.730 573.920 1048.870 ;
        RECT 573.780 999.330 573.920 1048.730 ;
        RECT 575.450 999.330 575.730 1000.000 ;
        RECT 573.780 999.190 575.730 999.330 ;
        RECT 575.450 996.000 575.730 999.190 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 3502.920 593.790 3502.980 ;
        RECT 2068.230 3502.920 2068.550 3502.980 ;
        RECT 593.470 3502.780 2068.550 3502.920 ;
        RECT 593.470 3502.720 593.790 3502.780 ;
        RECT 2068.230 3502.720 2068.550 3502.780 ;
      LAYER via ;
        RECT 593.500 3502.720 593.760 3502.980 ;
        RECT 2068.260 3502.720 2068.520 3502.980 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3503.010 2068.460 3517.600 ;
        RECT 593.500 3502.690 593.760 3503.010 ;
        RECT 2068.260 3502.690 2068.520 3503.010 ;
        RECT 593.560 1048.870 593.700 3502.690 ;
        RECT 593.560 1048.730 596.000 1048.870 ;
        RECT 595.860 999.330 596.000 1048.730 ;
        RECT 597.990 999.330 598.270 1000.000 ;
        RECT 595.860 999.190 598.270 999.330 ;
        RECT 597.990 996.000 598.270 999.190 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 3503.600 614.490 3503.660 ;
        RECT 1743.930 3503.600 1744.250 3503.660 ;
        RECT 614.170 3503.460 1744.250 3503.600 ;
        RECT 614.170 3503.400 614.490 3503.460 ;
        RECT 1743.930 3503.400 1744.250 3503.460 ;
      LAYER via ;
        RECT 614.200 3503.400 614.460 3503.660 ;
        RECT 1743.960 3503.400 1744.220 3503.660 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.690 1744.160 3517.600 ;
        RECT 614.200 3503.370 614.460 3503.690 ;
        RECT 1743.960 3503.370 1744.220 3503.690 ;
        RECT 614.260 1048.870 614.400 3503.370 ;
        RECT 614.260 1048.730 618.080 1048.870 ;
        RECT 617.940 999.330 618.080 1048.730 ;
        RECT 620.070 999.330 620.350 1000.000 ;
        RECT 617.940 999.190 620.350 999.330 ;
        RECT 620.070 996.000 620.350 999.190 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 3504.280 642.090 3504.340 ;
        RECT 1419.170 3504.280 1419.490 3504.340 ;
        RECT 641.770 3504.140 1419.490 3504.280 ;
        RECT 641.770 3504.080 642.090 3504.140 ;
        RECT 1419.170 3504.080 1419.490 3504.140 ;
      LAYER via ;
        RECT 641.800 3504.080 642.060 3504.340 ;
        RECT 1419.200 3504.080 1419.460 3504.340 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3504.370 1419.400 3517.600 ;
        RECT 641.800 3504.050 642.060 3504.370 ;
        RECT 1419.200 3504.050 1419.460 3504.370 ;
        RECT 641.860 999.330 642.000 3504.050 ;
        RECT 642.610 999.330 642.890 1000.000 ;
        RECT 641.860 999.190 642.890 999.330 ;
        RECT 642.610 996.000 642.890 999.190 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 242.490 998.140 242.810 998.200 ;
        RECT 281.130 998.140 281.450 998.200 ;
        RECT 242.490 998.000 281.450 998.140 ;
        RECT 242.490 997.940 242.810 998.000 ;
        RECT 281.130 997.940 281.450 998.000 ;
        RECT 281.130 997.260 281.450 997.520 ;
        RECT 281.220 997.120 281.360 997.260 ;
        RECT 281.220 996.980 281.820 997.120 ;
        RECT 281.680 995.420 281.820 996.980 ;
        RECT 281.680 995.280 303.670 995.420 ;
        RECT 303.530 994.400 303.670 995.280 ;
        RECT 2902.670 994.400 2902.990 994.460 ;
        RECT 303.530 994.260 2902.990 994.400 ;
        RECT 2902.670 994.200 2902.990 994.260 ;
      LAYER via ;
        RECT 242.520 997.940 242.780 998.200 ;
        RECT 281.160 997.940 281.420 998.200 ;
        RECT 281.160 997.260 281.420 997.520 ;
        RECT 2902.700 994.200 2902.960 994.460 ;
      LAYER met2 ;
        RECT 240.570 997.970 240.850 1000.000 ;
        RECT 242.520 997.970 242.780 998.230 ;
        RECT 240.570 997.910 242.780 997.970 ;
        RECT 281.160 997.910 281.420 998.230 ;
        RECT 240.570 997.830 242.720 997.910 ;
        RECT 240.570 996.000 240.850 997.830 ;
        RECT 281.220 997.550 281.360 997.910 ;
        RECT 281.160 997.230 281.420 997.550 ;
        RECT 2902.700 994.170 2902.960 994.490 ;
        RECT 2902.760 298.365 2902.900 994.170 ;
        RECT 2902.690 297.995 2902.970 298.365 ;
      LAYER via2 ;
        RECT 2902.690 298.040 2902.970 298.320 ;
      LAYER met3 ;
        RECT 2902.665 298.330 2902.995 298.345 ;
        RECT 2917.600 298.330 2924.800 298.780 ;
        RECT 2902.665 298.030 2924.800 298.330 ;
        RECT 2902.665 298.015 2902.995 298.030 ;
        RECT 2917.600 297.580 2924.800 298.030 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 3504.960 662.790 3505.020 ;
        RECT 1094.870 3504.960 1095.190 3505.020 ;
        RECT 662.470 3504.820 1095.190 3504.960 ;
        RECT 662.470 3504.760 662.790 3504.820 ;
        RECT 1094.870 3504.760 1095.190 3504.820 ;
      LAYER via ;
        RECT 662.500 3504.760 662.760 3505.020 ;
        RECT 1094.900 3504.760 1095.160 3505.020 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3505.050 1095.100 3517.600 ;
        RECT 662.500 3504.730 662.760 3505.050 ;
        RECT 1094.900 3504.730 1095.160 3505.050 ;
        RECT 662.560 1048.870 662.700 3504.730 ;
        RECT 662.560 1048.730 663.160 1048.870 ;
        RECT 663.020 999.330 663.160 1048.730 ;
        RECT 664.690 999.330 664.970 1000.000 ;
        RECT 663.020 999.190 664.970 999.330 ;
        RECT 664.690 996.000 664.970 999.190 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 3500.540 683.950 3500.600 ;
        RECT 770.570 3500.540 770.890 3500.600 ;
        RECT 683.630 3500.400 770.890 3500.540 ;
        RECT 683.630 3500.340 683.950 3500.400 ;
        RECT 770.570 3500.340 770.890 3500.400 ;
      LAYER via ;
        RECT 683.660 3500.340 683.920 3500.600 ;
        RECT 770.600 3500.340 770.860 3500.600 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3500.630 770.800 3517.600 ;
        RECT 683.660 3500.310 683.920 3500.630 ;
        RECT 770.600 3500.310 770.860 3500.630 ;
        RECT 683.720 1048.870 683.860 3500.310 ;
        RECT 683.720 1048.730 685.240 1048.870 ;
        RECT 685.100 999.330 685.240 1048.730 ;
        RECT 687.230 999.330 687.510 1000.000 ;
        RECT 685.100 999.190 687.510 999.330 ;
        RECT 687.230 996.000 687.510 999.190 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 445.810 3504.620 446.130 3504.680 ;
        RECT 686.390 3504.620 686.710 3504.680 ;
        RECT 445.810 3504.480 686.710 3504.620 ;
        RECT 445.810 3504.420 446.130 3504.480 ;
        RECT 686.390 3504.420 686.710 3504.480 ;
        RECT 686.390 1014.120 686.710 1014.180 ;
        RECT 707.550 1014.120 707.870 1014.180 ;
        RECT 686.390 1013.980 707.870 1014.120 ;
        RECT 686.390 1013.920 686.710 1013.980 ;
        RECT 707.550 1013.920 707.870 1013.980 ;
      LAYER via ;
        RECT 445.840 3504.420 446.100 3504.680 ;
        RECT 686.420 3504.420 686.680 3504.680 ;
        RECT 686.420 1013.920 686.680 1014.180 ;
        RECT 707.580 1013.920 707.840 1014.180 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3504.710 446.040 3517.600 ;
        RECT 445.840 3504.390 446.100 3504.710 ;
        RECT 686.420 3504.390 686.680 3504.710 ;
        RECT 686.480 1014.210 686.620 3504.390 ;
        RECT 686.420 1013.890 686.680 1014.210 ;
        RECT 707.580 1013.890 707.840 1014.210 ;
        RECT 707.640 999.330 707.780 1013.890 ;
        RECT 709.310 999.330 709.590 1000.000 ;
        RECT 707.640 999.190 709.590 999.330 ;
        RECT 709.310 996.000 709.590 999.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 121.510 3502.580 121.830 3502.640 ;
        RECT 731.470 3502.580 731.790 3502.640 ;
        RECT 121.510 3502.440 731.790 3502.580 ;
        RECT 121.510 3502.380 121.830 3502.440 ;
        RECT 731.470 3502.380 731.790 3502.440 ;
      LAYER via ;
        RECT 121.540 3502.380 121.800 3502.640 ;
        RECT 731.500 3502.380 731.760 3502.640 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3502.670 121.740 3517.600 ;
        RECT 121.540 3502.350 121.800 3502.670 ;
        RECT 731.500 3502.350 731.760 3502.670 ;
        RECT 731.560 999.330 731.700 3502.350 ;
        RECT 731.850 999.330 732.130 1000.000 ;
        RECT 731.560 999.190 732.130 999.330 ;
        RECT 731.850 996.000 732.130 999.190 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.630 3354.000 16.950 3354.060 ;
        RECT 752.170 3354.000 752.490 3354.060 ;
        RECT 16.630 3353.860 752.490 3354.000 ;
        RECT 16.630 3353.800 16.950 3353.860 ;
        RECT 752.170 3353.800 752.490 3353.860 ;
      LAYER via ;
        RECT 16.660 3353.800 16.920 3354.060 ;
        RECT 752.200 3353.800 752.460 3354.060 ;
      LAYER met2 ;
        RECT 16.650 3355.955 16.930 3356.325 ;
        RECT 16.720 3354.090 16.860 3355.955 ;
        RECT 16.660 3353.770 16.920 3354.090 ;
        RECT 752.200 3353.770 752.460 3354.090 ;
        RECT 752.260 999.330 752.400 3353.770 ;
        RECT 753.930 999.330 754.210 1000.000 ;
        RECT 752.260 999.190 754.210 999.330 ;
        RECT 753.930 996.000 754.210 999.190 ;
      LAYER via2 ;
        RECT 16.650 3356.000 16.930 3356.280 ;
      LAYER met3 ;
        RECT -4.800 3356.290 2.400 3356.740 ;
        RECT 16.625 3356.290 16.955 3356.305 ;
        RECT -4.800 3355.990 16.955 3356.290 ;
        RECT -4.800 3355.540 2.400 3355.990 ;
        RECT 16.625 3355.975 16.955 3355.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 3091.520 17.870 3091.580 ;
        RECT 772.870 3091.520 773.190 3091.580 ;
        RECT 17.550 3091.380 773.190 3091.520 ;
        RECT 17.550 3091.320 17.870 3091.380 ;
        RECT 772.870 3091.320 773.190 3091.380 ;
      LAYER via ;
        RECT 17.580 3091.320 17.840 3091.580 ;
        RECT 772.900 3091.320 773.160 3091.580 ;
      LAYER met2 ;
        RECT 17.570 3095.515 17.850 3095.885 ;
        RECT 17.640 3091.610 17.780 3095.515 ;
        RECT 17.580 3091.290 17.840 3091.610 ;
        RECT 772.900 3091.290 773.160 3091.610 ;
        RECT 772.960 1048.870 773.100 3091.290 ;
        RECT 772.960 1048.730 774.480 1048.870 ;
        RECT 774.340 999.330 774.480 1048.730 ;
        RECT 776.470 999.330 776.750 1000.000 ;
        RECT 774.340 999.190 776.750 999.330 ;
        RECT 776.470 996.000 776.750 999.190 ;
      LAYER via2 ;
        RECT 17.570 3095.560 17.850 3095.840 ;
      LAYER met3 ;
        RECT -4.800 3095.850 2.400 3096.300 ;
        RECT 17.545 3095.850 17.875 3095.865 ;
        RECT -4.800 3095.550 17.875 3095.850 ;
        RECT -4.800 3095.100 2.400 3095.550 ;
        RECT 17.545 3095.535 17.875 3095.550 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.170 2829.380 16.490 2829.440 ;
        RECT 793.570 2829.380 793.890 2829.440 ;
        RECT 16.170 2829.240 793.890 2829.380 ;
        RECT 16.170 2829.180 16.490 2829.240 ;
        RECT 793.570 2829.180 793.890 2829.240 ;
      LAYER via ;
        RECT 16.200 2829.180 16.460 2829.440 ;
        RECT 793.600 2829.180 793.860 2829.440 ;
      LAYER met2 ;
        RECT 16.190 2834.395 16.470 2834.765 ;
        RECT 16.260 2829.470 16.400 2834.395 ;
        RECT 16.200 2829.150 16.460 2829.470 ;
        RECT 793.600 2829.150 793.860 2829.470 ;
        RECT 793.660 1048.870 793.800 2829.150 ;
        RECT 793.660 1048.730 796.560 1048.870 ;
        RECT 796.420 999.330 796.560 1048.730 ;
        RECT 798.550 999.330 798.830 1000.000 ;
        RECT 796.420 999.190 798.830 999.330 ;
        RECT 798.550 996.000 798.830 999.190 ;
      LAYER via2 ;
        RECT 16.190 2834.440 16.470 2834.720 ;
      LAYER met3 ;
        RECT -4.800 2834.730 2.400 2835.180 ;
        RECT 16.165 2834.730 16.495 2834.745 ;
        RECT -4.800 2834.430 16.495 2834.730 ;
        RECT -4.800 2833.980 2.400 2834.430 ;
        RECT 16.165 2834.415 16.495 2834.430 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2574.040 17.870 2574.100 ;
        RECT 821.170 2574.040 821.490 2574.100 ;
        RECT 17.550 2573.900 821.490 2574.040 ;
        RECT 17.550 2573.840 17.870 2573.900 ;
        RECT 821.170 2573.840 821.490 2573.900 ;
      LAYER via ;
        RECT 17.580 2573.840 17.840 2574.100 ;
        RECT 821.200 2573.840 821.460 2574.100 ;
      LAYER met2 ;
        RECT 17.570 2573.955 17.850 2574.325 ;
        RECT 17.580 2573.810 17.840 2573.955 ;
        RECT 821.200 2573.810 821.460 2574.130 ;
        RECT 821.260 1048.870 821.400 2573.810 ;
        RECT 821.260 1048.730 821.860 1048.870 ;
        RECT 821.090 999.330 821.370 1000.000 ;
        RECT 821.720 999.330 821.860 1048.730 ;
        RECT 821.090 999.190 821.860 999.330 ;
        RECT 821.090 996.000 821.370 999.190 ;
      LAYER via2 ;
        RECT 17.570 2574.000 17.850 2574.280 ;
      LAYER met3 ;
        RECT -4.800 2574.290 2.400 2574.740 ;
        RECT 17.545 2574.290 17.875 2574.305 ;
        RECT -4.800 2573.990 17.875 2574.290 ;
        RECT -4.800 2573.540 2.400 2573.990 ;
        RECT 17.545 2573.975 17.875 2573.990 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 2311.900 17.870 2311.960 ;
        RECT 841.870 2311.900 842.190 2311.960 ;
        RECT 17.550 2311.760 842.190 2311.900 ;
        RECT 17.550 2311.700 17.870 2311.760 ;
        RECT 841.870 2311.700 842.190 2311.760 ;
      LAYER via ;
        RECT 17.580 2311.700 17.840 2311.960 ;
        RECT 841.900 2311.700 842.160 2311.960 ;
      LAYER met2 ;
        RECT 17.570 2312.835 17.850 2313.205 ;
        RECT 17.640 2311.990 17.780 2312.835 ;
        RECT 17.580 2311.670 17.840 2311.990 ;
        RECT 841.900 2311.670 842.160 2311.990 ;
        RECT 841.960 999.330 842.100 2311.670 ;
        RECT 843.170 999.330 843.450 1000.000 ;
        RECT 841.960 999.190 843.450 999.330 ;
        RECT 843.170 996.000 843.450 999.190 ;
      LAYER via2 ;
        RECT 17.570 2312.880 17.850 2313.160 ;
      LAYER met3 ;
        RECT -4.800 2313.170 2.400 2313.620 ;
        RECT 17.545 2313.170 17.875 2313.185 ;
        RECT -4.800 2312.870 17.875 2313.170 ;
        RECT -4.800 2312.420 2.400 2312.870 ;
        RECT 17.545 2312.855 17.875 2312.870 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.330 2049.420 14.650 2049.480 ;
        RECT 862.570 2049.420 862.890 2049.480 ;
        RECT 14.330 2049.280 862.890 2049.420 ;
        RECT 14.330 2049.220 14.650 2049.280 ;
        RECT 862.570 2049.220 862.890 2049.280 ;
      LAYER via ;
        RECT 14.360 2049.220 14.620 2049.480 ;
        RECT 862.600 2049.220 862.860 2049.480 ;
      LAYER met2 ;
        RECT 14.350 2052.395 14.630 2052.765 ;
        RECT 14.420 2049.510 14.560 2052.395 ;
        RECT 14.360 2049.190 14.620 2049.510 ;
        RECT 862.600 2049.190 862.860 2049.510 ;
        RECT 862.660 1048.870 862.800 2049.190 ;
        RECT 862.660 1048.730 863.720 1048.870 ;
        RECT 863.580 999.330 863.720 1048.730 ;
        RECT 865.710 999.330 865.990 1000.000 ;
        RECT 863.580 999.190 865.990 999.330 ;
        RECT 865.710 996.000 865.990 999.190 ;
      LAYER via2 ;
        RECT 14.350 2052.440 14.630 2052.720 ;
      LAYER met3 ;
        RECT -4.800 2052.730 2.400 2053.180 ;
        RECT 14.325 2052.730 14.655 2052.745 ;
        RECT -4.800 2052.430 14.655 2052.730 ;
        RECT -4.800 2051.980 2.400 2052.430 ;
        RECT 14.325 2052.415 14.655 2052.430 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 264.570 1009.360 264.890 1009.420 ;
        RECT 1100.390 1009.360 1100.710 1009.420 ;
        RECT 264.570 1009.220 1100.710 1009.360 ;
        RECT 264.570 1009.160 264.890 1009.220 ;
        RECT 1100.390 1009.160 1100.710 1009.220 ;
        RECT 1100.390 503.440 1100.710 503.500 ;
        RECT 2900.830 503.440 2901.150 503.500 ;
        RECT 1100.390 503.300 2901.150 503.440 ;
        RECT 1100.390 503.240 1100.710 503.300 ;
        RECT 2900.830 503.240 2901.150 503.300 ;
      LAYER via ;
        RECT 264.600 1009.160 264.860 1009.420 ;
        RECT 1100.420 1009.160 1100.680 1009.420 ;
        RECT 1100.420 503.240 1100.680 503.500 ;
        RECT 2900.860 503.240 2901.120 503.500 ;
      LAYER met2 ;
        RECT 264.600 1009.130 264.860 1009.450 ;
        RECT 1100.420 1009.130 1100.680 1009.450 ;
        RECT 263.110 999.330 263.390 1000.000 ;
        RECT 264.660 999.330 264.800 1009.130 ;
        RECT 263.110 999.190 264.800 999.330 ;
        RECT 263.110 996.000 263.390 999.190 ;
        RECT 1100.480 503.530 1100.620 1009.130 ;
        RECT 1100.420 503.210 1100.680 503.530 ;
        RECT 2900.860 503.210 2901.120 503.530 ;
        RECT 2900.920 497.605 2901.060 503.210 ;
        RECT 2900.850 497.235 2901.130 497.605 ;
      LAYER via2 ;
        RECT 2900.850 497.280 2901.130 497.560 ;
      LAYER met3 ;
        RECT 2900.825 497.570 2901.155 497.585 ;
        RECT 2917.600 497.570 2924.800 498.020 ;
        RECT 2900.825 497.270 2924.800 497.570 ;
        RECT 2900.825 497.255 2901.155 497.270 ;
        RECT 2917.600 496.820 2924.800 497.270 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1787.280 16.030 1787.340 ;
        RECT 883.270 1787.280 883.590 1787.340 ;
        RECT 15.710 1787.140 883.590 1787.280 ;
        RECT 15.710 1787.080 16.030 1787.140 ;
        RECT 883.270 1787.080 883.590 1787.140 ;
      LAYER via ;
        RECT 15.740 1787.080 16.000 1787.340 ;
        RECT 883.300 1787.080 883.560 1787.340 ;
      LAYER met2 ;
        RECT 15.730 1791.955 16.010 1792.325 ;
        RECT 15.800 1787.370 15.940 1791.955 ;
        RECT 15.740 1787.050 16.000 1787.370 ;
        RECT 883.300 1787.050 883.560 1787.370 ;
        RECT 883.360 1048.870 883.500 1787.050 ;
        RECT 883.360 1048.730 885.800 1048.870 ;
        RECT 885.660 999.330 885.800 1048.730 ;
        RECT 887.790 999.330 888.070 1000.000 ;
        RECT 885.660 999.190 888.070 999.330 ;
        RECT 887.790 996.000 888.070 999.190 ;
      LAYER via2 ;
        RECT 15.730 1792.000 16.010 1792.280 ;
      LAYER met3 ;
        RECT -4.800 1792.290 2.400 1792.740 ;
        RECT 15.705 1792.290 16.035 1792.305 ;
        RECT -4.800 1791.990 16.035 1792.290 ;
        RECT -4.800 1791.540 2.400 1791.990 ;
        RECT 15.705 1791.975 16.035 1791.990 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1525.140 17.870 1525.200 ;
        RECT 903.970 1525.140 904.290 1525.200 ;
        RECT 17.550 1525.000 904.290 1525.140 ;
        RECT 17.550 1524.940 17.870 1525.000 ;
        RECT 903.970 1524.940 904.290 1525.000 ;
      LAYER via ;
        RECT 17.580 1524.940 17.840 1525.200 ;
        RECT 904.000 1524.940 904.260 1525.200 ;
      LAYER met2 ;
        RECT 17.570 1530.835 17.850 1531.205 ;
        RECT 17.640 1525.230 17.780 1530.835 ;
        RECT 17.580 1524.910 17.840 1525.230 ;
        RECT 904.000 1524.910 904.260 1525.230 ;
        RECT 904.060 1048.870 904.200 1524.910 ;
        RECT 904.060 1048.730 908.800 1048.870 ;
        RECT 908.660 999.330 908.800 1048.730 ;
        RECT 910.330 999.330 910.610 1000.000 ;
        RECT 908.660 999.190 910.610 999.330 ;
        RECT 910.330 996.000 910.610 999.190 ;
      LAYER via2 ;
        RECT 17.570 1530.880 17.850 1531.160 ;
      LAYER met3 ;
        RECT -4.800 1531.170 2.400 1531.620 ;
        RECT 17.545 1531.170 17.875 1531.185 ;
        RECT -4.800 1530.870 17.875 1531.170 ;
        RECT -4.800 1530.420 2.400 1530.870 ;
        RECT 17.545 1530.855 17.875 1530.870 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 15.710 1269.800 16.030 1269.860 ;
        RECT 900.290 1269.800 900.610 1269.860 ;
        RECT 15.710 1269.660 900.610 1269.800 ;
        RECT 15.710 1269.600 16.030 1269.660 ;
        RECT 900.290 1269.600 900.610 1269.660 ;
        RECT 900.290 1011.740 900.610 1011.800 ;
        RECT 931.570 1011.740 931.890 1011.800 ;
        RECT 900.290 1011.600 931.890 1011.740 ;
        RECT 900.290 1011.540 900.610 1011.600 ;
        RECT 931.570 1011.540 931.890 1011.600 ;
      LAYER via ;
        RECT 15.740 1269.600 16.000 1269.860 ;
        RECT 900.320 1269.600 900.580 1269.860 ;
        RECT 900.320 1011.540 900.580 1011.800 ;
        RECT 931.600 1011.540 931.860 1011.800 ;
      LAYER met2 ;
        RECT 15.730 1270.395 16.010 1270.765 ;
        RECT 15.800 1269.890 15.940 1270.395 ;
        RECT 15.740 1269.570 16.000 1269.890 ;
        RECT 900.320 1269.570 900.580 1269.890 ;
        RECT 900.380 1011.830 900.520 1269.570 ;
        RECT 900.320 1011.510 900.580 1011.830 ;
        RECT 931.600 1011.510 931.860 1011.830 ;
        RECT 931.660 999.330 931.800 1011.510 ;
        RECT 932.870 999.330 933.150 1000.000 ;
        RECT 931.660 999.190 933.150 999.330 ;
        RECT 932.870 996.000 933.150 999.190 ;
      LAYER via2 ;
        RECT 15.730 1270.440 16.010 1270.720 ;
      LAYER met3 ;
        RECT -4.800 1270.730 2.400 1271.180 ;
        RECT 15.705 1270.730 16.035 1270.745 ;
        RECT -4.800 1270.430 16.035 1270.730 ;
        RECT -4.800 1269.980 2.400 1270.430 ;
        RECT 15.705 1270.415 16.035 1270.430 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 17.550 1009.020 17.870 1009.080 ;
        RECT 953.190 1009.020 953.510 1009.080 ;
        RECT 17.550 1008.880 953.510 1009.020 ;
        RECT 17.550 1008.820 17.870 1008.880 ;
        RECT 953.190 1008.820 953.510 1008.880 ;
      LAYER via ;
        RECT 17.580 1008.820 17.840 1009.080 ;
        RECT 953.220 1008.820 953.480 1009.080 ;
      LAYER met2 ;
        RECT 17.570 1009.275 17.850 1009.645 ;
        RECT 17.640 1009.110 17.780 1009.275 ;
        RECT 17.580 1008.790 17.840 1009.110 ;
        RECT 953.220 1008.790 953.480 1009.110 ;
        RECT 953.280 999.330 953.420 1008.790 ;
        RECT 954.950 999.330 955.230 1000.000 ;
        RECT 953.280 999.190 955.230 999.330 ;
        RECT 954.950 996.000 955.230 999.190 ;
      LAYER via2 ;
        RECT 17.570 1009.320 17.850 1009.600 ;
      LAYER met3 ;
        RECT -4.800 1009.610 2.400 1010.060 ;
        RECT 17.545 1009.610 17.875 1009.625 ;
        RECT -4.800 1009.310 17.875 1009.610 ;
        RECT -4.800 1008.860 2.400 1009.310 ;
        RECT 17.545 1009.295 17.875 1009.310 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 201.090 997.800 201.410 997.860 ;
        RECT 201.090 997.660 229.380 997.800 ;
        RECT 201.090 997.600 201.410 997.660 ;
        RECT 229.240 996.780 229.380 997.660 ;
        RECT 265.120 997.660 317.470 997.800 ;
        RECT 265.120 996.780 265.260 997.660 ;
        RECT 317.330 997.120 317.470 997.660 ;
        RECT 976.190 997.460 976.510 997.520 ;
        RECT 903.830 997.320 976.510 997.460 ;
        RECT 317.330 996.980 324.370 997.120 ;
        RECT 229.240 996.640 265.260 996.780 ;
        RECT 201.090 995.760 201.410 995.820 ;
        RECT 131.030 995.620 201.410 995.760 ;
        RECT 24.910 995.080 25.230 995.140 ;
        RECT 131.030 995.080 131.170 995.620 ;
        RECT 201.090 995.560 201.410 995.620 ;
        RECT 24.910 994.940 131.170 995.080 ;
        RECT 324.230 995.080 324.370 996.980 ;
        RECT 903.830 995.080 903.970 997.320 ;
        RECT 976.190 997.260 976.510 997.320 ;
        RECT 324.230 994.940 903.970 995.080 ;
        RECT 24.910 994.880 25.230 994.940 ;
        RECT 13.870 750.280 14.190 750.340 ;
        RECT 24.910 750.280 25.230 750.340 ;
        RECT 13.870 750.140 25.230 750.280 ;
        RECT 13.870 750.080 14.190 750.140 ;
        RECT 24.910 750.080 25.230 750.140 ;
      LAYER via ;
        RECT 201.120 997.600 201.380 997.860 ;
        RECT 24.940 994.880 25.200 995.140 ;
        RECT 201.120 995.560 201.380 995.820 ;
        RECT 976.220 997.260 976.480 997.520 ;
        RECT 13.900 750.080 14.160 750.340 ;
        RECT 24.940 750.080 25.200 750.340 ;
      LAYER met2 ;
        RECT 201.120 997.570 201.380 997.890 ;
        RECT 201.180 995.850 201.320 997.570 ;
        RECT 976.220 997.290 976.480 997.550 ;
        RECT 977.490 997.290 977.770 1000.000 ;
        RECT 976.220 997.230 977.770 997.290 ;
        RECT 976.280 997.150 977.770 997.230 ;
        RECT 977.490 996.000 977.770 997.150 ;
        RECT 201.120 995.530 201.380 995.850 ;
        RECT 24.940 994.850 25.200 995.170 ;
        RECT 25.000 750.370 25.140 994.850 ;
        RECT 13.900 750.050 14.160 750.370 ;
        RECT 24.940 750.050 25.200 750.370 ;
        RECT 13.960 749.205 14.100 750.050 ;
        RECT 13.890 748.835 14.170 749.205 ;
      LAYER via2 ;
        RECT 13.890 748.880 14.170 749.160 ;
      LAYER met3 ;
        RECT -4.800 749.170 2.400 749.620 ;
        RECT 13.865 749.170 14.195 749.185 ;
        RECT -4.800 748.870 14.195 749.170 ;
        RECT -4.800 748.420 2.400 748.870 ;
        RECT 13.865 748.855 14.195 748.870 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 20.310 1008.000 20.630 1008.060 ;
        RECT 998.270 1008.000 998.590 1008.060 ;
        RECT 20.310 1007.860 998.590 1008.000 ;
        RECT 20.310 1007.800 20.630 1007.860 ;
        RECT 998.270 1007.800 998.590 1007.860 ;
      LAYER via ;
        RECT 20.340 1007.800 20.600 1008.060 ;
        RECT 998.300 1007.800 998.560 1008.060 ;
      LAYER met2 ;
        RECT 20.340 1007.770 20.600 1008.090 ;
        RECT 998.300 1007.770 998.560 1008.090 ;
        RECT 20.400 488.085 20.540 1007.770 ;
        RECT 998.360 999.330 998.500 1007.770 ;
        RECT 999.570 999.330 999.850 1000.000 ;
        RECT 998.360 999.190 999.850 999.330 ;
        RECT 999.570 996.000 999.850 999.190 ;
        RECT 20.330 487.715 20.610 488.085 ;
      LAYER via2 ;
        RECT 20.330 487.760 20.610 488.040 ;
      LAYER met3 ;
        RECT -4.800 488.050 2.400 488.500 ;
        RECT 20.305 488.050 20.635 488.065 ;
        RECT -4.800 487.750 20.635 488.050 ;
        RECT -4.800 487.300 2.400 487.750 ;
        RECT 20.305 487.735 20.635 487.750 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 18.930 1007.660 19.250 1007.720 ;
        RECT 1021.270 1007.660 1021.590 1007.720 ;
        RECT 18.930 1007.520 1021.590 1007.660 ;
        RECT 18.930 1007.460 19.250 1007.520 ;
        RECT 1021.270 1007.460 1021.590 1007.520 ;
      LAYER via ;
        RECT 18.960 1007.460 19.220 1007.720 ;
        RECT 1021.300 1007.460 1021.560 1007.720 ;
      LAYER met2 ;
        RECT 18.960 1007.430 19.220 1007.750 ;
        RECT 1021.300 1007.430 1021.560 1007.750 ;
        RECT 19.020 292.925 19.160 1007.430 ;
        RECT 1021.360 999.330 1021.500 1007.430 ;
        RECT 1022.110 999.330 1022.390 1000.000 ;
        RECT 1021.360 999.190 1022.390 999.330 ;
        RECT 1022.110 996.000 1022.390 999.190 ;
        RECT 18.950 292.555 19.230 292.925 ;
      LAYER via2 ;
        RECT 18.950 292.600 19.230 292.880 ;
      LAYER met3 ;
        RECT -4.800 292.890 2.400 293.340 ;
        RECT 18.925 292.890 19.255 292.905 ;
        RECT -4.800 292.590 19.255 292.890 ;
        RECT -4.800 292.140 2.400 292.590 ;
        RECT 18.925 292.575 19.255 292.590 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.450 1002.220 24.770 1002.280 ;
        RECT 1042.430 1002.220 1042.750 1002.280 ;
        RECT 24.450 1002.080 1042.750 1002.220 ;
        RECT 24.450 1002.020 24.770 1002.080 ;
        RECT 1042.430 1002.020 1042.750 1002.080 ;
        RECT 14.330 101.900 14.650 101.960 ;
        RECT 24.450 101.900 24.770 101.960 ;
        RECT 14.330 101.760 24.770 101.900 ;
        RECT 14.330 101.700 14.650 101.760 ;
        RECT 24.450 101.700 24.770 101.760 ;
      LAYER via ;
        RECT 24.480 1002.020 24.740 1002.280 ;
        RECT 1042.460 1002.020 1042.720 1002.280 ;
        RECT 14.360 101.700 14.620 101.960 ;
        RECT 24.480 101.700 24.740 101.960 ;
      LAYER met2 ;
        RECT 24.480 1001.990 24.740 1002.310 ;
        RECT 1042.460 1001.990 1042.720 1002.310 ;
        RECT 24.540 101.990 24.680 1001.990 ;
        RECT 1042.520 999.330 1042.660 1001.990 ;
        RECT 1044.190 999.330 1044.470 1000.000 ;
        RECT 1042.520 999.190 1044.470 999.330 ;
        RECT 1044.190 996.000 1044.470 999.190 ;
        RECT 14.360 101.670 14.620 101.990 ;
        RECT 24.480 101.670 24.740 101.990 ;
        RECT 14.420 97.085 14.560 101.670 ;
        RECT 14.350 96.715 14.630 97.085 ;
      LAYER via2 ;
        RECT 14.350 96.760 14.630 97.040 ;
      LAYER met3 ;
        RECT -4.800 97.050 2.400 97.500 ;
        RECT 14.325 97.050 14.655 97.065 ;
        RECT -4.800 96.750 14.655 97.050 ;
        RECT -4.800 96.300 2.400 96.750 ;
        RECT 14.325 96.735 14.655 96.750 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 286.650 1010.380 286.970 1010.440 ;
        RECT 1101.310 1010.380 1101.630 1010.440 ;
        RECT 286.650 1010.240 1101.630 1010.380 ;
        RECT 286.650 1010.180 286.970 1010.240 ;
        RECT 1101.310 1010.180 1101.630 1010.240 ;
        RECT 1101.310 696.900 1101.630 696.960 ;
        RECT 2900.830 696.900 2901.150 696.960 ;
        RECT 1101.310 696.760 2901.150 696.900 ;
        RECT 1101.310 696.700 1101.630 696.760 ;
        RECT 2900.830 696.700 2901.150 696.760 ;
      LAYER via ;
        RECT 286.680 1010.180 286.940 1010.440 ;
        RECT 1101.340 1010.180 1101.600 1010.440 ;
        RECT 1101.340 696.700 1101.600 696.960 ;
        RECT 2900.860 696.700 2901.120 696.960 ;
      LAYER met2 ;
        RECT 286.680 1010.150 286.940 1010.470 ;
        RECT 1101.340 1010.150 1101.600 1010.470 ;
        RECT 285.190 999.330 285.470 1000.000 ;
        RECT 286.740 999.330 286.880 1010.150 ;
        RECT 285.190 999.190 286.880 999.330 ;
        RECT 285.190 996.000 285.470 999.190 ;
        RECT 1101.400 696.990 1101.540 1010.150 ;
        RECT 1101.340 696.670 1101.600 696.990 ;
        RECT 2900.860 696.845 2901.120 696.990 ;
        RECT 2900.850 696.475 2901.130 696.845 ;
      LAYER via2 ;
        RECT 2900.850 696.520 2901.130 696.800 ;
      LAYER met3 ;
        RECT 2900.825 696.810 2901.155 696.825 ;
        RECT 2917.600 696.810 2924.800 697.260 ;
        RECT 2900.825 696.510 2924.800 696.810 ;
        RECT 2900.825 696.495 2901.155 696.510 ;
        RECT 2917.600 696.060 2924.800 696.510 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 309.650 1011.400 309.970 1011.460 ;
        RECT 1102.690 1011.400 1103.010 1011.460 ;
        RECT 309.650 1011.260 1103.010 1011.400 ;
        RECT 309.650 1011.200 309.970 1011.260 ;
        RECT 1102.690 1011.200 1103.010 1011.260 ;
        RECT 1102.690 896.820 1103.010 896.880 ;
        RECT 2898.990 896.820 2899.310 896.880 ;
        RECT 1102.690 896.680 2899.310 896.820 ;
        RECT 1102.690 896.620 1103.010 896.680 ;
        RECT 2898.990 896.620 2899.310 896.680 ;
      LAYER via ;
        RECT 309.680 1011.200 309.940 1011.460 ;
        RECT 1102.720 1011.200 1102.980 1011.460 ;
        RECT 1102.720 896.620 1102.980 896.880 ;
        RECT 2899.020 896.620 2899.280 896.880 ;
      LAYER met2 ;
        RECT 309.680 1011.170 309.940 1011.490 ;
        RECT 1102.720 1011.170 1102.980 1011.490 ;
        RECT 307.730 999.330 308.010 1000.000 ;
        RECT 309.740 999.330 309.880 1011.170 ;
        RECT 307.730 999.190 309.880 999.330 ;
        RECT 307.730 996.000 308.010 999.190 ;
        RECT 1102.780 896.910 1102.920 1011.170 ;
        RECT 1102.720 896.590 1102.980 896.910 ;
        RECT 2899.020 896.590 2899.280 896.910 ;
        RECT 2899.080 896.085 2899.220 896.590 ;
        RECT 2899.010 895.715 2899.290 896.085 ;
      LAYER via2 ;
        RECT 2899.010 895.760 2899.290 896.040 ;
      LAYER met3 ;
        RECT 2898.985 896.050 2899.315 896.065 ;
        RECT 2917.600 896.050 2924.800 896.500 ;
        RECT 2898.985 895.750 2924.800 896.050 ;
        RECT 2898.985 895.735 2899.315 895.750 ;
        RECT 2917.600 895.300 2924.800 895.750 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 1090.280 324.690 1090.340 ;
        RECT 2900.830 1090.280 2901.150 1090.340 ;
        RECT 324.370 1090.140 2901.150 1090.280 ;
        RECT 324.370 1090.080 324.690 1090.140 ;
        RECT 2900.830 1090.080 2901.150 1090.140 ;
      LAYER via ;
        RECT 324.400 1090.080 324.660 1090.340 ;
        RECT 2900.860 1090.080 2901.120 1090.340 ;
      LAYER met2 ;
        RECT 2900.850 1094.955 2901.130 1095.325 ;
        RECT 2900.920 1090.370 2901.060 1094.955 ;
        RECT 324.400 1090.050 324.660 1090.370 ;
        RECT 2900.860 1090.050 2901.120 1090.370 ;
        RECT 324.460 1048.870 324.600 1090.050 ;
        RECT 324.460 1048.730 328.280 1048.870 ;
        RECT 328.140 999.330 328.280 1048.730 ;
        RECT 329.810 999.330 330.090 1000.000 ;
        RECT 328.140 999.190 330.090 999.330 ;
        RECT 329.810 996.000 330.090 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1095.000 2901.130 1095.280 ;
      LAYER met3 ;
        RECT 2900.825 1095.290 2901.155 1095.305 ;
        RECT 2917.600 1095.290 2924.800 1095.740 ;
        RECT 2900.825 1094.990 2924.800 1095.290 ;
        RECT 2900.825 1094.975 2901.155 1094.990 ;
        RECT 2917.600 1094.540 2924.800 1094.990 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.970 1290.540 352.290 1290.600 ;
        RECT 2900.830 1290.540 2901.150 1290.600 ;
        RECT 351.970 1290.400 2901.150 1290.540 ;
        RECT 351.970 1290.340 352.290 1290.400 ;
        RECT 2900.830 1290.340 2901.150 1290.400 ;
      LAYER via ;
        RECT 352.000 1290.340 352.260 1290.600 ;
        RECT 2900.860 1290.340 2901.120 1290.600 ;
      LAYER met2 ;
        RECT 2900.850 1294.195 2901.130 1294.565 ;
        RECT 2900.920 1290.630 2901.060 1294.195 ;
        RECT 352.000 1290.310 352.260 1290.630 ;
        RECT 2900.860 1290.310 2901.120 1290.630 ;
        RECT 352.060 999.330 352.200 1290.310 ;
        RECT 352.350 999.330 352.630 1000.000 ;
        RECT 352.060 999.190 352.630 999.330 ;
        RECT 352.350 996.000 352.630 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1294.240 2901.130 1294.520 ;
      LAYER met3 ;
        RECT 2900.825 1294.530 2901.155 1294.545 ;
        RECT 2917.600 1294.530 2924.800 1294.980 ;
        RECT 2900.825 1294.230 2924.800 1294.530 ;
        RECT 2900.825 1294.215 2901.155 1294.230 ;
        RECT 2917.600 1293.780 2924.800 1294.230 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 1559.480 372.990 1559.540 ;
        RECT 2900.830 1559.480 2901.150 1559.540 ;
        RECT 372.670 1559.340 2901.150 1559.480 ;
        RECT 372.670 1559.280 372.990 1559.340 ;
        RECT 2900.830 1559.280 2901.150 1559.340 ;
      LAYER via ;
        RECT 372.700 1559.280 372.960 1559.540 ;
        RECT 2900.860 1559.280 2901.120 1559.540 ;
      LAYER met2 ;
        RECT 2900.850 1560.075 2901.130 1560.445 ;
        RECT 2900.920 1559.570 2901.060 1560.075 ;
        RECT 372.700 1559.250 372.960 1559.570 ;
        RECT 2900.860 1559.250 2901.120 1559.570 ;
        RECT 372.760 999.330 372.900 1559.250 ;
        RECT 374.430 999.330 374.710 1000.000 ;
        RECT 372.760 999.190 374.710 999.330 ;
        RECT 374.430 996.000 374.710 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1560.120 2901.130 1560.400 ;
      LAYER met3 ;
        RECT 2900.825 1560.410 2901.155 1560.425 ;
        RECT 2917.600 1560.410 2924.800 1560.860 ;
        RECT 2900.825 1560.110 2924.800 1560.410 ;
        RECT 2900.825 1560.095 2901.155 1560.110 ;
        RECT 2917.600 1559.660 2924.800 1560.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.370 1821.960 393.690 1822.020 ;
        RECT 2900.830 1821.960 2901.150 1822.020 ;
        RECT 393.370 1821.820 2901.150 1821.960 ;
        RECT 393.370 1821.760 393.690 1821.820 ;
        RECT 2900.830 1821.760 2901.150 1821.820 ;
      LAYER via ;
        RECT 393.400 1821.760 393.660 1822.020 ;
        RECT 2900.860 1821.760 2901.120 1822.020 ;
      LAYER met2 ;
        RECT 2900.850 1825.275 2901.130 1825.645 ;
        RECT 2900.920 1822.050 2901.060 1825.275 ;
        RECT 393.400 1821.730 393.660 1822.050 ;
        RECT 2900.860 1821.730 2901.120 1822.050 ;
        RECT 393.460 1048.870 393.600 1821.730 ;
        RECT 393.460 1048.730 395.440 1048.870 ;
        RECT 395.300 999.330 395.440 1048.730 ;
        RECT 396.970 999.330 397.250 1000.000 ;
        RECT 395.300 999.190 397.250 999.330 ;
        RECT 396.970 996.000 397.250 999.190 ;
      LAYER via2 ;
        RECT 2900.850 1825.320 2901.130 1825.600 ;
      LAYER met3 ;
        RECT 2900.825 1825.610 2901.155 1825.625 ;
        RECT 2917.600 1825.610 2924.800 1826.060 ;
        RECT 2900.825 1825.310 2924.800 1825.610 ;
        RECT 2900.825 1825.295 2901.155 1825.310 ;
        RECT 2917.600 1824.860 2924.800 1825.310 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 2090.900 414.390 2090.960 ;
        RECT 2900.830 2090.900 2901.150 2090.960 ;
        RECT 414.070 2090.760 2901.150 2090.900 ;
        RECT 414.070 2090.700 414.390 2090.760 ;
        RECT 2900.830 2090.700 2901.150 2090.760 ;
      LAYER via ;
        RECT 414.100 2090.700 414.360 2090.960 ;
        RECT 2900.860 2090.700 2901.120 2090.960 ;
      LAYER met2 ;
        RECT 2900.850 2091.155 2901.130 2091.525 ;
        RECT 2900.920 2090.990 2901.060 2091.155 ;
        RECT 414.100 2090.670 414.360 2090.990 ;
        RECT 2900.860 2090.670 2901.120 2090.990 ;
        RECT 414.160 1048.870 414.300 2090.670 ;
        RECT 414.160 1048.730 417.520 1048.870 ;
        RECT 417.380 999.330 417.520 1048.730 ;
        RECT 419.510 999.330 419.790 1000.000 ;
        RECT 417.380 999.190 419.790 999.330 ;
        RECT 419.510 996.000 419.790 999.190 ;
      LAYER via2 ;
        RECT 2900.850 2091.200 2901.130 2091.480 ;
      LAYER met3 ;
        RECT 2900.825 2091.490 2901.155 2091.505 ;
        RECT 2917.600 2091.490 2924.800 2091.940 ;
        RECT 2900.825 2091.190 2924.800 2091.490 ;
        RECT 2900.825 2091.175 2901.155 2091.190 ;
        RECT 2917.600 2090.740 2924.800 2091.190 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1053.010 1008.000 1053.330 1008.060 ;
        RECT 1104.530 1008.000 1104.850 1008.060 ;
        RECT 1053.010 1007.860 1104.850 1008.000 ;
        RECT 1053.010 1007.800 1053.330 1007.860 ;
        RECT 1104.530 1007.800 1104.850 1007.860 ;
        RECT 1104.530 403.480 1104.850 403.540 ;
        RECT 627.600 403.340 1104.850 403.480 ;
        RECT 627.600 403.200 627.740 403.340 ;
        RECT 1104.530 403.280 1104.850 403.340 ;
        RECT 627.510 402.940 627.830 403.200 ;
        RECT 386.930 385.800 387.250 385.860 ;
        RECT 391.530 385.800 391.850 385.860 ;
        RECT 386.930 385.660 391.850 385.800 ;
        RECT 386.930 385.600 387.250 385.660 ;
        RECT 391.530 385.600 391.850 385.660 ;
        RECT 386.930 30.840 387.250 30.900 ;
        RECT 573.230 30.840 573.550 30.900 ;
        RECT 386.930 30.700 573.550 30.840 ;
        RECT 386.930 30.640 387.250 30.700 ;
        RECT 573.230 30.640 573.550 30.700 ;
        RECT 573.230 20.300 573.550 20.360 ;
        RECT 627.510 20.300 627.830 20.360 ;
        RECT 573.230 20.160 627.830 20.300 ;
        RECT 573.230 20.100 573.550 20.160 ;
        RECT 627.510 20.100 627.830 20.160 ;
      LAYER via ;
        RECT 1053.040 1007.800 1053.300 1008.060 ;
        RECT 1104.560 1007.800 1104.820 1008.060 ;
        RECT 1104.560 403.280 1104.820 403.540 ;
        RECT 627.540 402.940 627.800 403.200 ;
        RECT 386.960 385.600 387.220 385.860 ;
        RECT 391.560 385.600 391.820 385.860 ;
        RECT 386.960 30.640 387.220 30.900 ;
        RECT 573.260 30.640 573.520 30.900 ;
        RECT 573.260 20.100 573.520 20.360 ;
        RECT 627.540 20.100 627.800 20.360 ;
      LAYER met2 ;
        RECT 1053.040 1007.770 1053.300 1008.090 ;
        RECT 1104.560 1007.770 1104.820 1008.090 ;
        RECT 1051.550 999.330 1051.830 1000.000 ;
        RECT 1053.100 999.330 1053.240 1007.770 ;
        RECT 1051.550 999.190 1053.240 999.330 ;
        RECT 1051.550 996.000 1051.830 999.190 ;
        RECT 392.830 400.250 393.110 404.000 ;
        RECT 1104.620 403.570 1104.760 1007.770 ;
        RECT 1104.560 403.250 1104.820 403.570 ;
        RECT 627.540 402.910 627.800 403.230 ;
        RECT 391.620 400.110 393.110 400.250 ;
        RECT 391.620 385.890 391.760 400.110 ;
        RECT 392.830 400.000 393.110 400.110 ;
        RECT 386.960 385.570 387.220 385.890 ;
        RECT 391.560 385.570 391.820 385.890 ;
        RECT 387.020 30.930 387.160 385.570 ;
        RECT 386.960 30.610 387.220 30.930 ;
        RECT 573.260 30.610 573.520 30.930 ;
        RECT 573.320 20.390 573.460 30.610 ;
        RECT 627.600 20.390 627.740 402.910 ;
        RECT 573.260 20.070 573.520 20.390 ;
        RECT 627.540 20.070 627.800 20.390 ;
        RECT 627.600 18.090 627.740 20.070 ;
        RECT 627.600 17.950 628.200 18.090 ;
        RECT 628.060 1.770 628.200 17.950 ;
        RECT 629.230 1.770 629.790 2.400 ;
        RECT 628.060 1.630 629.790 1.770 ;
        RECT 629.230 -4.800 629.790 1.630 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.950 109.040 933.270 109.100 ;
        RECT 2401.270 109.040 2401.590 109.100 ;
        RECT 932.950 108.900 2401.590 109.040 ;
        RECT 932.950 108.840 933.270 108.900 ;
        RECT 2401.270 108.840 2401.590 108.900 ;
      LAYER via ;
        RECT 932.980 108.840 933.240 109.100 ;
        RECT 2401.300 108.840 2401.560 109.100 ;
      LAYER met2 ;
        RECT 937.010 400.250 937.290 404.000 ;
        RECT 935.800 400.110 937.290 400.250 ;
        RECT 935.800 324.370 935.940 400.110 ;
        RECT 937.010 400.000 937.290 400.110 ;
        RECT 933.040 324.230 935.940 324.370 ;
        RECT 933.040 109.130 933.180 324.230 ;
        RECT 932.980 108.810 933.240 109.130 ;
        RECT 2401.300 108.810 2401.560 109.130 ;
        RECT 2401.360 82.870 2401.500 108.810 ;
        RECT 2401.360 82.730 2402.880 82.870 ;
        RECT 2402.740 2.400 2402.880 82.730 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 939.850 108.700 940.170 108.760 ;
        RECT 2415.070 108.700 2415.390 108.760 ;
        RECT 939.850 108.560 2415.390 108.700 ;
        RECT 939.850 108.500 940.170 108.560 ;
        RECT 2415.070 108.500 2415.390 108.560 ;
      LAYER via ;
        RECT 939.880 108.500 940.140 108.760 ;
        RECT 2415.100 108.500 2415.360 108.760 ;
      LAYER met2 ;
        RECT 942.530 400.250 942.810 404.000 ;
        RECT 941.320 400.110 942.810 400.250 ;
        RECT 941.320 324.370 941.460 400.110 ;
        RECT 942.530 400.000 942.810 400.110 ;
        RECT 939.940 324.230 941.460 324.370 ;
        RECT 939.940 108.790 940.080 324.230 ;
        RECT 939.880 108.470 940.140 108.790 ;
        RECT 2415.100 108.470 2415.360 108.790 ;
        RECT 2415.160 82.870 2415.300 108.470 ;
        RECT 2415.160 82.730 2420.360 82.870 ;
        RECT 2420.220 2.400 2420.360 82.730 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.750 108.360 947.070 108.420 ;
        RECT 2435.770 108.360 2436.090 108.420 ;
        RECT 946.750 108.220 2436.090 108.360 ;
        RECT 946.750 108.160 947.070 108.220 ;
        RECT 2435.770 108.160 2436.090 108.220 ;
      LAYER via ;
        RECT 946.780 108.160 947.040 108.420 ;
        RECT 2435.800 108.160 2436.060 108.420 ;
      LAYER met2 ;
        RECT 948.050 400.250 948.330 404.000 ;
        RECT 946.840 400.110 948.330 400.250 ;
        RECT 946.840 108.450 946.980 400.110 ;
        RECT 948.050 400.000 948.330 400.110 ;
        RECT 946.780 108.130 947.040 108.450 ;
        RECT 2435.800 108.130 2436.060 108.450 ;
        RECT 2435.860 1.770 2436.000 108.130 ;
        RECT 2437.950 1.770 2438.510 2.400 ;
        RECT 2435.860 1.630 2438.510 1.770 ;
        RECT 2437.950 -4.800 2438.510 1.630 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 953.190 108.020 953.510 108.080 ;
        RECT 2449.570 108.020 2449.890 108.080 ;
        RECT 953.190 107.880 2449.890 108.020 ;
        RECT 953.190 107.820 953.510 107.880 ;
        RECT 2449.570 107.820 2449.890 107.880 ;
        RECT 2449.570 17.580 2449.890 17.640 ;
        RECT 2453.710 17.580 2454.030 17.640 ;
        RECT 2449.570 17.440 2454.030 17.580 ;
        RECT 2449.570 17.380 2449.890 17.440 ;
        RECT 2453.710 17.380 2454.030 17.440 ;
      LAYER via ;
        RECT 953.220 107.820 953.480 108.080 ;
        RECT 2449.600 107.820 2449.860 108.080 ;
        RECT 2449.600 17.380 2449.860 17.640 ;
        RECT 2453.740 17.380 2454.000 17.640 ;
      LAYER met2 ;
        RECT 953.570 400.180 953.850 404.000 ;
        RECT 953.570 400.000 953.880 400.180 ;
        RECT 953.740 324.370 953.880 400.000 ;
        RECT 953.280 324.230 953.880 324.370 ;
        RECT 953.280 108.110 953.420 324.230 ;
        RECT 953.220 107.790 953.480 108.110 ;
        RECT 2449.600 107.790 2449.860 108.110 ;
        RECT 2449.660 17.670 2449.800 107.790 ;
        RECT 2449.600 17.350 2449.860 17.670 ;
        RECT 2453.740 17.350 2454.000 17.670 ;
        RECT 2453.800 1.770 2453.940 17.350 ;
        RECT 2455.430 1.770 2455.990 2.400 ;
        RECT 2453.800 1.630 2455.990 1.770 ;
        RECT 2455.430 -4.800 2455.990 1.630 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.170 22.340 959.490 22.400 ;
        RECT 2473.490 22.340 2473.810 22.400 ;
        RECT 959.170 22.200 2473.810 22.340 ;
        RECT 959.170 22.140 959.490 22.200 ;
        RECT 2473.490 22.140 2473.810 22.200 ;
      LAYER via ;
        RECT 959.200 22.140 959.460 22.400 ;
        RECT 2473.520 22.140 2473.780 22.400 ;
      LAYER met2 ;
        RECT 959.090 400.180 959.370 404.000 ;
        RECT 959.090 400.000 959.400 400.180 ;
        RECT 959.260 22.430 959.400 400.000 ;
        RECT 959.200 22.110 959.460 22.430 ;
        RECT 2473.520 22.110 2473.780 22.430 ;
        RECT 2473.580 2.400 2473.720 22.110 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 959.630 386.480 959.950 386.540 ;
        RECT 963.310 386.480 963.630 386.540 ;
        RECT 959.630 386.340 963.630 386.480 ;
        RECT 959.630 386.280 959.950 386.340 ;
        RECT 963.310 386.280 963.630 386.340 ;
        RECT 959.630 22.680 959.950 22.740 ;
        RECT 2490.970 22.680 2491.290 22.740 ;
        RECT 959.630 22.540 2491.290 22.680 ;
        RECT 959.630 22.480 959.950 22.540 ;
        RECT 2490.970 22.480 2491.290 22.540 ;
      LAYER via ;
        RECT 959.660 386.280 959.920 386.540 ;
        RECT 963.340 386.280 963.600 386.540 ;
        RECT 959.660 22.480 959.920 22.740 ;
        RECT 2491.000 22.480 2491.260 22.740 ;
      LAYER met2 ;
        RECT 964.610 400.250 964.890 404.000 ;
        RECT 963.400 400.110 964.890 400.250 ;
        RECT 963.400 386.570 963.540 400.110 ;
        RECT 964.610 400.000 964.890 400.110 ;
        RECT 959.660 386.250 959.920 386.570 ;
        RECT 963.340 386.250 963.600 386.570 ;
        RECT 959.720 22.770 959.860 386.250 ;
        RECT 959.660 22.450 959.920 22.770 ;
        RECT 2491.000 22.450 2491.260 22.770 ;
        RECT 2491.060 2.400 2491.200 22.450 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.070 386.480 966.390 386.540 ;
        RECT 968.370 386.480 968.690 386.540 ;
        RECT 966.070 386.340 968.690 386.480 ;
        RECT 966.070 386.280 966.390 386.340 ;
        RECT 968.370 386.280 968.690 386.340 ;
        RECT 966.530 23.020 966.850 23.080 ;
        RECT 2508.910 23.020 2509.230 23.080 ;
        RECT 966.530 22.880 2509.230 23.020 ;
        RECT 966.530 22.820 966.850 22.880 ;
        RECT 2508.910 22.820 2509.230 22.880 ;
      LAYER via ;
        RECT 966.100 386.280 966.360 386.540 ;
        RECT 968.400 386.280 968.660 386.540 ;
        RECT 966.560 22.820 966.820 23.080 ;
        RECT 2508.940 22.820 2509.200 23.080 ;
      LAYER met2 ;
        RECT 969.670 400.250 969.950 404.000 ;
        RECT 968.460 400.110 969.950 400.250 ;
        RECT 968.460 386.570 968.600 400.110 ;
        RECT 969.670 400.000 969.950 400.110 ;
        RECT 966.100 386.250 966.360 386.570 ;
        RECT 968.400 386.250 968.660 386.570 ;
        RECT 966.160 34.570 966.300 386.250 ;
        RECT 966.160 34.430 966.760 34.570 ;
        RECT 966.620 23.110 966.760 34.430 ;
        RECT 966.560 22.790 966.820 23.110 ;
        RECT 2508.940 22.790 2509.200 23.110 ;
        RECT 2509.000 2.400 2509.140 22.790 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 972.970 23.360 973.290 23.420 ;
        RECT 2526.850 23.360 2527.170 23.420 ;
        RECT 972.970 23.220 2527.170 23.360 ;
        RECT 972.970 23.160 973.290 23.220 ;
        RECT 2526.850 23.160 2527.170 23.220 ;
      LAYER via ;
        RECT 973.000 23.160 973.260 23.420 ;
        RECT 2526.880 23.160 2527.140 23.420 ;
      LAYER met2 ;
        RECT 975.190 400.250 975.470 404.000 ;
        RECT 973.980 400.110 975.470 400.250 ;
        RECT 973.980 387.330 974.120 400.110 ;
        RECT 975.190 400.000 975.470 400.110 ;
        RECT 973.060 387.190 974.120 387.330 ;
        RECT 973.060 23.450 973.200 387.190 ;
        RECT 973.000 23.130 973.260 23.450 ;
        RECT 2526.880 23.130 2527.140 23.450 ;
        RECT 2526.940 2.400 2527.080 23.130 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 979.870 23.700 980.190 23.760 ;
        RECT 2544.330 23.700 2544.650 23.760 ;
        RECT 979.870 23.560 2544.650 23.700 ;
        RECT 979.870 23.500 980.190 23.560 ;
        RECT 2544.330 23.500 2544.650 23.560 ;
      LAYER via ;
        RECT 979.900 23.500 980.160 23.760 ;
        RECT 2544.360 23.500 2544.620 23.760 ;
      LAYER met2 ;
        RECT 980.710 400.250 980.990 404.000 ;
        RECT 979.960 400.110 980.990 400.250 ;
        RECT 979.960 23.790 980.100 400.110 ;
        RECT 980.710 400.000 980.990 400.110 ;
        RECT 979.900 23.470 980.160 23.790 ;
        RECT 2544.360 23.470 2544.620 23.790 ;
        RECT 2544.420 2.400 2544.560 23.470 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.330 386.140 980.650 386.200 ;
        RECT 984.930 386.140 985.250 386.200 ;
        RECT 980.330 386.000 985.250 386.140 ;
        RECT 980.330 385.940 980.650 386.000 ;
        RECT 984.930 385.940 985.250 386.000 ;
        RECT 980.330 27.440 980.650 27.500 ;
        RECT 2562.270 27.440 2562.590 27.500 ;
        RECT 980.330 27.300 2562.590 27.440 ;
        RECT 980.330 27.240 980.650 27.300 ;
        RECT 2562.270 27.240 2562.590 27.300 ;
      LAYER via ;
        RECT 980.360 385.940 980.620 386.200 ;
        RECT 984.960 385.940 985.220 386.200 ;
        RECT 980.360 27.240 980.620 27.500 ;
        RECT 2562.300 27.240 2562.560 27.500 ;
      LAYER met2 ;
        RECT 986.230 400.250 986.510 404.000 ;
        RECT 985.020 400.110 986.510 400.250 ;
        RECT 985.020 386.230 985.160 400.110 ;
        RECT 986.230 400.000 986.510 400.110 ;
        RECT 980.360 385.910 980.620 386.230 ;
        RECT 984.960 385.910 985.220 386.230 ;
        RECT 980.420 27.530 980.560 385.910 ;
        RECT 980.360 27.210 980.620 27.530 ;
        RECT 2562.300 27.210 2562.560 27.530 ;
        RECT 2562.360 2.400 2562.500 27.210 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.130 386.480 442.450 386.540 ;
        RECT 445.810 386.480 446.130 386.540 ;
        RECT 442.130 386.340 446.130 386.480 ;
        RECT 442.130 386.280 442.450 386.340 ;
        RECT 445.810 386.280 446.130 386.340 ;
        RECT 442.130 28.460 442.450 28.520 ;
        RECT 586.110 28.460 586.430 28.520 ;
        RECT 442.130 28.320 586.430 28.460 ;
        RECT 442.130 28.260 442.450 28.320 ;
        RECT 586.110 28.260 586.430 28.320 ;
        RECT 586.110 19.960 586.430 20.020 ;
        RECT 806.450 19.960 806.770 20.020 ;
        RECT 586.110 19.820 806.770 19.960 ;
        RECT 586.110 19.760 586.430 19.820 ;
        RECT 806.450 19.760 806.770 19.820 ;
      LAYER via ;
        RECT 442.160 386.280 442.420 386.540 ;
        RECT 445.840 386.280 446.100 386.540 ;
        RECT 442.160 28.260 442.420 28.520 ;
        RECT 586.140 28.260 586.400 28.520 ;
        RECT 586.140 19.760 586.400 20.020 ;
        RECT 806.480 19.760 806.740 20.020 ;
      LAYER met2 ;
        RECT 447.110 400.250 447.390 404.000 ;
        RECT 445.900 400.110 447.390 400.250 ;
        RECT 445.900 386.570 446.040 400.110 ;
        RECT 447.110 400.000 447.390 400.110 ;
        RECT 442.160 386.250 442.420 386.570 ;
        RECT 445.840 386.250 446.100 386.570 ;
        RECT 442.220 28.550 442.360 386.250 ;
        RECT 442.160 28.230 442.420 28.550 ;
        RECT 586.140 28.230 586.400 28.550 ;
        RECT 586.200 20.050 586.340 28.230 ;
        RECT 586.140 19.730 586.400 20.050 ;
        RECT 806.480 19.730 806.740 20.050 ;
        RECT 806.540 2.400 806.680 19.730 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 986.770 386.140 987.090 386.200 ;
        RECT 990.450 386.140 990.770 386.200 ;
        RECT 986.770 386.000 990.770 386.140 ;
        RECT 986.770 385.940 987.090 386.000 ;
        RECT 990.450 385.940 990.770 386.000 ;
        RECT 986.770 27.100 987.090 27.160 ;
        RECT 2579.750 27.100 2580.070 27.160 ;
        RECT 986.770 26.960 2580.070 27.100 ;
        RECT 986.770 26.900 987.090 26.960 ;
        RECT 2579.750 26.900 2580.070 26.960 ;
      LAYER via ;
        RECT 986.800 385.940 987.060 386.200 ;
        RECT 990.480 385.940 990.740 386.200 ;
        RECT 986.800 26.900 987.060 27.160 ;
        RECT 2579.780 26.900 2580.040 27.160 ;
      LAYER met2 ;
        RECT 991.750 400.250 992.030 404.000 ;
        RECT 990.540 400.110 992.030 400.250 ;
        RECT 990.540 386.230 990.680 400.110 ;
        RECT 991.750 400.000 992.030 400.110 ;
        RECT 986.800 385.910 987.060 386.230 ;
        RECT 990.480 385.910 990.740 386.230 ;
        RECT 986.860 27.190 987.000 385.910 ;
        RECT 986.800 26.870 987.060 27.190 ;
        RECT 2579.780 26.870 2580.040 27.190 ;
        RECT 2579.840 2.400 2579.980 26.870 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 993.670 386.140 993.990 386.200 ;
        RECT 995.970 386.140 996.290 386.200 ;
        RECT 993.670 386.000 996.290 386.140 ;
        RECT 993.670 385.940 993.990 386.000 ;
        RECT 995.970 385.940 996.290 386.000 ;
        RECT 993.670 26.760 993.990 26.820 ;
        RECT 2597.690 26.760 2598.010 26.820 ;
        RECT 993.670 26.620 2598.010 26.760 ;
        RECT 993.670 26.560 993.990 26.620 ;
        RECT 2597.690 26.560 2598.010 26.620 ;
      LAYER via ;
        RECT 993.700 385.940 993.960 386.200 ;
        RECT 996.000 385.940 996.260 386.200 ;
        RECT 993.700 26.560 993.960 26.820 ;
        RECT 2597.720 26.560 2597.980 26.820 ;
      LAYER met2 ;
        RECT 997.270 400.250 997.550 404.000 ;
        RECT 996.060 400.110 997.550 400.250 ;
        RECT 996.060 386.230 996.200 400.110 ;
        RECT 997.270 400.000 997.550 400.110 ;
        RECT 993.700 385.910 993.960 386.230 ;
        RECT 996.000 385.910 996.260 386.230 ;
        RECT 993.760 26.850 993.900 385.910 ;
        RECT 993.700 26.530 993.960 26.850 ;
        RECT 2597.720 26.530 2597.980 26.850 ;
        RECT 2597.780 2.400 2597.920 26.530 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.570 386.140 1000.890 386.200 ;
        RECT 1001.950 386.140 1002.270 386.200 ;
        RECT 1000.570 386.000 1002.270 386.140 ;
        RECT 1000.570 385.940 1000.890 386.000 ;
        RECT 1001.950 385.940 1002.270 386.000 ;
        RECT 1000.570 26.420 1000.890 26.480 ;
        RECT 2615.170 26.420 2615.490 26.480 ;
        RECT 1000.570 26.280 2615.490 26.420 ;
        RECT 1000.570 26.220 1000.890 26.280 ;
        RECT 2615.170 26.220 2615.490 26.280 ;
      LAYER via ;
        RECT 1000.600 385.940 1000.860 386.200 ;
        RECT 1001.980 385.940 1002.240 386.200 ;
        RECT 1000.600 26.220 1000.860 26.480 ;
        RECT 2615.200 26.220 2615.460 26.480 ;
      LAYER met2 ;
        RECT 1002.330 400.250 1002.610 404.000 ;
        RECT 1002.040 400.110 1002.610 400.250 ;
        RECT 1002.040 386.230 1002.180 400.110 ;
        RECT 1002.330 400.000 1002.610 400.110 ;
        RECT 1000.600 385.910 1000.860 386.230 ;
        RECT 1001.980 385.910 1002.240 386.230 ;
        RECT 1000.660 26.510 1000.800 385.910 ;
        RECT 1000.600 26.190 1000.860 26.510 ;
        RECT 2615.200 26.190 2615.460 26.510 ;
        RECT 2615.260 2.400 2615.400 26.190 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.470 26.080 1007.790 26.140 ;
        RECT 2633.110 26.080 2633.430 26.140 ;
        RECT 1007.470 25.940 2633.430 26.080 ;
        RECT 1007.470 25.880 1007.790 25.940 ;
        RECT 2633.110 25.880 2633.430 25.940 ;
      LAYER via ;
        RECT 1007.500 25.880 1007.760 26.140 ;
        RECT 2633.140 25.880 2633.400 26.140 ;
      LAYER met2 ;
        RECT 1007.850 400.250 1008.130 404.000 ;
        RECT 1007.560 400.110 1008.130 400.250 ;
        RECT 1007.560 26.170 1007.700 400.110 ;
        RECT 1007.850 400.000 1008.130 400.110 ;
        RECT 1007.500 25.850 1007.760 26.170 ;
        RECT 2633.140 25.850 2633.400 26.170 ;
        RECT 2633.200 2.400 2633.340 25.850 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1007.930 386.480 1008.250 386.540 ;
        RECT 1012.070 386.480 1012.390 386.540 ;
        RECT 1007.930 386.340 1012.390 386.480 ;
        RECT 1007.930 386.280 1008.250 386.340 ;
        RECT 1012.070 386.280 1012.390 386.340 ;
        RECT 1007.930 25.740 1008.250 25.800 ;
        RECT 2650.590 25.740 2650.910 25.800 ;
        RECT 1007.930 25.600 2650.910 25.740 ;
        RECT 1007.930 25.540 1008.250 25.600 ;
        RECT 2650.590 25.540 2650.910 25.600 ;
      LAYER via ;
        RECT 1007.960 386.280 1008.220 386.540 ;
        RECT 1012.100 386.280 1012.360 386.540 ;
        RECT 1007.960 25.540 1008.220 25.800 ;
        RECT 2650.620 25.540 2650.880 25.800 ;
      LAYER met2 ;
        RECT 1013.370 400.250 1013.650 404.000 ;
        RECT 1012.160 400.110 1013.650 400.250 ;
        RECT 1012.160 386.570 1012.300 400.110 ;
        RECT 1013.370 400.000 1013.650 400.110 ;
        RECT 1007.960 386.250 1008.220 386.570 ;
        RECT 1012.100 386.250 1012.360 386.570 ;
        RECT 1008.020 25.830 1008.160 386.250 ;
        RECT 1007.960 25.510 1008.220 25.830 ;
        RECT 2650.620 25.510 2650.880 25.830 ;
        RECT 2650.680 2.400 2650.820 25.510 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.370 386.140 1014.690 386.200 ;
        RECT 1017.590 386.140 1017.910 386.200 ;
        RECT 1014.370 386.000 1017.910 386.140 ;
        RECT 1014.370 385.940 1014.690 386.000 ;
        RECT 1017.590 385.940 1017.910 386.000 ;
        RECT 1014.370 25.400 1014.690 25.460 ;
        RECT 2668.530 25.400 2668.850 25.460 ;
        RECT 1014.370 25.260 2668.850 25.400 ;
        RECT 1014.370 25.200 1014.690 25.260 ;
        RECT 2668.530 25.200 2668.850 25.260 ;
      LAYER via ;
        RECT 1014.400 385.940 1014.660 386.200 ;
        RECT 1017.620 385.940 1017.880 386.200 ;
        RECT 1014.400 25.200 1014.660 25.460 ;
        RECT 2668.560 25.200 2668.820 25.460 ;
      LAYER met2 ;
        RECT 1018.890 400.250 1019.170 404.000 ;
        RECT 1017.680 400.110 1019.170 400.250 ;
        RECT 1017.680 386.230 1017.820 400.110 ;
        RECT 1018.890 400.000 1019.170 400.110 ;
        RECT 1014.400 385.910 1014.660 386.230 ;
        RECT 1017.620 385.910 1017.880 386.230 ;
        RECT 1014.460 25.490 1014.600 385.910 ;
        RECT 1014.400 25.170 1014.660 25.490 ;
        RECT 2668.560 25.170 2668.820 25.490 ;
        RECT 2668.620 2.400 2668.760 25.170 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.270 386.480 1021.590 386.540 ;
        RECT 1023.110 386.480 1023.430 386.540 ;
        RECT 1021.270 386.340 1023.430 386.480 ;
        RECT 1021.270 386.280 1021.590 386.340 ;
        RECT 1023.110 386.280 1023.430 386.340 ;
        RECT 1021.270 25.060 1021.590 25.120 ;
        RECT 2686.010 25.060 2686.330 25.120 ;
        RECT 1021.270 24.920 2686.330 25.060 ;
        RECT 1021.270 24.860 1021.590 24.920 ;
        RECT 2686.010 24.860 2686.330 24.920 ;
      LAYER via ;
        RECT 1021.300 386.280 1021.560 386.540 ;
        RECT 1023.140 386.280 1023.400 386.540 ;
        RECT 1021.300 24.860 1021.560 25.120 ;
        RECT 2686.040 24.860 2686.300 25.120 ;
      LAYER met2 ;
        RECT 1024.410 400.250 1024.690 404.000 ;
        RECT 1023.200 400.110 1024.690 400.250 ;
        RECT 1023.200 386.570 1023.340 400.110 ;
        RECT 1024.410 400.000 1024.690 400.110 ;
        RECT 1021.300 386.250 1021.560 386.570 ;
        RECT 1023.140 386.250 1023.400 386.570 ;
        RECT 1021.360 25.150 1021.500 386.250 ;
        RECT 1021.300 24.830 1021.560 25.150 ;
        RECT 2686.040 24.830 2686.300 25.150 ;
        RECT 2686.100 2.400 2686.240 24.830 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.170 24.720 1028.490 24.780 ;
        RECT 2703.950 24.720 2704.270 24.780 ;
        RECT 1028.170 24.580 2704.270 24.720 ;
        RECT 1028.170 24.520 1028.490 24.580 ;
        RECT 2703.950 24.520 2704.270 24.580 ;
      LAYER via ;
        RECT 1028.200 24.520 1028.460 24.780 ;
        RECT 2703.980 24.520 2704.240 24.780 ;
      LAYER met2 ;
        RECT 1029.930 401.610 1030.210 404.000 ;
        RECT 1029.180 401.470 1030.210 401.610 ;
        RECT 1029.180 389.370 1029.320 401.470 ;
        RECT 1029.930 400.000 1030.210 401.470 ;
        RECT 1028.720 389.230 1029.320 389.370 ;
        RECT 1028.720 388.010 1028.860 389.230 ;
        RECT 1028.260 387.870 1028.860 388.010 ;
        RECT 1028.260 24.810 1028.400 387.870 ;
        RECT 1028.200 24.490 1028.460 24.810 ;
        RECT 2703.980 24.490 2704.240 24.810 ;
        RECT 2704.040 2.400 2704.180 24.490 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.070 24.380 1035.390 24.440 ;
        RECT 2721.890 24.380 2722.210 24.440 ;
        RECT 1035.070 24.240 2722.210 24.380 ;
        RECT 1035.070 24.180 1035.390 24.240 ;
        RECT 2721.890 24.180 2722.210 24.240 ;
      LAYER via ;
        RECT 1035.100 24.180 1035.360 24.440 ;
        RECT 2721.920 24.180 2722.180 24.440 ;
      LAYER met2 ;
        RECT 1034.990 400.180 1035.270 404.000 ;
        RECT 1034.990 400.000 1035.300 400.180 ;
        RECT 1035.160 24.470 1035.300 400.000 ;
        RECT 1035.100 24.150 1035.360 24.470 ;
        RECT 2721.920 24.150 2722.180 24.470 ;
        RECT 2721.980 2.400 2722.120 24.150 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.530 376.280 1035.850 376.340 ;
        RECT 1039.210 376.280 1039.530 376.340 ;
        RECT 1035.530 376.140 1039.530 376.280 ;
        RECT 1035.530 376.080 1035.850 376.140 ;
        RECT 1039.210 376.080 1039.530 376.140 ;
      LAYER via ;
        RECT 1035.560 376.080 1035.820 376.340 ;
        RECT 1039.240 376.080 1039.500 376.340 ;
      LAYER met2 ;
        RECT 1040.510 400.250 1040.790 404.000 ;
        RECT 1039.300 400.110 1040.790 400.250 ;
        RECT 1039.300 376.370 1039.440 400.110 ;
        RECT 1040.510 400.000 1040.790 400.110 ;
        RECT 1035.560 376.050 1035.820 376.370 ;
        RECT 1039.240 376.050 1039.500 376.370 ;
        RECT 1035.620 24.325 1035.760 376.050 ;
        RECT 1035.550 23.955 1035.830 24.325 ;
        RECT 2739.390 23.955 2739.670 24.325 ;
        RECT 2739.460 2.400 2739.600 23.955 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
      LAYER via2 ;
        RECT 1035.550 24.000 1035.830 24.280 ;
        RECT 2739.390 24.000 2739.670 24.280 ;
      LAYER met3 ;
        RECT 1035.525 24.290 1035.855 24.305 ;
        RECT 2739.365 24.290 2739.695 24.305 ;
        RECT 1035.525 23.990 2739.695 24.290 ;
        RECT 1035.525 23.975 1035.855 23.990 ;
        RECT 2739.365 23.975 2739.695 23.990 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 452.710 389.540 453.030 389.600 ;
        RECT 596.690 389.540 597.010 389.600 ;
        RECT 452.710 389.400 597.010 389.540 ;
        RECT 452.710 389.340 453.030 389.400 ;
        RECT 596.690 389.340 597.010 389.400 ;
        RECT 596.690 19.620 597.010 19.680 ;
        RECT 824.390 19.620 824.710 19.680 ;
        RECT 596.690 19.480 824.710 19.620 ;
        RECT 596.690 19.420 597.010 19.480 ;
        RECT 824.390 19.420 824.710 19.480 ;
      LAYER via ;
        RECT 452.740 389.340 453.000 389.600 ;
        RECT 596.720 389.340 596.980 389.600 ;
        RECT 596.720 19.420 596.980 19.680 ;
        RECT 824.420 19.420 824.680 19.680 ;
      LAYER met2 ;
        RECT 452.630 400.180 452.910 404.000 ;
        RECT 452.630 400.000 452.940 400.180 ;
        RECT 452.800 389.630 452.940 400.000 ;
        RECT 452.740 389.310 453.000 389.630 ;
        RECT 596.720 389.310 596.980 389.630 ;
        RECT 596.780 19.710 596.920 389.310 ;
        RECT 596.720 19.390 596.980 19.710 ;
        RECT 824.420 19.390 824.680 19.710 ;
        RECT 824.480 2.400 824.620 19.390 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.970 376.280 1042.290 376.340 ;
        RECT 1044.730 376.280 1045.050 376.340 ;
        RECT 1041.970 376.140 1045.050 376.280 ;
        RECT 1041.970 376.080 1042.290 376.140 ;
        RECT 1044.730 376.080 1045.050 376.140 ;
        RECT 1041.970 24.040 1042.290 24.100 ;
        RECT 2757.310 24.040 2757.630 24.100 ;
        RECT 1041.970 23.900 2757.630 24.040 ;
        RECT 1041.970 23.840 1042.290 23.900 ;
        RECT 2757.310 23.840 2757.630 23.900 ;
      LAYER via ;
        RECT 1042.000 376.080 1042.260 376.340 ;
        RECT 1044.760 376.080 1045.020 376.340 ;
        RECT 1042.000 23.840 1042.260 24.100 ;
        RECT 2757.340 23.840 2757.600 24.100 ;
      LAYER met2 ;
        RECT 1046.030 400.250 1046.310 404.000 ;
        RECT 1044.820 400.110 1046.310 400.250 ;
        RECT 1044.820 376.370 1044.960 400.110 ;
        RECT 1046.030 400.000 1046.310 400.110 ;
        RECT 1042.000 376.050 1042.260 376.370 ;
        RECT 1044.760 376.050 1045.020 376.370 ;
        RECT 1042.060 24.130 1042.200 376.050 ;
        RECT 1042.000 23.810 1042.260 24.130 ;
        RECT 2757.340 23.810 2757.600 24.130 ;
        RECT 2757.400 2.400 2757.540 23.810 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1050.250 107.680 1050.570 107.740 ;
        RECT 2773.870 107.680 2774.190 107.740 ;
        RECT 1050.250 107.540 2774.190 107.680 ;
        RECT 1050.250 107.480 1050.570 107.540 ;
        RECT 2773.870 107.480 2774.190 107.540 ;
      LAYER via ;
        RECT 1050.280 107.480 1050.540 107.740 ;
        RECT 2773.900 107.480 2774.160 107.740 ;
      LAYER met2 ;
        RECT 1051.550 400.250 1051.830 404.000 ;
        RECT 1050.340 400.110 1051.830 400.250 ;
        RECT 1050.340 107.770 1050.480 400.110 ;
        RECT 1051.550 400.000 1051.830 400.110 ;
        RECT 1050.280 107.450 1050.540 107.770 ;
        RECT 2773.900 107.450 2774.160 107.770 ;
        RECT 2773.960 1.770 2774.100 107.450 ;
        RECT 2774.670 1.770 2775.230 2.400 ;
        RECT 2773.960 1.630 2775.230 1.770 ;
        RECT 2774.670 -4.800 2775.230 1.630 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1056.690 107.340 1057.010 107.400 ;
        RECT 2787.670 107.340 2787.990 107.400 ;
        RECT 1056.690 107.200 2787.990 107.340 ;
        RECT 1056.690 107.140 1057.010 107.200 ;
        RECT 2787.670 107.140 2787.990 107.200 ;
      LAYER via ;
        RECT 1056.720 107.140 1056.980 107.400 ;
        RECT 2787.700 107.140 2787.960 107.400 ;
      LAYER met2 ;
        RECT 1057.070 400.250 1057.350 404.000 ;
        RECT 1056.780 400.110 1057.350 400.250 ;
        RECT 1056.780 107.430 1056.920 400.110 ;
        RECT 1057.070 400.000 1057.350 400.110 ;
        RECT 1056.720 107.110 1056.980 107.430 ;
        RECT 2787.700 107.110 2787.960 107.430 ;
        RECT 2787.760 82.870 2787.900 107.110 ;
        RECT 2787.760 82.730 2792.960 82.870 ;
        RECT 2792.820 2.400 2792.960 82.730 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.590 327.800 1063.910 328.060 ;
        RECT 1063.680 327.040 1063.820 327.800 ;
        RECT 1063.590 326.780 1063.910 327.040 ;
        RECT 1063.590 107.000 1063.910 107.060 ;
        RECT 2808.370 107.000 2808.690 107.060 ;
        RECT 1063.590 106.860 2808.690 107.000 ;
        RECT 1063.590 106.800 1063.910 106.860 ;
        RECT 2808.370 106.800 2808.690 106.860 ;
      LAYER via ;
        RECT 1063.620 327.800 1063.880 328.060 ;
        RECT 1063.620 326.780 1063.880 327.040 ;
        RECT 1063.620 106.800 1063.880 107.060 ;
        RECT 2808.400 106.800 2808.660 107.060 ;
      LAYER met2 ;
        RECT 1062.590 400.250 1062.870 404.000 ;
        RECT 1062.590 400.110 1063.820 400.250 ;
        RECT 1062.590 400.000 1062.870 400.110 ;
        RECT 1063.680 328.090 1063.820 400.110 ;
        RECT 1063.620 327.770 1063.880 328.090 ;
        RECT 1063.620 326.750 1063.880 327.070 ;
        RECT 1063.680 107.090 1063.820 326.750 ;
        RECT 1063.620 106.770 1063.880 107.090 ;
        RECT 2808.400 106.770 2808.660 107.090 ;
        RECT 2808.460 82.870 2808.600 106.770 ;
        RECT 2808.460 82.730 2810.440 82.870 ;
        RECT 2810.300 2.400 2810.440 82.730 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1067.730 391.920 1068.050 391.980 ;
        RECT 2218.190 391.920 2218.510 391.980 ;
        RECT 1067.730 391.780 2218.510 391.920 ;
        RECT 1067.730 391.720 1068.050 391.780 ;
        RECT 2218.190 391.720 2218.510 391.780 ;
        RECT 2828.150 16.900 2828.470 16.960 ;
        RECT 2256.230 16.760 2828.470 16.900 ;
        RECT 2218.190 16.560 2218.510 16.620 ;
        RECT 2256.230 16.560 2256.370 16.760 ;
        RECT 2828.150 16.700 2828.470 16.760 ;
        RECT 2218.190 16.420 2256.370 16.560 ;
        RECT 2218.190 16.360 2218.510 16.420 ;
      LAYER via ;
        RECT 1067.760 391.720 1068.020 391.980 ;
        RECT 2218.220 391.720 2218.480 391.980 ;
        RECT 2218.220 16.360 2218.480 16.620 ;
        RECT 2828.180 16.700 2828.440 16.960 ;
      LAYER met2 ;
        RECT 1067.650 400.180 1067.930 404.000 ;
        RECT 1067.650 400.000 1067.960 400.180 ;
        RECT 1067.820 392.010 1067.960 400.000 ;
        RECT 1067.760 391.690 1068.020 392.010 ;
        RECT 2218.220 391.690 2218.480 392.010 ;
        RECT 2218.280 16.650 2218.420 391.690 ;
        RECT 2828.180 16.670 2828.440 16.990 ;
        RECT 2218.220 16.330 2218.480 16.650 ;
        RECT 2828.240 2.400 2828.380 16.670 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1069.570 375.940 1069.890 376.000 ;
        RECT 1071.870 375.940 1072.190 376.000 ;
        RECT 1069.570 375.800 1072.190 375.940 ;
        RECT 1069.570 375.740 1069.890 375.800 ;
        RECT 1071.870 375.740 1072.190 375.800 ;
        RECT 1069.570 32.200 1069.890 32.260 ;
        RECT 2845.630 32.200 2845.950 32.260 ;
        RECT 1069.570 32.060 2845.950 32.200 ;
        RECT 1069.570 32.000 1069.890 32.060 ;
        RECT 2845.630 32.000 2845.950 32.060 ;
      LAYER via ;
        RECT 1069.600 375.740 1069.860 376.000 ;
        RECT 1071.900 375.740 1072.160 376.000 ;
        RECT 1069.600 32.000 1069.860 32.260 ;
        RECT 2845.660 32.000 2845.920 32.260 ;
      LAYER met2 ;
        RECT 1073.170 400.250 1073.450 404.000 ;
        RECT 1071.960 400.110 1073.450 400.250 ;
        RECT 1071.960 376.030 1072.100 400.110 ;
        RECT 1073.170 400.000 1073.450 400.110 ;
        RECT 1069.600 375.710 1069.860 376.030 ;
        RECT 1071.900 375.710 1072.160 376.030 ;
        RECT 1069.660 32.290 1069.800 375.710 ;
        RECT 1069.600 31.970 1069.860 32.290 ;
        RECT 2845.660 31.970 2845.920 32.290 ;
        RECT 2845.720 2.400 2845.860 31.970 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.470 376.280 1076.790 376.340 ;
        RECT 1077.850 376.280 1078.170 376.340 ;
        RECT 1076.470 376.140 1078.170 376.280 ;
        RECT 1076.470 376.080 1076.790 376.140 ;
        RECT 1077.850 376.080 1078.170 376.140 ;
        RECT 1076.470 31.520 1076.790 31.580 ;
        RECT 2863.570 31.520 2863.890 31.580 ;
        RECT 1076.470 31.380 2863.890 31.520 ;
        RECT 1076.470 31.320 1076.790 31.380 ;
        RECT 2863.570 31.320 2863.890 31.380 ;
      LAYER via ;
        RECT 1076.500 376.080 1076.760 376.340 ;
        RECT 1077.880 376.080 1078.140 376.340 ;
        RECT 1076.500 31.320 1076.760 31.580 ;
        RECT 2863.600 31.320 2863.860 31.580 ;
      LAYER met2 ;
        RECT 1078.690 400.250 1078.970 404.000 ;
        RECT 1077.940 400.110 1078.970 400.250 ;
        RECT 1077.940 376.370 1078.080 400.110 ;
        RECT 1078.690 400.000 1078.970 400.110 ;
        RECT 1076.500 376.050 1076.760 376.370 ;
        RECT 1077.880 376.050 1078.140 376.370 ;
        RECT 1076.560 31.610 1076.700 376.050 ;
        RECT 1076.500 31.290 1076.760 31.610 ;
        RECT 2863.600 31.290 2863.860 31.610 ;
        RECT 2863.660 2.400 2863.800 31.290 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.750 31.180 1085.070 31.240 ;
        RECT 2881.510 31.180 2881.830 31.240 ;
        RECT 1084.750 31.040 2881.830 31.180 ;
        RECT 1084.750 30.980 1085.070 31.040 ;
        RECT 2881.510 30.980 2881.830 31.040 ;
      LAYER via ;
        RECT 1084.780 30.980 1085.040 31.240 ;
        RECT 2881.540 30.980 2881.800 31.240 ;
      LAYER met2 ;
        RECT 1084.210 400.180 1084.490 404.000 ;
        RECT 1084.210 400.000 1084.520 400.180 ;
        RECT 1084.380 34.570 1084.520 400.000 ;
        RECT 1084.380 34.430 1084.980 34.570 ;
        RECT 1084.840 31.270 1084.980 34.430 ;
        RECT 1084.780 30.950 1085.040 31.270 ;
        RECT 2881.540 30.950 2881.800 31.270 ;
        RECT 2881.600 2.400 2881.740 30.950 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 458.230 388.860 458.550 388.920 ;
        RECT 597.150 388.860 597.470 388.920 ;
        RECT 458.230 388.720 597.470 388.860 ;
        RECT 458.230 388.660 458.550 388.720 ;
        RECT 597.150 388.660 597.470 388.720 ;
        RECT 597.150 17.920 597.470 17.980 ;
        RECT 841.870 17.920 842.190 17.980 ;
        RECT 597.150 17.780 842.190 17.920 ;
        RECT 597.150 17.720 597.470 17.780 ;
        RECT 841.870 17.720 842.190 17.780 ;
      LAYER via ;
        RECT 458.260 388.660 458.520 388.920 ;
        RECT 597.180 388.660 597.440 388.920 ;
        RECT 597.180 17.720 597.440 17.980 ;
        RECT 841.900 17.720 842.160 17.980 ;
      LAYER met2 ;
        RECT 458.150 400.180 458.430 404.000 ;
        RECT 458.150 400.000 458.460 400.180 ;
        RECT 458.320 388.950 458.460 400.000 ;
        RECT 458.260 388.630 458.520 388.950 ;
        RECT 597.180 388.630 597.440 388.950 ;
        RECT 597.240 18.010 597.380 388.630 ;
        RECT 597.180 17.690 597.440 18.010 ;
        RECT 841.900 17.690 842.160 18.010 ;
        RECT 841.960 2.400 842.100 17.690 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 388.520 462.690 388.580 ;
        RECT 597.610 388.520 597.930 388.580 ;
        RECT 462.370 388.380 597.930 388.520 ;
        RECT 462.370 388.320 462.690 388.380 ;
        RECT 597.610 388.320 597.930 388.380 ;
        RECT 597.610 17.580 597.930 17.640 ;
        RECT 859.810 17.580 860.130 17.640 ;
        RECT 597.610 17.440 860.130 17.580 ;
        RECT 597.610 17.380 597.930 17.440 ;
        RECT 859.810 17.380 860.130 17.440 ;
      LAYER via ;
        RECT 462.400 388.320 462.660 388.580 ;
        RECT 597.640 388.320 597.900 388.580 ;
        RECT 597.640 17.380 597.900 17.640 ;
        RECT 859.840 17.380 860.100 17.640 ;
      LAYER met2 ;
        RECT 463.670 400.250 463.950 404.000 ;
        RECT 462.460 400.110 463.950 400.250 ;
        RECT 462.460 388.610 462.600 400.110 ;
        RECT 463.670 400.000 463.950 400.110 ;
        RECT 462.400 388.290 462.660 388.610 ;
        RECT 597.640 388.290 597.900 388.610 ;
        RECT 597.700 17.670 597.840 388.290 ;
        RECT 597.640 17.350 597.900 17.670 ;
        RECT 859.840 17.350 860.100 17.670 ;
        RECT 859.900 2.400 860.040 17.350 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.370 376.280 462.690 376.340 ;
        RECT 467.430 376.280 467.750 376.340 ;
        RECT 462.370 376.140 467.750 376.280 ;
        RECT 462.370 376.080 462.690 376.140 ;
        RECT 467.430 376.080 467.750 376.140 ;
        RECT 462.370 26.420 462.690 26.480 ;
        RECT 877.290 26.420 877.610 26.480 ;
        RECT 462.370 26.280 877.610 26.420 ;
        RECT 462.370 26.220 462.690 26.280 ;
        RECT 877.290 26.220 877.610 26.280 ;
      LAYER via ;
        RECT 462.400 376.080 462.660 376.340 ;
        RECT 467.460 376.080 467.720 376.340 ;
        RECT 462.400 26.220 462.660 26.480 ;
        RECT 877.320 26.220 877.580 26.480 ;
      LAYER met2 ;
        RECT 468.730 400.250 469.010 404.000 ;
        RECT 467.520 400.110 469.010 400.250 ;
        RECT 467.520 376.370 467.660 400.110 ;
        RECT 468.730 400.000 469.010 400.110 ;
        RECT 462.400 376.050 462.660 376.370 ;
        RECT 467.460 376.050 467.720 376.370 ;
        RECT 462.460 26.510 462.600 376.050 ;
        RECT 462.400 26.190 462.660 26.510 ;
        RECT 877.320 26.190 877.580 26.510 ;
        RECT 877.380 2.400 877.520 26.190 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 474.330 392.940 474.650 393.000 ;
        RECT 516.190 392.940 516.510 393.000 ;
        RECT 474.330 392.800 516.510 392.940 ;
        RECT 474.330 392.740 474.650 392.800 ;
        RECT 516.190 392.740 516.510 392.800 ;
        RECT 516.190 389.200 516.510 389.260 ;
        RECT 610.030 389.200 610.350 389.260 ;
        RECT 516.190 389.060 610.350 389.200 ;
        RECT 516.190 389.000 516.510 389.060 ;
        RECT 610.030 389.000 610.350 389.060 ;
        RECT 610.490 17.240 610.810 17.300 ;
        RECT 895.230 17.240 895.550 17.300 ;
        RECT 610.490 17.100 895.550 17.240 ;
        RECT 610.490 17.040 610.810 17.100 ;
        RECT 895.230 17.040 895.550 17.100 ;
      LAYER via ;
        RECT 474.360 392.740 474.620 393.000 ;
        RECT 516.220 392.740 516.480 393.000 ;
        RECT 516.220 389.000 516.480 389.260 ;
        RECT 610.060 389.000 610.320 389.260 ;
        RECT 610.520 17.040 610.780 17.300 ;
        RECT 895.260 17.040 895.520 17.300 ;
      LAYER met2 ;
        RECT 474.250 400.180 474.530 404.000 ;
        RECT 474.250 400.000 474.560 400.180 ;
        RECT 474.420 393.030 474.560 400.000 ;
        RECT 474.360 392.710 474.620 393.030 ;
        RECT 516.220 392.710 516.480 393.030 ;
        RECT 516.280 389.290 516.420 392.710 ;
        RECT 516.220 388.970 516.480 389.290 ;
        RECT 610.060 388.970 610.320 389.290 ;
        RECT 610.120 351.970 610.260 388.970 ;
        RECT 610.120 351.830 610.720 351.970 ;
        RECT 610.580 17.330 610.720 351.830 ;
        RECT 610.520 17.010 610.780 17.330 ;
        RECT 895.260 17.010 895.520 17.330 ;
        RECT 895.320 2.400 895.460 17.010 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 376.280 476.490 376.340 ;
        RECT 478.470 376.280 478.790 376.340 ;
        RECT 476.170 376.140 478.790 376.280 ;
        RECT 476.170 376.080 476.490 376.140 ;
        RECT 478.470 376.080 478.790 376.140 ;
        RECT 476.170 26.080 476.490 26.140 ;
        RECT 912.710 26.080 913.030 26.140 ;
        RECT 476.170 25.940 913.030 26.080 ;
        RECT 476.170 25.880 476.490 25.940 ;
        RECT 912.710 25.880 913.030 25.940 ;
      LAYER via ;
        RECT 476.200 376.080 476.460 376.340 ;
        RECT 478.500 376.080 478.760 376.340 ;
        RECT 476.200 25.880 476.460 26.140 ;
        RECT 912.740 25.880 913.000 26.140 ;
      LAYER met2 ;
        RECT 479.770 400.250 480.050 404.000 ;
        RECT 478.560 400.110 480.050 400.250 ;
        RECT 478.560 376.370 478.700 400.110 ;
        RECT 479.770 400.000 480.050 400.110 ;
        RECT 476.200 376.050 476.460 376.370 ;
        RECT 478.500 376.050 478.760 376.370 ;
        RECT 476.260 26.170 476.400 376.050 ;
        RECT 476.200 25.850 476.460 26.170 ;
        RECT 912.740 25.850 913.000 26.170 ;
        RECT 912.800 2.400 912.940 25.850 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.070 382.060 483.390 382.120 ;
        RECT 485.370 382.060 485.690 382.120 ;
        RECT 483.070 381.920 485.690 382.060 ;
        RECT 483.070 381.860 483.390 381.920 ;
        RECT 485.370 381.860 485.690 381.920 ;
        RECT 483.070 25.740 483.390 25.800 ;
        RECT 930.650 25.740 930.970 25.800 ;
        RECT 483.070 25.600 930.970 25.740 ;
        RECT 483.070 25.540 483.390 25.600 ;
        RECT 930.650 25.540 930.970 25.600 ;
      LAYER via ;
        RECT 483.100 381.860 483.360 382.120 ;
        RECT 485.400 381.860 485.660 382.120 ;
        RECT 483.100 25.540 483.360 25.800 ;
        RECT 930.680 25.540 930.940 25.800 ;
      LAYER met2 ;
        RECT 485.290 400.180 485.570 404.000 ;
        RECT 485.290 400.000 485.600 400.180 ;
        RECT 485.460 382.150 485.600 400.000 ;
        RECT 483.100 381.830 483.360 382.150 ;
        RECT 485.400 381.830 485.660 382.150 ;
        RECT 483.160 25.830 483.300 381.830 ;
        RECT 483.100 25.510 483.360 25.830 ;
        RECT 930.680 25.510 930.940 25.830 ;
        RECT 930.740 2.400 930.880 25.510 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 25.400 490.290 25.460 ;
        RECT 948.590 25.400 948.910 25.460 ;
        RECT 489.970 25.260 948.910 25.400 ;
        RECT 489.970 25.200 490.290 25.260 ;
        RECT 948.590 25.200 948.910 25.260 ;
      LAYER via ;
        RECT 490.000 25.200 490.260 25.460 ;
        RECT 948.620 25.200 948.880 25.460 ;
      LAYER met2 ;
        RECT 490.810 400.250 491.090 404.000 ;
        RECT 490.060 400.110 491.090 400.250 ;
        RECT 490.060 25.490 490.200 400.110 ;
        RECT 490.810 400.000 491.090 400.110 ;
        RECT 490.000 25.170 490.260 25.490 ;
        RECT 948.620 25.170 948.880 25.490 ;
        RECT 948.680 2.400 948.820 25.170 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.430 376.280 490.750 376.340 ;
        RECT 495.030 376.280 495.350 376.340 ;
        RECT 490.430 376.140 495.350 376.280 ;
        RECT 490.430 376.080 490.750 376.140 ;
        RECT 495.030 376.080 495.350 376.140 ;
        RECT 490.430 25.060 490.750 25.120 ;
        RECT 966.070 25.060 966.390 25.120 ;
        RECT 490.430 24.920 966.390 25.060 ;
        RECT 490.430 24.860 490.750 24.920 ;
        RECT 966.070 24.860 966.390 24.920 ;
      LAYER via ;
        RECT 490.460 376.080 490.720 376.340 ;
        RECT 495.060 376.080 495.320 376.340 ;
        RECT 490.460 24.860 490.720 25.120 ;
        RECT 966.100 24.860 966.360 25.120 ;
      LAYER met2 ;
        RECT 496.330 400.250 496.610 404.000 ;
        RECT 495.120 400.110 496.610 400.250 ;
        RECT 495.120 376.370 495.260 400.110 ;
        RECT 496.330 400.000 496.610 400.110 ;
        RECT 490.460 376.050 490.720 376.370 ;
        RECT 495.060 376.050 495.320 376.370 ;
        RECT 490.520 25.150 490.660 376.050 ;
        RECT 490.460 24.830 490.720 25.150 ;
        RECT 966.100 24.830 966.360 25.150 ;
        RECT 966.160 2.400 966.300 24.830 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 393.830 386.480 394.150 386.540 ;
        RECT 397.050 386.480 397.370 386.540 ;
        RECT 393.830 386.340 397.370 386.480 ;
        RECT 393.830 386.280 394.150 386.340 ;
        RECT 397.050 386.280 397.370 386.340 ;
        RECT 393.830 22.340 394.150 22.400 ;
        RECT 646.830 22.340 647.150 22.400 ;
        RECT 393.830 22.200 647.150 22.340 ;
        RECT 393.830 22.140 394.150 22.200 ;
        RECT 646.830 22.140 647.150 22.200 ;
      LAYER via ;
        RECT 393.860 386.280 394.120 386.540 ;
        RECT 397.080 386.280 397.340 386.540 ;
        RECT 393.860 22.140 394.120 22.400 ;
        RECT 646.860 22.140 647.120 22.400 ;
      LAYER met2 ;
        RECT 398.350 400.250 398.630 404.000 ;
        RECT 397.140 400.110 398.630 400.250 ;
        RECT 397.140 386.570 397.280 400.110 ;
        RECT 398.350 400.000 398.630 400.110 ;
        RECT 393.860 386.250 394.120 386.570 ;
        RECT 397.080 386.250 397.340 386.570 ;
        RECT 393.920 22.430 394.060 386.250 ;
        RECT 393.860 22.110 394.120 22.430 ;
        RECT 646.860 22.110 647.120 22.430 ;
        RECT 646.920 2.400 647.060 22.110 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 496.870 386.480 497.190 386.540 ;
        RECT 500.550 386.480 500.870 386.540 ;
        RECT 496.870 386.340 500.870 386.480 ;
        RECT 496.870 386.280 497.190 386.340 ;
        RECT 500.550 386.280 500.870 386.340 ;
        RECT 496.870 24.720 497.190 24.780 ;
        RECT 984.010 24.720 984.330 24.780 ;
        RECT 496.870 24.580 984.330 24.720 ;
        RECT 496.870 24.520 497.190 24.580 ;
        RECT 984.010 24.520 984.330 24.580 ;
      LAYER via ;
        RECT 496.900 386.280 497.160 386.540 ;
        RECT 500.580 386.280 500.840 386.540 ;
        RECT 496.900 24.520 497.160 24.780 ;
        RECT 984.040 24.520 984.300 24.780 ;
      LAYER met2 ;
        RECT 501.390 400.250 501.670 404.000 ;
        RECT 500.640 400.110 501.670 400.250 ;
        RECT 500.640 386.570 500.780 400.110 ;
        RECT 501.390 400.000 501.670 400.110 ;
        RECT 496.900 386.250 497.160 386.570 ;
        RECT 500.580 386.250 500.840 386.570 ;
        RECT 496.960 24.810 497.100 386.250 ;
        RECT 496.900 24.490 497.160 24.810 ;
        RECT 984.040 24.490 984.300 24.810 ;
        RECT 984.100 2.400 984.240 24.490 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 503.770 386.480 504.090 386.540 ;
        RECT 505.610 386.480 505.930 386.540 ;
        RECT 503.770 386.340 505.930 386.480 ;
        RECT 503.770 386.280 504.090 386.340 ;
        RECT 505.610 386.280 505.930 386.340 ;
        RECT 503.770 24.380 504.090 24.440 ;
        RECT 1001.490 24.380 1001.810 24.440 ;
        RECT 503.770 24.240 1001.810 24.380 ;
        RECT 503.770 24.180 504.090 24.240 ;
        RECT 1001.490 24.180 1001.810 24.240 ;
      LAYER via ;
        RECT 503.800 386.280 504.060 386.540 ;
        RECT 505.640 386.280 505.900 386.540 ;
        RECT 503.800 24.180 504.060 24.440 ;
        RECT 1001.520 24.180 1001.780 24.440 ;
      LAYER met2 ;
        RECT 506.910 400.250 507.190 404.000 ;
        RECT 505.700 400.110 507.190 400.250 ;
        RECT 505.700 386.570 505.840 400.110 ;
        RECT 506.910 400.000 507.190 400.110 ;
        RECT 503.800 386.250 504.060 386.570 ;
        RECT 505.640 386.250 505.900 386.570 ;
        RECT 503.860 24.470 504.000 386.250 ;
        RECT 503.800 24.150 504.060 24.470 ;
        RECT 1001.520 24.150 1001.780 24.470 ;
        RECT 1001.580 2.400 1001.720 24.150 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 510.670 386.480 510.990 386.540 ;
        RECT 511.590 386.480 511.910 386.540 ;
        RECT 510.670 386.340 511.910 386.480 ;
        RECT 510.670 386.280 510.990 386.340 ;
        RECT 511.590 386.280 511.910 386.340 ;
        RECT 510.670 24.040 510.990 24.100 ;
        RECT 1019.430 24.040 1019.750 24.100 ;
        RECT 510.670 23.900 1019.750 24.040 ;
        RECT 510.670 23.840 510.990 23.900 ;
        RECT 1019.430 23.840 1019.750 23.900 ;
      LAYER via ;
        RECT 510.700 386.280 510.960 386.540 ;
        RECT 511.620 386.280 511.880 386.540 ;
        RECT 510.700 23.840 510.960 24.100 ;
        RECT 1019.460 23.840 1019.720 24.100 ;
      LAYER met2 ;
        RECT 512.430 400.250 512.710 404.000 ;
        RECT 511.680 400.110 512.710 400.250 ;
        RECT 511.680 386.570 511.820 400.110 ;
        RECT 512.430 400.000 512.710 400.110 ;
        RECT 510.700 386.250 510.960 386.570 ;
        RECT 511.620 386.250 511.880 386.570 ;
        RECT 510.760 24.130 510.900 386.250 ;
        RECT 510.700 23.810 510.960 24.130 ;
        RECT 1019.460 23.810 1019.720 24.130 ;
        RECT 1019.520 2.400 1019.660 23.810 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.950 400.250 518.230 404.000 ;
        RECT 517.950 400.110 518.720 400.250 ;
        RECT 517.950 400.000 518.230 400.110 ;
        RECT 518.580 25.685 518.720 400.110 ;
        RECT 518.510 25.315 518.790 25.685 ;
        RECT 1036.930 25.315 1037.210 25.685 ;
        RECT 1037.000 2.400 1037.140 25.315 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
      LAYER via2 ;
        RECT 518.510 25.360 518.790 25.640 ;
        RECT 1036.930 25.360 1037.210 25.640 ;
      LAYER met3 ;
        RECT 518.485 25.650 518.815 25.665 ;
        RECT 1036.905 25.650 1037.235 25.665 ;
        RECT 518.485 25.350 1037.235 25.650 ;
        RECT 518.485 25.335 518.815 25.350 ;
        RECT 1036.905 25.335 1037.235 25.350 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.570 386.140 517.890 386.200 ;
        RECT 522.170 386.140 522.490 386.200 ;
        RECT 517.570 386.000 522.490 386.140 ;
        RECT 517.570 385.940 517.890 386.000 ;
        RECT 522.170 385.940 522.490 386.000 ;
      LAYER via ;
        RECT 517.600 385.940 517.860 386.200 ;
        RECT 522.200 385.940 522.460 386.200 ;
      LAYER met2 ;
        RECT 523.470 400.250 523.750 404.000 ;
        RECT 522.260 400.110 523.750 400.250 ;
        RECT 522.260 386.230 522.400 400.110 ;
        RECT 523.470 400.000 523.750 400.110 ;
        RECT 517.600 385.910 517.860 386.230 ;
        RECT 522.200 385.910 522.460 386.230 ;
        RECT 517.660 25.005 517.800 385.910 ;
        RECT 517.590 24.635 517.870 25.005 ;
        RECT 1054.870 24.635 1055.150 25.005 ;
        RECT 1054.940 2.400 1055.080 24.635 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
      LAYER via2 ;
        RECT 517.590 24.680 517.870 24.960 ;
        RECT 1054.870 24.680 1055.150 24.960 ;
      LAYER met3 ;
        RECT 517.565 24.970 517.895 24.985 ;
        RECT 1054.845 24.970 1055.175 24.985 ;
        RECT 517.565 24.670 1055.175 24.970 ;
        RECT 517.565 24.655 517.895 24.670 ;
        RECT 1054.845 24.655 1055.175 24.670 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 529.070 389.880 529.390 389.940 ;
        RECT 776.090 389.880 776.410 389.940 ;
        RECT 529.070 389.740 776.410 389.880 ;
        RECT 529.070 389.680 529.390 389.740 ;
        RECT 776.090 389.680 776.410 389.740 ;
        RECT 776.090 28.800 776.410 28.860 ;
        RECT 1072.330 28.800 1072.650 28.860 ;
        RECT 776.090 28.660 1072.650 28.800 ;
        RECT 776.090 28.600 776.410 28.660 ;
        RECT 1072.330 28.600 1072.650 28.660 ;
      LAYER via ;
        RECT 529.100 389.680 529.360 389.940 ;
        RECT 776.120 389.680 776.380 389.940 ;
        RECT 776.120 28.600 776.380 28.860 ;
        RECT 1072.360 28.600 1072.620 28.860 ;
      LAYER met2 ;
        RECT 528.990 400.180 529.270 404.000 ;
        RECT 528.990 400.000 529.300 400.180 ;
        RECT 529.160 389.970 529.300 400.000 ;
        RECT 529.100 389.650 529.360 389.970 ;
        RECT 776.120 389.650 776.380 389.970 ;
        RECT 776.180 28.890 776.320 389.650 ;
        RECT 776.120 28.570 776.380 28.890 ;
        RECT 1072.360 28.570 1072.620 28.890 ;
        RECT 1072.420 2.400 1072.560 28.570 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 534.130 390.900 534.450 390.960 ;
        RECT 534.130 390.760 545.170 390.900 ;
        RECT 534.130 390.700 534.450 390.760 ;
        RECT 545.030 390.560 545.170 390.760 ;
        RECT 769.190 390.560 769.510 390.620 ;
        RECT 545.030 390.420 769.510 390.560 ;
        RECT 769.190 390.360 769.510 390.420 ;
        RECT 769.190 29.480 769.510 29.540 ;
        RECT 1090.730 29.480 1091.050 29.540 ;
        RECT 769.190 29.340 1091.050 29.480 ;
        RECT 769.190 29.280 769.510 29.340 ;
        RECT 1090.730 29.280 1091.050 29.340 ;
      LAYER via ;
        RECT 534.160 390.700 534.420 390.960 ;
        RECT 769.220 390.360 769.480 390.620 ;
        RECT 769.220 29.280 769.480 29.540 ;
        RECT 1090.760 29.280 1091.020 29.540 ;
      LAYER met2 ;
        RECT 534.050 400.180 534.330 404.000 ;
        RECT 534.050 400.000 534.360 400.180 ;
        RECT 534.220 390.990 534.360 400.000 ;
        RECT 534.160 390.670 534.420 390.990 ;
        RECT 769.220 390.330 769.480 390.650 ;
        RECT 769.280 29.570 769.420 390.330 ;
        RECT 769.220 29.250 769.480 29.570 ;
        RECT 1090.760 29.250 1091.020 29.570 ;
        RECT 1090.820 14.690 1090.960 29.250 ;
        RECT 1090.360 14.550 1090.960 14.690 ;
        RECT 1090.360 2.400 1090.500 14.550 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 539.650 390.220 539.970 390.280 ;
        RECT 782.990 390.220 783.310 390.280 ;
        RECT 539.650 390.080 783.310 390.220 ;
        RECT 539.650 390.020 539.970 390.080 ;
        RECT 782.990 390.020 783.310 390.080 ;
        RECT 782.990 29.140 783.310 29.200 ;
        RECT 1107.750 29.140 1108.070 29.200 ;
        RECT 782.990 29.000 1108.070 29.140 ;
        RECT 782.990 28.940 783.310 29.000 ;
        RECT 1107.750 28.940 1108.070 29.000 ;
      LAYER via ;
        RECT 539.680 390.020 539.940 390.280 ;
        RECT 783.020 390.020 783.280 390.280 ;
        RECT 783.020 28.940 783.280 29.200 ;
        RECT 1107.780 28.940 1108.040 29.200 ;
      LAYER met2 ;
        RECT 539.570 400.180 539.850 404.000 ;
        RECT 539.570 400.000 539.880 400.180 ;
        RECT 539.740 390.310 539.880 400.000 ;
        RECT 539.680 389.990 539.940 390.310 ;
        RECT 783.020 389.990 783.280 390.310 ;
        RECT 783.080 29.230 783.220 389.990 ;
        RECT 783.020 28.910 783.280 29.230 ;
        RECT 1107.780 28.910 1108.040 29.230 ;
        RECT 1107.840 2.400 1107.980 28.910 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.170 31.860 545.490 31.920 ;
        RECT 1125.690 31.860 1126.010 31.920 ;
        RECT 545.170 31.720 1126.010 31.860 ;
        RECT 545.170 31.660 545.490 31.720 ;
        RECT 1125.690 31.660 1126.010 31.720 ;
      LAYER via ;
        RECT 545.200 31.660 545.460 31.920 ;
        RECT 1125.720 31.660 1125.980 31.920 ;
      LAYER met2 ;
        RECT 545.090 400.180 545.370 404.000 ;
        RECT 545.090 400.000 545.400 400.180 ;
        RECT 545.260 31.950 545.400 400.000 ;
        RECT 545.200 31.630 545.460 31.950 ;
        RECT 1125.720 31.630 1125.980 31.950 ;
        RECT 1125.780 2.400 1125.920 31.630 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 545.630 375.940 545.950 376.000 ;
        RECT 549.310 375.940 549.630 376.000 ;
        RECT 545.630 375.800 549.630 375.940 ;
        RECT 545.630 375.740 545.950 375.800 ;
        RECT 549.310 375.740 549.630 375.800 ;
        RECT 545.630 29.820 545.950 29.880 ;
        RECT 1143.630 29.820 1143.950 29.880 ;
        RECT 545.630 29.680 1143.950 29.820 ;
        RECT 545.630 29.620 545.950 29.680 ;
        RECT 1143.630 29.620 1143.950 29.680 ;
      LAYER via ;
        RECT 545.660 375.740 545.920 376.000 ;
        RECT 549.340 375.740 549.600 376.000 ;
        RECT 545.660 29.620 545.920 29.880 ;
        RECT 1143.660 29.620 1143.920 29.880 ;
      LAYER met2 ;
        RECT 550.610 400.250 550.890 404.000 ;
        RECT 549.400 400.110 550.890 400.250 ;
        RECT 549.400 376.030 549.540 400.110 ;
        RECT 550.610 400.000 550.890 400.110 ;
        RECT 545.660 375.710 545.920 376.030 ;
        RECT 549.340 375.710 549.600 376.030 ;
        RECT 545.720 29.910 545.860 375.710 ;
        RECT 545.660 29.590 545.920 29.910 ;
        RECT 1143.660 29.590 1143.920 29.910 ;
        RECT 1143.720 2.400 1143.860 29.590 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.270 387.160 400.590 387.220 ;
        RECT 402.110 387.160 402.430 387.220 ;
        RECT 400.270 387.020 402.430 387.160 ;
        RECT 400.270 386.960 400.590 387.020 ;
        RECT 402.110 386.960 402.430 387.020 ;
        RECT 400.270 23.020 400.590 23.080 ;
        RECT 664.770 23.020 665.090 23.080 ;
        RECT 400.270 22.880 665.090 23.020 ;
        RECT 400.270 22.820 400.590 22.880 ;
        RECT 664.770 22.820 665.090 22.880 ;
      LAYER via ;
        RECT 400.300 386.960 400.560 387.220 ;
        RECT 402.140 386.960 402.400 387.220 ;
        RECT 400.300 22.820 400.560 23.080 ;
        RECT 664.800 22.820 665.060 23.080 ;
      LAYER met2 ;
        RECT 403.410 400.250 403.690 404.000 ;
        RECT 402.200 400.110 403.690 400.250 ;
        RECT 402.200 387.250 402.340 400.110 ;
        RECT 403.410 400.000 403.690 400.110 ;
        RECT 400.300 386.930 400.560 387.250 ;
        RECT 402.140 386.930 402.400 387.250 ;
        RECT 400.360 23.110 400.500 386.930 ;
        RECT 400.300 22.790 400.560 23.110 ;
        RECT 664.800 22.790 665.060 23.110 ;
        RECT 664.860 2.400 665.000 22.790 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.070 375.940 552.390 376.000 ;
        RECT 554.830 375.940 555.150 376.000 ;
        RECT 552.070 375.800 555.150 375.940 ;
        RECT 552.070 375.740 552.390 375.800 ;
        RECT 554.830 375.740 555.150 375.800 ;
        RECT 552.070 30.160 552.390 30.220 ;
        RECT 1161.110 30.160 1161.430 30.220 ;
        RECT 552.070 30.020 1161.430 30.160 ;
        RECT 552.070 29.960 552.390 30.020 ;
        RECT 1161.110 29.960 1161.430 30.020 ;
      LAYER via ;
        RECT 552.100 375.740 552.360 376.000 ;
        RECT 554.860 375.740 555.120 376.000 ;
        RECT 552.100 29.960 552.360 30.220 ;
        RECT 1161.140 29.960 1161.400 30.220 ;
      LAYER met2 ;
        RECT 556.130 400.250 556.410 404.000 ;
        RECT 554.920 400.110 556.410 400.250 ;
        RECT 554.920 376.030 555.060 400.110 ;
        RECT 556.130 400.000 556.410 400.110 ;
        RECT 552.100 375.710 552.360 376.030 ;
        RECT 554.860 375.710 555.120 376.030 ;
        RECT 552.160 30.250 552.300 375.710 ;
        RECT 552.100 29.930 552.360 30.250 ;
        RECT 1161.140 29.930 1161.400 30.250 ;
        RECT 1161.200 2.400 1161.340 29.930 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 558.970 393.960 559.290 394.020 ;
        RECT 561.730 393.960 562.050 394.020 ;
        RECT 558.970 393.820 562.050 393.960 ;
        RECT 558.970 393.760 559.290 393.820 ;
        RECT 561.730 393.760 562.050 393.820 ;
        RECT 558.970 30.500 559.290 30.560 ;
        RECT 1179.050 30.500 1179.370 30.560 ;
        RECT 558.970 30.360 1179.370 30.500 ;
        RECT 558.970 30.300 559.290 30.360 ;
        RECT 1179.050 30.300 1179.370 30.360 ;
      LAYER via ;
        RECT 559.000 393.760 559.260 394.020 ;
        RECT 561.760 393.760 562.020 394.020 ;
        RECT 559.000 30.300 559.260 30.560 ;
        RECT 1179.080 30.300 1179.340 30.560 ;
      LAYER met2 ;
        RECT 561.650 400.180 561.930 404.000 ;
        RECT 561.650 400.000 561.960 400.180 ;
        RECT 561.820 394.050 561.960 400.000 ;
        RECT 559.000 393.730 559.260 394.050 ;
        RECT 561.760 393.730 562.020 394.050 ;
        RECT 559.060 30.590 559.200 393.730 ;
        RECT 559.000 30.270 559.260 30.590 ;
        RECT 1179.080 30.270 1179.340 30.590 ;
        RECT 1179.140 2.400 1179.280 30.270 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 565.870 34.240 566.190 34.300 ;
        RECT 1196.530 34.240 1196.850 34.300 ;
        RECT 565.870 34.100 1196.850 34.240 ;
        RECT 565.870 34.040 566.190 34.100 ;
        RECT 1196.530 34.040 1196.850 34.100 ;
      LAYER via ;
        RECT 565.900 34.040 566.160 34.300 ;
        RECT 1196.560 34.040 1196.820 34.300 ;
      LAYER met2 ;
        RECT 567.170 400.250 567.450 404.000 ;
        RECT 565.960 400.110 567.450 400.250 ;
        RECT 565.960 34.330 566.100 400.110 ;
        RECT 567.170 400.000 567.450 400.110 ;
        RECT 565.900 34.010 566.160 34.330 ;
        RECT 1196.560 34.010 1196.820 34.330 ;
        RECT 1196.620 2.400 1196.760 34.010 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.330 376.280 566.650 376.340 ;
        RECT 570.930 376.280 571.250 376.340 ;
        RECT 566.330 376.140 571.250 376.280 ;
        RECT 566.330 376.080 566.650 376.140 ;
        RECT 570.930 376.080 571.250 376.140 ;
        RECT 566.330 33.900 566.650 33.960 ;
        RECT 1214.930 33.900 1215.250 33.960 ;
        RECT 566.330 33.760 1215.250 33.900 ;
        RECT 566.330 33.700 566.650 33.760 ;
        RECT 1214.930 33.700 1215.250 33.760 ;
      LAYER via ;
        RECT 566.360 376.080 566.620 376.340 ;
        RECT 570.960 376.080 571.220 376.340 ;
        RECT 566.360 33.700 566.620 33.960 ;
        RECT 1214.960 33.700 1215.220 33.960 ;
      LAYER met2 ;
        RECT 572.230 400.250 572.510 404.000 ;
        RECT 571.020 400.110 572.510 400.250 ;
        RECT 571.020 376.370 571.160 400.110 ;
        RECT 572.230 400.000 572.510 400.110 ;
        RECT 566.360 376.050 566.620 376.370 ;
        RECT 570.960 376.050 571.220 376.370 ;
        RECT 566.420 33.990 566.560 376.050 ;
        RECT 566.360 33.670 566.620 33.990 ;
        RECT 1214.960 33.670 1215.220 33.990 ;
        RECT 1215.020 14.690 1215.160 33.670 ;
        RECT 1214.560 14.550 1215.160 14.690 ;
        RECT 1214.560 2.400 1214.700 14.550 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 572.770 376.280 573.090 376.340 ;
        RECT 576.450 376.280 576.770 376.340 ;
        RECT 572.770 376.140 576.770 376.280 ;
        RECT 572.770 376.080 573.090 376.140 ;
        RECT 576.450 376.080 576.770 376.140 ;
        RECT 572.770 33.560 573.090 33.620 ;
        RECT 1231.950 33.560 1232.270 33.620 ;
        RECT 572.770 33.420 1232.270 33.560 ;
        RECT 572.770 33.360 573.090 33.420 ;
        RECT 1231.950 33.360 1232.270 33.420 ;
      LAYER via ;
        RECT 572.800 376.080 573.060 376.340 ;
        RECT 576.480 376.080 576.740 376.340 ;
        RECT 572.800 33.360 573.060 33.620 ;
        RECT 1231.980 33.360 1232.240 33.620 ;
      LAYER met2 ;
        RECT 577.750 400.250 578.030 404.000 ;
        RECT 576.540 400.110 578.030 400.250 ;
        RECT 576.540 376.370 576.680 400.110 ;
        RECT 577.750 400.000 578.030 400.110 ;
        RECT 572.800 376.050 573.060 376.370 ;
        RECT 576.480 376.050 576.740 376.370 ;
        RECT 572.860 33.650 573.000 376.050 ;
        RECT 572.800 33.330 573.060 33.650 ;
        RECT 1231.980 33.330 1232.240 33.650 ;
        RECT 1232.040 2.400 1232.180 33.330 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 579.670 375.940 579.990 376.000 ;
        RECT 581.970 375.940 582.290 376.000 ;
        RECT 579.670 375.800 582.290 375.940 ;
        RECT 579.670 375.740 579.990 375.800 ;
        RECT 581.970 375.740 582.290 375.800 ;
        RECT 579.670 33.220 579.990 33.280 ;
        RECT 1249.890 33.220 1250.210 33.280 ;
        RECT 579.670 33.080 1250.210 33.220 ;
        RECT 579.670 33.020 579.990 33.080 ;
        RECT 1249.890 33.020 1250.210 33.080 ;
      LAYER via ;
        RECT 579.700 375.740 579.960 376.000 ;
        RECT 582.000 375.740 582.260 376.000 ;
        RECT 579.700 33.020 579.960 33.280 ;
        RECT 1249.920 33.020 1250.180 33.280 ;
      LAYER met2 ;
        RECT 583.270 400.250 583.550 404.000 ;
        RECT 582.060 400.110 583.550 400.250 ;
        RECT 582.060 376.030 582.200 400.110 ;
        RECT 583.270 400.000 583.550 400.110 ;
        RECT 579.700 375.710 579.960 376.030 ;
        RECT 582.000 375.710 582.260 376.030 ;
        RECT 579.760 33.310 579.900 375.710 ;
        RECT 579.700 32.990 579.960 33.310 ;
        RECT 1249.920 32.990 1250.180 33.310 ;
        RECT 1249.980 2.400 1250.120 32.990 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 586.570 381.720 586.890 381.780 ;
        RECT 588.870 381.720 589.190 381.780 ;
        RECT 586.570 381.580 589.190 381.720 ;
        RECT 586.570 381.520 586.890 381.580 ;
        RECT 588.870 381.520 589.190 381.580 ;
        RECT 586.570 32.880 586.890 32.940 ;
        RECT 1267.370 32.880 1267.690 32.940 ;
        RECT 586.570 32.740 1267.690 32.880 ;
        RECT 586.570 32.680 586.890 32.740 ;
        RECT 1267.370 32.680 1267.690 32.740 ;
      LAYER via ;
        RECT 586.600 381.520 586.860 381.780 ;
        RECT 588.900 381.520 589.160 381.780 ;
        RECT 586.600 32.680 586.860 32.940 ;
        RECT 1267.400 32.680 1267.660 32.940 ;
      LAYER met2 ;
        RECT 588.790 400.180 589.070 404.000 ;
        RECT 588.790 400.000 589.100 400.180 ;
        RECT 588.960 381.810 589.100 400.000 ;
        RECT 586.600 381.490 586.860 381.810 ;
        RECT 588.900 381.490 589.160 381.810 ;
        RECT 586.660 32.970 586.800 381.490 ;
        RECT 586.600 32.650 586.860 32.970 ;
        RECT 1267.400 32.650 1267.660 32.970 ;
        RECT 1267.460 2.400 1267.600 32.650 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.930 32.540 594.250 32.600 ;
        RECT 1285.310 32.540 1285.630 32.600 ;
        RECT 593.930 32.400 1285.630 32.540 ;
        RECT 593.930 32.340 594.250 32.400 ;
        RECT 1285.310 32.340 1285.630 32.400 ;
      LAYER via ;
        RECT 593.960 32.340 594.220 32.600 ;
        RECT 1285.340 32.340 1285.600 32.600 ;
      LAYER met2 ;
        RECT 594.310 400.250 594.590 404.000 ;
        RECT 594.020 400.110 594.590 400.250 ;
        RECT 594.020 32.630 594.160 400.110 ;
        RECT 594.310 400.000 594.590 400.110 ;
        RECT 593.960 32.310 594.220 32.630 ;
        RECT 1285.340 32.310 1285.600 32.630 ;
        RECT 1285.400 2.400 1285.540 32.310 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 593.470 376.280 593.790 376.340 ;
        RECT 598.530 376.280 598.850 376.340 ;
        RECT 593.470 376.140 598.850 376.280 ;
        RECT 593.470 376.080 593.790 376.140 ;
        RECT 598.530 376.080 598.850 376.140 ;
      LAYER via ;
        RECT 593.500 376.080 593.760 376.340 ;
        RECT 598.560 376.080 598.820 376.340 ;
      LAYER met2 ;
        RECT 599.830 400.250 600.110 404.000 ;
        RECT 598.620 400.110 600.110 400.250 ;
        RECT 598.620 376.370 598.760 400.110 ;
        RECT 599.830 400.000 600.110 400.110 ;
        RECT 593.500 376.050 593.760 376.370 ;
        RECT 598.560 376.050 598.820 376.370 ;
        RECT 593.560 31.805 593.700 376.050 ;
        RECT 593.490 31.435 593.770 31.805 ;
        RECT 1303.270 31.435 1303.550 31.805 ;
        RECT 1303.340 2.400 1303.480 31.435 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
      LAYER via2 ;
        RECT 593.490 31.480 593.770 31.760 ;
        RECT 1303.270 31.480 1303.550 31.760 ;
      LAYER met3 ;
        RECT 593.465 31.770 593.795 31.785 ;
        RECT 1303.245 31.770 1303.575 31.785 ;
        RECT 593.465 31.470 1303.575 31.770 ;
        RECT 593.465 31.455 593.795 31.470 ;
        RECT 1303.245 31.455 1303.575 31.470 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.370 375.940 600.690 376.000 ;
        RECT 603.590 375.940 603.910 376.000 ;
        RECT 600.370 375.800 603.910 375.940 ;
        RECT 600.370 375.740 600.690 375.800 ;
        RECT 603.590 375.740 603.910 375.800 ;
      LAYER via ;
        RECT 600.400 375.740 600.660 376.000 ;
        RECT 603.620 375.740 603.880 376.000 ;
      LAYER met2 ;
        RECT 604.890 400.250 605.170 404.000 ;
        RECT 603.680 400.110 605.170 400.250 ;
        RECT 603.680 376.030 603.820 400.110 ;
        RECT 604.890 400.000 605.170 400.110 ;
        RECT 600.400 375.710 600.660 376.030 ;
        RECT 603.620 375.710 603.880 376.030 ;
        RECT 600.460 31.125 600.600 375.710 ;
        RECT 600.390 30.755 600.670 31.125 ;
        RECT 1320.750 30.755 1321.030 31.125 ;
        RECT 1320.820 2.400 1320.960 30.755 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
      LAYER via2 ;
        RECT 600.390 30.800 600.670 31.080 ;
        RECT 1320.750 30.800 1321.030 31.080 ;
      LAYER met3 ;
        RECT 600.365 31.090 600.695 31.105 ;
        RECT 1320.725 31.090 1321.055 31.105 ;
        RECT 600.365 30.790 1321.055 31.090 ;
        RECT 600.365 30.775 600.695 30.790 ;
        RECT 1320.725 30.775 1321.055 30.790 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.170 386.480 407.490 386.540 ;
        RECT 408.550 386.480 408.870 386.540 ;
        RECT 407.170 386.340 408.870 386.480 ;
        RECT 407.170 386.280 407.490 386.340 ;
        RECT 408.550 386.280 408.870 386.340 ;
        RECT 407.170 23.360 407.490 23.420 ;
        RECT 682.250 23.360 682.570 23.420 ;
        RECT 407.170 23.220 682.570 23.360 ;
        RECT 407.170 23.160 407.490 23.220 ;
        RECT 682.250 23.160 682.570 23.220 ;
      LAYER via ;
        RECT 407.200 386.280 407.460 386.540 ;
        RECT 408.580 386.280 408.840 386.540 ;
        RECT 407.200 23.160 407.460 23.420 ;
        RECT 682.280 23.160 682.540 23.420 ;
      LAYER met2 ;
        RECT 408.930 400.250 409.210 404.000 ;
        RECT 408.640 400.110 409.210 400.250 ;
        RECT 408.640 386.570 408.780 400.110 ;
        RECT 408.930 400.000 409.210 400.110 ;
        RECT 407.200 386.250 407.460 386.570 ;
        RECT 408.580 386.250 408.840 386.570 ;
        RECT 407.260 23.450 407.400 386.250 ;
        RECT 407.200 23.130 407.460 23.450 ;
        RECT 682.280 23.130 682.540 23.450 ;
        RECT 682.340 2.400 682.480 23.130 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 608.190 105.640 608.510 105.700 ;
        RECT 1338.670 105.640 1338.990 105.700 ;
        RECT 608.190 105.500 1338.990 105.640 ;
        RECT 608.190 105.440 608.510 105.500 ;
        RECT 1338.670 105.440 1338.990 105.500 ;
      LAYER via ;
        RECT 608.220 105.440 608.480 105.700 ;
        RECT 1338.700 105.440 1338.960 105.700 ;
      LAYER met2 ;
        RECT 610.410 400.250 610.690 404.000 ;
        RECT 609.200 400.110 610.690 400.250 ;
        RECT 609.200 324.370 609.340 400.110 ;
        RECT 610.410 400.000 610.690 400.110 ;
        RECT 608.280 324.230 609.340 324.370 ;
        RECT 608.280 105.730 608.420 324.230 ;
        RECT 608.220 105.410 608.480 105.730 ;
        RECT 1338.700 105.410 1338.960 105.730 ;
        RECT 1338.760 2.400 1338.900 105.410 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.550 105.980 615.870 106.040 ;
        RECT 1352.470 105.980 1352.790 106.040 ;
        RECT 615.550 105.840 1352.790 105.980 ;
        RECT 615.550 105.780 615.870 105.840 ;
        RECT 1352.470 105.780 1352.790 105.840 ;
      LAYER via ;
        RECT 615.580 105.780 615.840 106.040 ;
        RECT 1352.500 105.780 1352.760 106.040 ;
      LAYER met2 ;
        RECT 615.930 400.250 616.210 404.000 ;
        RECT 615.640 400.110 616.210 400.250 ;
        RECT 615.640 106.070 615.780 400.110 ;
        RECT 615.930 400.000 616.210 400.110 ;
        RECT 615.580 105.750 615.840 106.070 ;
        RECT 1352.500 105.750 1352.760 106.070 ;
        RECT 1352.560 82.870 1352.700 105.750 ;
        RECT 1352.560 82.730 1354.080 82.870 ;
        RECT 1353.940 1.770 1354.080 82.730 ;
        RECT 1356.030 1.770 1356.590 2.400 ;
        RECT 1353.940 1.630 1356.590 1.770 ;
        RECT 1356.030 -4.800 1356.590 1.630 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.990 106.320 622.310 106.380 ;
        RECT 1373.170 106.320 1373.490 106.380 ;
        RECT 621.990 106.180 1373.490 106.320 ;
        RECT 621.990 106.120 622.310 106.180 ;
        RECT 1373.170 106.120 1373.490 106.180 ;
      LAYER via ;
        RECT 622.020 106.120 622.280 106.380 ;
        RECT 1373.200 106.120 1373.460 106.380 ;
      LAYER met2 ;
        RECT 621.450 400.250 621.730 404.000 ;
        RECT 621.450 400.110 622.220 400.250 ;
        RECT 621.450 400.000 621.730 400.110 ;
        RECT 622.080 106.410 622.220 400.110 ;
        RECT 622.020 106.090 622.280 106.410 ;
        RECT 1373.200 106.090 1373.460 106.410 ;
        RECT 1373.260 82.870 1373.400 106.090 ;
        RECT 1373.260 82.730 1374.320 82.870 ;
        RECT 1374.180 2.400 1374.320 82.730 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 622.450 106.660 622.770 106.720 ;
        RECT 1386.970 106.660 1387.290 106.720 ;
        RECT 622.450 106.520 1387.290 106.660 ;
        RECT 622.450 106.460 622.770 106.520 ;
        RECT 1386.970 106.460 1387.290 106.520 ;
      LAYER via ;
        RECT 622.480 106.460 622.740 106.720 ;
        RECT 1387.000 106.460 1387.260 106.720 ;
      LAYER met2 ;
        RECT 626.970 400.250 627.250 404.000 ;
        RECT 625.760 400.110 627.250 400.250 ;
        RECT 625.760 324.370 625.900 400.110 ;
        RECT 626.970 400.000 627.250 400.110 ;
        RECT 622.540 324.230 625.900 324.370 ;
        RECT 622.540 106.750 622.680 324.230 ;
        RECT 622.480 106.430 622.740 106.750 ;
        RECT 1387.000 106.430 1387.260 106.750 ;
        RECT 1387.060 82.870 1387.200 106.430 ;
        RECT 1387.060 82.730 1391.800 82.870 ;
        RECT 1391.660 2.400 1391.800 82.730 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 629.350 110.400 629.670 110.460 ;
        RECT 1407.670 110.400 1407.990 110.460 ;
        RECT 629.350 110.260 1407.990 110.400 ;
        RECT 629.350 110.200 629.670 110.260 ;
        RECT 1407.670 110.200 1407.990 110.260 ;
      LAYER via ;
        RECT 629.380 110.200 629.640 110.460 ;
        RECT 1407.700 110.200 1407.960 110.460 ;
      LAYER met2 ;
        RECT 632.490 400.250 632.770 404.000 ;
        RECT 631.280 400.110 632.770 400.250 ;
        RECT 631.280 324.370 631.420 400.110 ;
        RECT 632.490 400.000 632.770 400.110 ;
        RECT 629.440 324.230 631.420 324.370 ;
        RECT 629.440 110.490 629.580 324.230 ;
        RECT 629.380 110.170 629.640 110.490 ;
        RECT 1407.700 110.170 1407.960 110.490 ;
        RECT 1407.760 1.770 1407.900 110.170 ;
        RECT 1409.390 1.770 1409.950 2.400 ;
        RECT 1407.760 1.630 1409.950 1.770 ;
        RECT 1409.390 -4.800 1409.950 1.630 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 634.870 399.740 635.190 399.800 ;
        RECT 636.250 399.740 636.570 399.800 ;
        RECT 634.870 399.600 636.570 399.740 ;
        RECT 634.870 399.540 635.190 399.600 ;
        RECT 636.250 399.540 636.570 399.600 ;
        RECT 634.870 36.280 635.190 36.340 ;
        RECT 1426.990 36.280 1427.310 36.340 ;
        RECT 634.870 36.140 1427.310 36.280 ;
        RECT 634.870 36.080 635.190 36.140 ;
        RECT 1426.990 36.080 1427.310 36.140 ;
      LAYER via ;
        RECT 634.900 399.540 635.160 399.800 ;
        RECT 636.280 399.540 636.540 399.800 ;
        RECT 634.900 36.080 635.160 36.340 ;
        RECT 1427.020 36.080 1427.280 36.340 ;
      LAYER met2 ;
        RECT 637.550 400.250 637.830 404.000 ;
        RECT 636.340 400.110 637.830 400.250 ;
        RECT 636.340 399.830 636.480 400.110 ;
        RECT 637.550 400.000 637.830 400.110 ;
        RECT 634.900 399.510 635.160 399.830 ;
        RECT 636.280 399.510 636.540 399.830 ;
        RECT 634.960 36.370 635.100 399.510 ;
        RECT 634.900 36.050 635.160 36.370 ;
        RECT 1427.020 36.050 1427.280 36.370 ;
        RECT 1427.080 2.400 1427.220 36.050 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 641.770 36.620 642.090 36.680 ;
        RECT 1444.930 36.620 1445.250 36.680 ;
        RECT 641.770 36.480 1445.250 36.620 ;
        RECT 641.770 36.420 642.090 36.480 ;
        RECT 1444.930 36.420 1445.250 36.480 ;
      LAYER via ;
        RECT 641.800 36.420 642.060 36.680 ;
        RECT 1444.960 36.420 1445.220 36.680 ;
      LAYER met2 ;
        RECT 643.070 400.250 643.350 404.000 ;
        RECT 641.860 400.110 643.350 400.250 ;
        RECT 641.860 36.710 642.000 400.110 ;
        RECT 643.070 400.000 643.350 400.110 ;
        RECT 641.800 36.390 642.060 36.710 ;
        RECT 1444.960 36.390 1445.220 36.710 ;
        RECT 1445.020 2.400 1445.160 36.390 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 649.130 36.960 649.450 37.020 ;
        RECT 1462.870 36.960 1463.190 37.020 ;
        RECT 649.130 36.820 1463.190 36.960 ;
        RECT 649.130 36.760 649.450 36.820 ;
        RECT 1462.870 36.760 1463.190 36.820 ;
      LAYER via ;
        RECT 649.160 36.760 649.420 37.020 ;
        RECT 1462.900 36.760 1463.160 37.020 ;
      LAYER met2 ;
        RECT 648.590 400.250 648.870 404.000 ;
        RECT 648.590 400.110 649.360 400.250 ;
        RECT 648.590 400.000 648.870 400.110 ;
        RECT 649.220 37.050 649.360 400.110 ;
        RECT 649.160 36.730 649.420 37.050 ;
        RECT 1462.900 36.730 1463.160 37.050 ;
        RECT 1462.960 2.400 1463.100 36.730 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 648.670 386.480 648.990 386.540 ;
        RECT 652.810 386.480 653.130 386.540 ;
        RECT 648.670 386.340 653.130 386.480 ;
        RECT 648.670 386.280 648.990 386.340 ;
        RECT 652.810 386.280 653.130 386.340 ;
        RECT 648.670 37.300 648.990 37.360 ;
        RECT 1480.350 37.300 1480.670 37.360 ;
        RECT 648.670 37.160 1480.670 37.300 ;
        RECT 648.670 37.100 648.990 37.160 ;
        RECT 1480.350 37.100 1480.670 37.160 ;
      LAYER via ;
        RECT 648.700 386.280 648.960 386.540 ;
        RECT 652.840 386.280 653.100 386.540 ;
        RECT 648.700 37.100 648.960 37.360 ;
        RECT 1480.380 37.100 1480.640 37.360 ;
      LAYER met2 ;
        RECT 654.110 400.250 654.390 404.000 ;
        RECT 652.900 400.110 654.390 400.250 ;
        RECT 652.900 386.570 653.040 400.110 ;
        RECT 654.110 400.000 654.390 400.110 ;
        RECT 648.700 386.250 648.960 386.570 ;
        RECT 652.840 386.250 653.100 386.570 ;
        RECT 648.760 37.390 648.900 386.250 ;
        RECT 648.700 37.070 648.960 37.390 ;
        RECT 1480.380 37.070 1480.640 37.390 ;
        RECT 1480.440 2.400 1480.580 37.070 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 655.570 375.940 655.890 376.000 ;
        RECT 658.330 375.940 658.650 376.000 ;
        RECT 655.570 375.800 658.650 375.940 ;
        RECT 655.570 375.740 655.890 375.800 ;
        RECT 658.330 375.740 658.650 375.800 ;
        RECT 655.570 37.640 655.890 37.700 ;
        RECT 1498.290 37.640 1498.610 37.700 ;
        RECT 655.570 37.500 1498.610 37.640 ;
        RECT 655.570 37.440 655.890 37.500 ;
        RECT 1498.290 37.440 1498.610 37.500 ;
      LAYER via ;
        RECT 655.600 375.740 655.860 376.000 ;
        RECT 658.360 375.740 658.620 376.000 ;
        RECT 655.600 37.440 655.860 37.700 ;
        RECT 1498.320 37.440 1498.580 37.700 ;
      LAYER met2 ;
        RECT 659.630 400.250 659.910 404.000 ;
        RECT 658.420 400.110 659.910 400.250 ;
        RECT 658.420 376.030 658.560 400.110 ;
        RECT 659.630 400.000 659.910 400.110 ;
        RECT 655.600 375.710 655.860 376.030 ;
        RECT 658.360 375.710 658.620 376.030 ;
        RECT 655.660 37.730 655.800 375.710 ;
        RECT 655.600 37.410 655.860 37.730 ;
        RECT 1498.320 37.410 1498.580 37.730 ;
        RECT 1498.380 2.400 1498.520 37.410 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.530 23.700 414.850 23.760 ;
        RECT 700.190 23.700 700.510 23.760 ;
        RECT 414.530 23.560 700.510 23.700 ;
        RECT 414.530 23.500 414.850 23.560 ;
        RECT 700.190 23.500 700.510 23.560 ;
      LAYER via ;
        RECT 414.560 23.500 414.820 23.760 ;
        RECT 700.220 23.500 700.480 23.760 ;
      LAYER met2 ;
        RECT 414.450 400.180 414.730 404.000 ;
        RECT 414.450 400.000 414.760 400.180 ;
        RECT 414.620 23.790 414.760 400.000 ;
        RECT 414.560 23.470 414.820 23.790 ;
        RECT 700.220 23.470 700.480 23.790 ;
        RECT 700.280 2.400 700.420 23.470 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.470 41.380 662.790 41.440 ;
        RECT 1515.770 41.380 1516.090 41.440 ;
        RECT 662.470 41.240 1516.090 41.380 ;
        RECT 662.470 41.180 662.790 41.240 ;
        RECT 1515.770 41.180 1516.090 41.240 ;
      LAYER via ;
        RECT 662.500 41.180 662.760 41.440 ;
        RECT 1515.800 41.180 1516.060 41.440 ;
      LAYER met2 ;
        RECT 665.150 400.250 665.430 404.000 ;
        RECT 663.940 400.110 665.430 400.250 ;
        RECT 663.940 387.330 664.080 400.110 ;
        RECT 665.150 400.000 665.430 400.110 ;
        RECT 662.560 387.190 664.080 387.330 ;
        RECT 662.560 41.470 662.700 387.190 ;
        RECT 662.500 41.150 662.760 41.470 ;
        RECT 1515.800 41.150 1516.060 41.470 ;
        RECT 1515.860 2.400 1516.000 41.150 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.370 41.040 669.690 41.100 ;
        RECT 1533.710 41.040 1534.030 41.100 ;
        RECT 669.370 40.900 1534.030 41.040 ;
        RECT 669.370 40.840 669.690 40.900 ;
        RECT 1533.710 40.840 1534.030 40.900 ;
      LAYER via ;
        RECT 669.400 40.840 669.660 41.100 ;
        RECT 1533.740 40.840 1534.000 41.100 ;
      LAYER met2 ;
        RECT 670.210 400.250 670.490 404.000 ;
        RECT 669.460 400.110 670.490 400.250 ;
        RECT 669.460 41.130 669.600 400.110 ;
        RECT 670.210 400.000 670.490 400.110 ;
        RECT 669.400 40.810 669.660 41.130 ;
        RECT 1533.740 40.810 1534.000 41.130 ;
        RECT 1533.800 2.400 1533.940 40.810 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 669.830 386.140 670.150 386.200 ;
        RECT 674.430 386.140 674.750 386.200 ;
        RECT 669.830 386.000 674.750 386.140 ;
        RECT 669.830 385.940 670.150 386.000 ;
        RECT 674.430 385.940 674.750 386.000 ;
        RECT 669.830 40.700 670.150 40.760 ;
        RECT 1551.190 40.700 1551.510 40.760 ;
        RECT 669.830 40.560 1551.510 40.700 ;
        RECT 669.830 40.500 670.150 40.560 ;
        RECT 1551.190 40.500 1551.510 40.560 ;
      LAYER via ;
        RECT 669.860 385.940 670.120 386.200 ;
        RECT 674.460 385.940 674.720 386.200 ;
        RECT 669.860 40.500 670.120 40.760 ;
        RECT 1551.220 40.500 1551.480 40.760 ;
      LAYER met2 ;
        RECT 675.730 400.250 676.010 404.000 ;
        RECT 674.520 400.110 676.010 400.250 ;
        RECT 674.520 386.230 674.660 400.110 ;
        RECT 675.730 400.000 676.010 400.110 ;
        RECT 669.860 385.910 670.120 386.230 ;
        RECT 674.460 385.910 674.720 386.230 ;
        RECT 669.920 40.790 670.060 385.910 ;
        RECT 669.860 40.470 670.120 40.790 ;
        RECT 1551.220 40.470 1551.480 40.790 ;
        RECT 1551.280 2.400 1551.420 40.470 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.270 373.560 676.590 373.620 ;
        RECT 679.950 373.560 680.270 373.620 ;
        RECT 676.270 373.420 680.270 373.560 ;
        RECT 676.270 373.360 676.590 373.420 ;
        RECT 679.950 373.360 680.270 373.420 ;
        RECT 676.270 40.360 676.590 40.420 ;
        RECT 1569.130 40.360 1569.450 40.420 ;
        RECT 676.270 40.220 1569.450 40.360 ;
        RECT 676.270 40.160 676.590 40.220 ;
        RECT 1569.130 40.160 1569.450 40.220 ;
      LAYER via ;
        RECT 676.300 373.360 676.560 373.620 ;
        RECT 679.980 373.360 680.240 373.620 ;
        RECT 676.300 40.160 676.560 40.420 ;
        RECT 1569.160 40.160 1569.420 40.420 ;
      LAYER met2 ;
        RECT 681.250 400.250 681.530 404.000 ;
        RECT 680.040 400.110 681.530 400.250 ;
        RECT 680.040 373.650 680.180 400.110 ;
        RECT 681.250 400.000 681.530 400.110 ;
        RECT 676.300 373.330 676.560 373.650 ;
        RECT 679.980 373.330 680.240 373.650 ;
        RECT 676.360 40.450 676.500 373.330 ;
        RECT 676.300 40.130 676.560 40.450 ;
        RECT 1569.160 40.130 1569.420 40.450 ;
        RECT 1569.220 2.400 1569.360 40.130 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.170 386.140 683.490 386.200 ;
        RECT 685.470 386.140 685.790 386.200 ;
        RECT 683.170 386.000 685.790 386.140 ;
        RECT 683.170 385.940 683.490 386.000 ;
        RECT 685.470 385.940 685.790 386.000 ;
        RECT 683.170 40.020 683.490 40.080 ;
        RECT 1586.610 40.020 1586.930 40.080 ;
        RECT 683.170 39.880 1586.930 40.020 ;
        RECT 683.170 39.820 683.490 39.880 ;
        RECT 1586.610 39.820 1586.930 39.880 ;
      LAYER via ;
        RECT 683.200 385.940 683.460 386.200 ;
        RECT 685.500 385.940 685.760 386.200 ;
        RECT 683.200 39.820 683.460 40.080 ;
        RECT 1586.640 39.820 1586.900 40.080 ;
      LAYER met2 ;
        RECT 686.770 400.250 687.050 404.000 ;
        RECT 685.560 400.110 687.050 400.250 ;
        RECT 685.560 386.230 685.700 400.110 ;
        RECT 686.770 400.000 687.050 400.110 ;
        RECT 683.200 385.910 683.460 386.230 ;
        RECT 685.500 385.910 685.760 386.230 ;
        RECT 683.260 40.110 683.400 385.910 ;
        RECT 683.200 39.790 683.460 40.110 ;
        RECT 1586.640 39.790 1586.900 40.110 ;
        RECT 1586.700 2.400 1586.840 39.790 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.070 386.480 690.390 386.540 ;
        RECT 691.910 386.480 692.230 386.540 ;
        RECT 690.070 386.340 692.230 386.480 ;
        RECT 690.070 386.280 690.390 386.340 ;
        RECT 691.910 386.280 692.230 386.340 ;
        RECT 690.070 39.680 690.390 39.740 ;
        RECT 1604.550 39.680 1604.870 39.740 ;
        RECT 690.070 39.540 1604.870 39.680 ;
        RECT 690.070 39.480 690.390 39.540 ;
        RECT 1604.550 39.480 1604.870 39.540 ;
      LAYER via ;
        RECT 690.100 386.280 690.360 386.540 ;
        RECT 691.940 386.280 692.200 386.540 ;
        RECT 690.100 39.480 690.360 39.740 ;
        RECT 1604.580 39.480 1604.840 39.740 ;
      LAYER met2 ;
        RECT 692.290 400.250 692.570 404.000 ;
        RECT 692.000 400.110 692.570 400.250 ;
        RECT 692.000 386.570 692.140 400.110 ;
        RECT 692.290 400.000 692.570 400.110 ;
        RECT 690.100 386.250 690.360 386.570 ;
        RECT 691.940 386.250 692.200 386.570 ;
        RECT 690.160 39.770 690.300 386.250 ;
        RECT 690.100 39.450 690.360 39.770 ;
        RECT 1604.580 39.450 1604.840 39.770 ;
        RECT 1604.640 2.400 1604.780 39.450 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 696.970 39.340 697.290 39.400 ;
        RECT 1622.030 39.340 1622.350 39.400 ;
        RECT 696.970 39.200 1622.350 39.340 ;
        RECT 696.970 39.140 697.290 39.200 ;
        RECT 1622.030 39.140 1622.350 39.200 ;
      LAYER via ;
        RECT 697.000 39.140 697.260 39.400 ;
        RECT 1622.060 39.140 1622.320 39.400 ;
      LAYER met2 ;
        RECT 697.810 400.250 698.090 404.000 ;
        RECT 697.060 400.110 698.090 400.250 ;
        RECT 697.060 39.430 697.200 400.110 ;
        RECT 697.810 400.000 698.090 400.110 ;
        RECT 697.000 39.110 697.260 39.430 ;
        RECT 1622.060 39.110 1622.320 39.430 ;
        RECT 1622.120 2.400 1622.260 39.110 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.430 386.480 697.750 386.540 ;
        RECT 701.570 386.480 701.890 386.540 ;
        RECT 697.430 386.340 701.890 386.480 ;
        RECT 697.430 386.280 697.750 386.340 ;
        RECT 701.570 386.280 701.890 386.340 ;
        RECT 697.430 39.000 697.750 39.060 ;
        RECT 1639.970 39.000 1640.290 39.060 ;
        RECT 697.430 38.860 1640.290 39.000 ;
        RECT 697.430 38.800 697.750 38.860 ;
        RECT 1639.970 38.800 1640.290 38.860 ;
      LAYER via ;
        RECT 697.460 386.280 697.720 386.540 ;
        RECT 701.600 386.280 701.860 386.540 ;
        RECT 697.460 38.800 697.720 39.060 ;
        RECT 1640.000 38.800 1640.260 39.060 ;
      LAYER met2 ;
        RECT 702.870 400.250 703.150 404.000 ;
        RECT 701.660 400.110 703.150 400.250 ;
        RECT 701.660 386.570 701.800 400.110 ;
        RECT 702.870 400.000 703.150 400.110 ;
        RECT 697.460 386.250 697.720 386.570 ;
        RECT 701.600 386.250 701.860 386.570 ;
        RECT 697.520 39.090 697.660 386.250 ;
        RECT 697.460 38.770 697.720 39.090 ;
        RECT 1640.000 38.770 1640.260 39.090 ;
        RECT 1640.060 2.400 1640.200 38.770 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 703.870 386.140 704.190 386.200 ;
        RECT 707.090 386.140 707.410 386.200 ;
        RECT 703.870 386.000 707.410 386.140 ;
        RECT 703.870 385.940 704.190 386.000 ;
        RECT 707.090 385.940 707.410 386.000 ;
        RECT 703.870 38.660 704.190 38.720 ;
        RECT 1657.910 38.660 1658.230 38.720 ;
        RECT 703.870 38.520 1658.230 38.660 ;
        RECT 703.870 38.460 704.190 38.520 ;
        RECT 1657.910 38.460 1658.230 38.520 ;
      LAYER via ;
        RECT 703.900 385.940 704.160 386.200 ;
        RECT 707.120 385.940 707.380 386.200 ;
        RECT 703.900 38.460 704.160 38.720 ;
        RECT 1657.940 38.460 1658.200 38.720 ;
      LAYER met2 ;
        RECT 708.390 400.250 708.670 404.000 ;
        RECT 707.180 400.110 708.670 400.250 ;
        RECT 707.180 386.230 707.320 400.110 ;
        RECT 708.390 400.000 708.670 400.110 ;
        RECT 703.900 385.910 704.160 386.230 ;
        RECT 707.120 385.910 707.380 386.230 ;
        RECT 703.960 38.750 704.100 385.910 ;
        RECT 703.900 38.430 704.160 38.750 ;
        RECT 1657.940 38.430 1658.200 38.750 ;
        RECT 1658.000 2.400 1658.140 38.430 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 710.770 386.480 711.090 386.540 ;
        RECT 712.610 386.480 712.930 386.540 ;
        RECT 710.770 386.340 712.930 386.480 ;
        RECT 710.770 386.280 711.090 386.340 ;
        RECT 712.610 386.280 712.930 386.340 ;
        RECT 710.770 38.320 711.090 38.380 ;
        RECT 1675.390 38.320 1675.710 38.380 ;
        RECT 710.770 38.180 1675.710 38.320 ;
        RECT 710.770 38.120 711.090 38.180 ;
        RECT 1675.390 38.120 1675.710 38.180 ;
      LAYER via ;
        RECT 710.800 386.280 711.060 386.540 ;
        RECT 712.640 386.280 712.900 386.540 ;
        RECT 710.800 38.120 711.060 38.380 ;
        RECT 1675.420 38.120 1675.680 38.380 ;
      LAYER met2 ;
        RECT 713.910 400.250 714.190 404.000 ;
        RECT 712.700 400.110 714.190 400.250 ;
        RECT 712.700 386.570 712.840 400.110 ;
        RECT 713.910 400.000 714.190 400.110 ;
        RECT 710.800 386.250 711.060 386.570 ;
        RECT 712.640 386.250 712.900 386.570 ;
        RECT 710.860 38.410 711.000 386.250 ;
        RECT 710.800 38.090 711.060 38.410 ;
        RECT 1675.420 38.090 1675.680 38.410 ;
        RECT 1675.480 2.400 1675.620 38.090 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.070 384.440 414.390 384.500 ;
        RECT 418.670 384.440 418.990 384.500 ;
        RECT 414.070 384.300 418.990 384.440 ;
        RECT 414.070 384.240 414.390 384.300 ;
        RECT 418.670 384.240 418.990 384.300 ;
        RECT 414.070 27.440 414.390 27.500 ;
        RECT 717.670 27.440 717.990 27.500 ;
        RECT 414.070 27.300 717.990 27.440 ;
        RECT 414.070 27.240 414.390 27.300 ;
        RECT 717.670 27.240 717.990 27.300 ;
      LAYER via ;
        RECT 414.100 384.240 414.360 384.500 ;
        RECT 418.700 384.240 418.960 384.500 ;
        RECT 414.100 27.240 414.360 27.500 ;
        RECT 717.700 27.240 717.960 27.500 ;
      LAYER met2 ;
        RECT 419.970 400.250 420.250 404.000 ;
        RECT 418.760 400.110 420.250 400.250 ;
        RECT 418.760 384.530 418.900 400.110 ;
        RECT 419.970 400.000 420.250 400.110 ;
        RECT 414.100 384.210 414.360 384.530 ;
        RECT 418.700 384.210 418.960 384.530 ;
        RECT 414.160 27.530 414.300 384.210 ;
        RECT 414.100 27.210 414.360 27.530 ;
        RECT 717.700 27.210 717.960 27.530 ;
        RECT 717.760 2.400 717.900 27.210 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 717.670 386.140 717.990 386.200 ;
        RECT 719.510 386.140 719.830 386.200 ;
        RECT 717.670 386.000 719.830 386.140 ;
        RECT 717.670 385.940 717.990 386.000 ;
        RECT 719.510 385.940 719.830 386.000 ;
        RECT 717.670 37.980 717.990 38.040 ;
        RECT 1693.330 37.980 1693.650 38.040 ;
        RECT 717.670 37.840 1693.650 37.980 ;
        RECT 717.670 37.780 717.990 37.840 ;
        RECT 1693.330 37.780 1693.650 37.840 ;
      LAYER via ;
        RECT 717.700 385.940 717.960 386.200 ;
        RECT 719.540 385.940 719.800 386.200 ;
        RECT 717.700 37.780 717.960 38.040 ;
        RECT 1693.360 37.780 1693.620 38.040 ;
      LAYER met2 ;
        RECT 719.430 400.180 719.710 404.000 ;
        RECT 719.430 400.000 719.740 400.180 ;
        RECT 719.600 386.230 719.740 400.000 ;
        RECT 717.700 385.910 717.960 386.230 ;
        RECT 719.540 385.910 719.800 386.230 ;
        RECT 717.760 38.070 717.900 385.910 ;
        RECT 717.700 37.750 717.960 38.070 ;
        RECT 1693.360 37.750 1693.620 38.070 ;
        RECT 1693.420 2.400 1693.560 37.750 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.950 400.250 725.230 404.000 ;
        RECT 724.660 400.110 725.230 400.250 ;
        RECT 724.660 37.925 724.800 400.110 ;
        RECT 724.950 400.000 725.230 400.110 ;
        RECT 724.590 37.555 724.870 37.925 ;
        RECT 1710.830 37.555 1711.110 37.925 ;
        RECT 1710.900 2.400 1711.040 37.555 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
      LAYER via2 ;
        RECT 724.590 37.600 724.870 37.880 ;
        RECT 1710.830 37.600 1711.110 37.880 ;
      LAYER met3 ;
        RECT 724.565 37.890 724.895 37.905 ;
        RECT 1710.805 37.890 1711.135 37.905 ;
        RECT 724.565 37.590 1711.135 37.890 ;
        RECT 724.565 37.575 724.895 37.590 ;
        RECT 1710.805 37.575 1711.135 37.590 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.490 385.800 725.810 385.860 ;
        RECT 729.170 385.800 729.490 385.860 ;
        RECT 725.490 385.660 729.490 385.800 ;
        RECT 725.490 385.600 725.810 385.660 ;
        RECT 729.170 385.600 729.490 385.660 ;
        RECT 725.490 110.060 725.810 110.120 ;
        RECT 1725.070 110.060 1725.390 110.120 ;
        RECT 725.490 109.920 1725.390 110.060 ;
        RECT 725.490 109.860 725.810 109.920 ;
        RECT 1725.070 109.860 1725.390 109.920 ;
      LAYER via ;
        RECT 725.520 385.600 725.780 385.860 ;
        RECT 729.200 385.600 729.460 385.860 ;
        RECT 725.520 109.860 725.780 110.120 ;
        RECT 1725.100 109.860 1725.360 110.120 ;
      LAYER met2 ;
        RECT 730.470 400.250 730.750 404.000 ;
        RECT 729.260 400.110 730.750 400.250 ;
        RECT 729.260 385.890 729.400 400.110 ;
        RECT 730.470 400.000 730.750 400.110 ;
        RECT 725.520 385.570 725.780 385.890 ;
        RECT 729.200 385.570 729.460 385.890 ;
        RECT 725.580 110.150 725.720 385.570 ;
        RECT 725.520 109.830 725.780 110.150 ;
        RECT 1725.100 109.830 1725.360 110.150 ;
        RECT 1725.160 82.870 1725.300 109.830 ;
        RECT 1725.160 82.730 1726.680 82.870 ;
        RECT 1726.540 1.770 1726.680 82.730 ;
        RECT 1728.630 1.770 1729.190 2.400 ;
        RECT 1726.540 1.630 1729.190 1.770 ;
        RECT 1728.630 -4.800 1729.190 1.630 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.390 386.480 732.710 386.540 ;
        RECT 734.230 386.480 734.550 386.540 ;
        RECT 732.390 386.340 734.550 386.480 ;
        RECT 732.390 386.280 732.710 386.340 ;
        RECT 734.230 386.280 734.550 386.340 ;
        RECT 732.390 109.720 732.710 109.780 ;
        RECT 1745.770 109.720 1746.090 109.780 ;
        RECT 732.390 109.580 1746.090 109.720 ;
        RECT 732.390 109.520 732.710 109.580 ;
        RECT 1745.770 109.520 1746.090 109.580 ;
      LAYER via ;
        RECT 732.420 386.280 732.680 386.540 ;
        RECT 734.260 386.280 734.520 386.540 ;
        RECT 732.420 109.520 732.680 109.780 ;
        RECT 1745.800 109.520 1746.060 109.780 ;
      LAYER met2 ;
        RECT 735.530 400.250 735.810 404.000 ;
        RECT 734.320 400.110 735.810 400.250 ;
        RECT 734.320 386.570 734.460 400.110 ;
        RECT 735.530 400.000 735.810 400.110 ;
        RECT 732.420 386.250 732.680 386.570 ;
        RECT 734.260 386.250 734.520 386.570 ;
        RECT 732.480 109.810 732.620 386.250 ;
        RECT 732.420 109.490 732.680 109.810 ;
        RECT 1745.800 109.490 1746.060 109.810 ;
        RECT 1745.860 14.690 1746.000 109.490 ;
        RECT 1745.860 14.550 1746.460 14.690 ;
        RECT 1746.320 2.400 1746.460 14.550 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.830 386.480 739.150 386.540 ;
        RECT 739.750 386.480 740.070 386.540 ;
        RECT 738.830 386.340 740.070 386.480 ;
        RECT 738.830 386.280 739.150 386.340 ;
        RECT 739.750 386.280 740.070 386.340 ;
        RECT 738.830 109.380 739.150 109.440 ;
        RECT 1759.570 109.380 1759.890 109.440 ;
        RECT 738.830 109.240 1759.890 109.380 ;
        RECT 738.830 109.180 739.150 109.240 ;
        RECT 1759.570 109.180 1759.890 109.240 ;
      LAYER via ;
        RECT 738.860 386.280 739.120 386.540 ;
        RECT 739.780 386.280 740.040 386.540 ;
        RECT 738.860 109.180 739.120 109.440 ;
        RECT 1759.600 109.180 1759.860 109.440 ;
      LAYER met2 ;
        RECT 741.050 400.250 741.330 404.000 ;
        RECT 739.840 400.110 741.330 400.250 ;
        RECT 739.840 386.570 739.980 400.110 ;
        RECT 741.050 400.000 741.330 400.110 ;
        RECT 738.860 386.250 739.120 386.570 ;
        RECT 739.780 386.250 740.040 386.570 ;
        RECT 738.920 109.470 739.060 386.250 ;
        RECT 738.860 109.150 739.120 109.470 ;
        RECT 1759.600 109.150 1759.860 109.470 ;
        RECT 1759.660 82.870 1759.800 109.150 ;
        RECT 1759.660 82.730 1764.400 82.870 ;
        RECT 1764.260 2.400 1764.400 82.730 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.730 117.200 746.050 117.260 ;
        RECT 1780.270 117.200 1780.590 117.260 ;
        RECT 745.730 117.060 1780.590 117.200 ;
        RECT 745.730 117.000 746.050 117.060 ;
        RECT 1780.270 117.000 1780.590 117.060 ;
      LAYER via ;
        RECT 745.760 117.000 746.020 117.260 ;
        RECT 1780.300 117.000 1780.560 117.260 ;
      LAYER met2 ;
        RECT 746.570 400.250 746.850 404.000 ;
        RECT 745.820 400.110 746.850 400.250 ;
        RECT 745.820 117.290 745.960 400.110 ;
        RECT 746.570 400.000 746.850 400.110 ;
        RECT 745.760 116.970 746.020 117.290 ;
        RECT 1780.300 116.970 1780.560 117.290 ;
        RECT 1780.360 82.870 1780.500 116.970 ;
        RECT 1780.360 82.730 1781.880 82.870 ;
        RECT 1781.740 2.400 1781.880 82.730 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.170 387.160 752.490 387.220 ;
        RECT 753.090 387.160 753.410 387.220 ;
        RECT 752.170 387.020 753.410 387.160 ;
        RECT 752.170 386.960 752.490 387.020 ;
        RECT 753.090 386.960 753.410 387.020 ;
        RECT 753.090 116.860 753.410 116.920 ;
        RECT 1794.070 116.860 1794.390 116.920 ;
        RECT 753.090 116.720 1794.390 116.860 ;
        RECT 753.090 116.660 753.410 116.720 ;
        RECT 1794.070 116.660 1794.390 116.720 ;
      LAYER via ;
        RECT 752.200 386.960 752.460 387.220 ;
        RECT 753.120 386.960 753.380 387.220 ;
        RECT 753.120 116.660 753.380 116.920 ;
        RECT 1794.100 116.660 1794.360 116.920 ;
      LAYER met2 ;
        RECT 752.090 400.180 752.370 404.000 ;
        RECT 752.090 400.000 752.400 400.180 ;
        RECT 752.260 387.250 752.400 400.000 ;
        RECT 752.200 386.930 752.460 387.250 ;
        RECT 753.120 386.930 753.380 387.250 ;
        RECT 753.180 116.950 753.320 386.930 ;
        RECT 753.120 116.630 753.380 116.950 ;
        RECT 1794.100 116.630 1794.360 116.950 ;
        RECT 1794.160 82.870 1794.300 116.630 ;
        RECT 1794.160 82.730 1797.520 82.870 ;
        RECT 1797.380 1.770 1797.520 82.730 ;
        RECT 1799.470 1.770 1800.030 2.400 ;
        RECT 1797.380 1.630 1800.030 1.770 ;
        RECT 1799.470 -4.800 1800.030 1.630 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.170 386.480 752.490 386.540 ;
        RECT 756.310 386.480 756.630 386.540 ;
        RECT 752.170 386.340 756.630 386.480 ;
        RECT 752.170 386.280 752.490 386.340 ;
        RECT 756.310 386.280 756.630 386.340 ;
        RECT 752.170 43.420 752.490 43.480 ;
        RECT 1817.530 43.420 1817.850 43.480 ;
        RECT 752.170 43.280 1817.850 43.420 ;
        RECT 752.170 43.220 752.490 43.280 ;
        RECT 1817.530 43.220 1817.850 43.280 ;
      LAYER via ;
        RECT 752.200 386.280 752.460 386.540 ;
        RECT 756.340 386.280 756.600 386.540 ;
        RECT 752.200 43.220 752.460 43.480 ;
        RECT 1817.560 43.220 1817.820 43.480 ;
      LAYER met2 ;
        RECT 757.610 400.250 757.890 404.000 ;
        RECT 756.400 400.110 757.890 400.250 ;
        RECT 756.400 386.570 756.540 400.110 ;
        RECT 757.610 400.000 757.890 400.110 ;
        RECT 752.200 386.250 752.460 386.570 ;
        RECT 756.340 386.250 756.600 386.570 ;
        RECT 752.260 43.510 752.400 386.250 ;
        RECT 752.200 43.190 752.460 43.510 ;
        RECT 1817.560 43.190 1817.820 43.510 ;
        RECT 1817.620 2.400 1817.760 43.190 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.070 386.480 759.390 386.540 ;
        RECT 761.830 386.480 762.150 386.540 ;
        RECT 759.070 386.340 762.150 386.480 ;
        RECT 759.070 386.280 759.390 386.340 ;
        RECT 761.830 386.280 762.150 386.340 ;
        RECT 759.530 43.760 759.850 43.820 ;
        RECT 1835.010 43.760 1835.330 43.820 ;
        RECT 759.530 43.620 1835.330 43.760 ;
        RECT 759.530 43.560 759.850 43.620 ;
        RECT 1835.010 43.560 1835.330 43.620 ;
      LAYER via ;
        RECT 759.100 386.280 759.360 386.540 ;
        RECT 761.860 386.280 762.120 386.540 ;
        RECT 759.560 43.560 759.820 43.820 ;
        RECT 1835.040 43.560 1835.300 43.820 ;
      LAYER met2 ;
        RECT 763.130 400.250 763.410 404.000 ;
        RECT 761.920 400.110 763.410 400.250 ;
        RECT 761.920 386.570 762.060 400.110 ;
        RECT 763.130 400.000 763.410 400.110 ;
        RECT 759.100 386.250 759.360 386.570 ;
        RECT 761.860 386.250 762.120 386.570 ;
        RECT 759.160 63.650 759.300 386.250 ;
        RECT 759.160 63.510 759.760 63.650 ;
        RECT 759.620 43.850 759.760 63.510 ;
        RECT 759.560 43.530 759.820 43.850 ;
        RECT 1835.040 43.530 1835.300 43.850 ;
        RECT 1835.100 2.400 1835.240 43.530 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 765.970 44.100 766.290 44.160 ;
        RECT 1852.950 44.100 1853.270 44.160 ;
        RECT 765.970 43.960 1853.270 44.100 ;
        RECT 765.970 43.900 766.290 43.960 ;
        RECT 1852.950 43.900 1853.270 43.960 ;
      LAYER via ;
        RECT 766.000 43.900 766.260 44.160 ;
        RECT 1852.980 43.900 1853.240 44.160 ;
      LAYER met2 ;
        RECT 768.190 400.250 768.470 404.000 ;
        RECT 767.440 400.110 768.470 400.250 ;
        RECT 767.440 386.650 767.580 400.110 ;
        RECT 768.190 400.000 768.470 400.110 ;
        RECT 766.060 386.510 767.580 386.650 ;
        RECT 766.060 44.190 766.200 386.510 ;
        RECT 766.000 43.870 766.260 44.190 ;
        RECT 1852.980 43.870 1853.240 44.190 ;
        RECT 1853.040 2.400 1853.180 43.870 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 420.970 374.240 421.290 374.300 ;
        RECT 424.190 374.240 424.510 374.300 ;
        RECT 420.970 374.100 424.510 374.240 ;
        RECT 420.970 374.040 421.290 374.100 ;
        RECT 424.190 374.040 424.510 374.100 ;
        RECT 420.970 27.100 421.290 27.160 ;
        RECT 735.610 27.100 735.930 27.160 ;
        RECT 420.970 26.960 735.930 27.100 ;
        RECT 420.970 26.900 421.290 26.960 ;
        RECT 735.610 26.900 735.930 26.960 ;
      LAYER via ;
        RECT 421.000 374.040 421.260 374.300 ;
        RECT 424.220 374.040 424.480 374.300 ;
        RECT 421.000 26.900 421.260 27.160 ;
        RECT 735.640 26.900 735.900 27.160 ;
      LAYER met2 ;
        RECT 425.490 400.250 425.770 404.000 ;
        RECT 424.280 400.110 425.770 400.250 ;
        RECT 424.280 374.330 424.420 400.110 ;
        RECT 425.490 400.000 425.770 400.110 ;
        RECT 421.000 374.010 421.260 374.330 ;
        RECT 424.220 374.010 424.480 374.330 ;
        RECT 421.060 27.190 421.200 374.010 ;
        RECT 421.000 26.870 421.260 27.190 ;
        RECT 735.640 26.870 735.900 27.190 ;
        RECT 735.700 2.400 735.840 26.870 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 772.870 44.440 773.190 44.500 ;
        RECT 1870.430 44.440 1870.750 44.500 ;
        RECT 772.870 44.300 1870.750 44.440 ;
        RECT 772.870 44.240 773.190 44.300 ;
        RECT 1870.430 44.240 1870.750 44.300 ;
      LAYER via ;
        RECT 772.900 44.240 773.160 44.500 ;
        RECT 1870.460 44.240 1870.720 44.500 ;
      LAYER met2 ;
        RECT 773.710 400.250 773.990 404.000 ;
        RECT 772.960 400.110 773.990 400.250 ;
        RECT 772.960 44.530 773.100 400.110 ;
        RECT 773.710 400.000 773.990 400.110 ;
        RECT 772.900 44.210 773.160 44.530 ;
        RECT 1870.460 44.210 1870.720 44.530 ;
        RECT 1870.520 2.400 1870.660 44.210 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.330 386.480 773.650 386.540 ;
        RECT 777.930 386.480 778.250 386.540 ;
        RECT 773.330 386.340 778.250 386.480 ;
        RECT 773.330 386.280 773.650 386.340 ;
        RECT 777.930 386.280 778.250 386.340 ;
        RECT 773.330 48.180 773.650 48.240 ;
        RECT 1888.370 48.180 1888.690 48.240 ;
        RECT 773.330 48.040 1888.690 48.180 ;
        RECT 773.330 47.980 773.650 48.040 ;
        RECT 1888.370 47.980 1888.690 48.040 ;
      LAYER via ;
        RECT 773.360 386.280 773.620 386.540 ;
        RECT 777.960 386.280 778.220 386.540 ;
        RECT 773.360 47.980 773.620 48.240 ;
        RECT 1888.400 47.980 1888.660 48.240 ;
      LAYER met2 ;
        RECT 779.230 400.250 779.510 404.000 ;
        RECT 778.020 400.110 779.510 400.250 ;
        RECT 778.020 386.570 778.160 400.110 ;
        RECT 779.230 400.000 779.510 400.110 ;
        RECT 773.360 386.250 773.620 386.570 ;
        RECT 777.960 386.250 778.220 386.570 ;
        RECT 773.420 48.270 773.560 386.250 ;
        RECT 773.360 47.950 773.620 48.270 ;
        RECT 1888.400 47.950 1888.660 48.270 ;
        RECT 1888.460 2.400 1888.600 47.950 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 779.770 386.480 780.090 386.540 ;
        RECT 783.450 386.480 783.770 386.540 ;
        RECT 779.770 386.340 783.770 386.480 ;
        RECT 779.770 386.280 780.090 386.340 ;
        RECT 783.450 386.280 783.770 386.340 ;
        RECT 779.770 47.840 780.090 47.900 ;
        RECT 1905.850 47.840 1906.170 47.900 ;
        RECT 779.770 47.700 1906.170 47.840 ;
        RECT 779.770 47.640 780.090 47.700 ;
        RECT 1905.850 47.640 1906.170 47.700 ;
      LAYER via ;
        RECT 779.800 386.280 780.060 386.540 ;
        RECT 783.480 386.280 783.740 386.540 ;
        RECT 779.800 47.640 780.060 47.900 ;
        RECT 1905.880 47.640 1906.140 47.900 ;
      LAYER met2 ;
        RECT 784.750 400.250 785.030 404.000 ;
        RECT 783.540 400.110 785.030 400.250 ;
        RECT 783.540 386.570 783.680 400.110 ;
        RECT 784.750 400.000 785.030 400.110 ;
        RECT 779.800 386.250 780.060 386.570 ;
        RECT 783.480 386.250 783.740 386.570 ;
        RECT 779.860 47.930 780.000 386.250 ;
        RECT 779.800 47.610 780.060 47.930 ;
        RECT 1905.880 47.610 1906.140 47.930 ;
        RECT 1905.940 2.400 1906.080 47.610 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 786.670 376.280 786.990 376.340 ;
        RECT 788.970 376.280 789.290 376.340 ;
        RECT 786.670 376.140 789.290 376.280 ;
        RECT 786.670 376.080 786.990 376.140 ;
        RECT 788.970 376.080 789.290 376.140 ;
        RECT 786.670 47.500 786.990 47.560 ;
        RECT 1923.790 47.500 1924.110 47.560 ;
        RECT 786.670 47.360 1924.110 47.500 ;
        RECT 786.670 47.300 786.990 47.360 ;
        RECT 1923.790 47.300 1924.110 47.360 ;
      LAYER via ;
        RECT 786.700 376.080 786.960 376.340 ;
        RECT 789.000 376.080 789.260 376.340 ;
        RECT 786.700 47.300 786.960 47.560 ;
        RECT 1923.820 47.300 1924.080 47.560 ;
      LAYER met2 ;
        RECT 790.270 400.250 790.550 404.000 ;
        RECT 789.060 400.110 790.550 400.250 ;
        RECT 789.060 376.370 789.200 400.110 ;
        RECT 790.270 400.000 790.550 400.110 ;
        RECT 786.700 376.050 786.960 376.370 ;
        RECT 789.000 376.050 789.260 376.370 ;
        RECT 786.760 47.590 786.900 376.050 ;
        RECT 786.700 47.270 786.960 47.590 ;
        RECT 1923.820 47.270 1924.080 47.590 ;
        RECT 1923.880 2.400 1924.020 47.270 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 793.570 377.640 793.890 377.700 ;
        RECT 794.490 377.640 794.810 377.700 ;
        RECT 793.570 377.500 794.810 377.640 ;
        RECT 793.570 377.440 793.890 377.500 ;
        RECT 794.490 377.440 794.810 377.500 ;
        RECT 793.570 47.160 793.890 47.220 ;
        RECT 1941.270 47.160 1941.590 47.220 ;
        RECT 793.570 47.020 1941.590 47.160 ;
        RECT 793.570 46.960 793.890 47.020 ;
        RECT 1941.270 46.960 1941.590 47.020 ;
      LAYER via ;
        RECT 793.600 377.440 793.860 377.700 ;
        RECT 794.520 377.440 794.780 377.700 ;
        RECT 793.600 46.960 793.860 47.220 ;
        RECT 1941.300 46.960 1941.560 47.220 ;
      LAYER met2 ;
        RECT 795.790 400.250 796.070 404.000 ;
        RECT 794.580 400.110 796.070 400.250 ;
        RECT 794.580 377.730 794.720 400.110 ;
        RECT 795.790 400.000 796.070 400.110 ;
        RECT 793.600 377.410 793.860 377.730 ;
        RECT 794.520 377.410 794.780 377.730 ;
        RECT 793.660 47.250 793.800 377.410 ;
        RECT 793.600 46.930 793.860 47.250 ;
        RECT 1941.300 46.930 1941.560 47.250 ;
        RECT 1941.360 2.400 1941.500 46.930 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.470 46.820 800.790 46.880 ;
        RECT 1959.210 46.820 1959.530 46.880 ;
        RECT 800.470 46.680 1959.530 46.820 ;
        RECT 800.470 46.620 800.790 46.680 ;
        RECT 1959.210 46.620 1959.530 46.680 ;
      LAYER via ;
        RECT 800.500 46.620 800.760 46.880 ;
        RECT 1959.240 46.620 1959.500 46.880 ;
      LAYER met2 ;
        RECT 800.850 400.250 801.130 404.000 ;
        RECT 800.560 400.110 801.130 400.250 ;
        RECT 800.560 46.910 800.700 400.110 ;
        RECT 800.850 400.000 801.130 400.110 ;
        RECT 800.500 46.590 800.760 46.910 ;
        RECT 1959.240 46.590 1959.500 46.910 ;
        RECT 1959.300 2.400 1959.440 46.590 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 800.930 376.280 801.250 376.340 ;
        RECT 805.070 376.280 805.390 376.340 ;
        RECT 800.930 376.140 805.390 376.280 ;
        RECT 800.930 376.080 801.250 376.140 ;
        RECT 805.070 376.080 805.390 376.140 ;
        RECT 800.930 46.480 801.250 46.540 ;
        RECT 1976.690 46.480 1977.010 46.540 ;
        RECT 800.930 46.340 1977.010 46.480 ;
        RECT 800.930 46.280 801.250 46.340 ;
        RECT 1976.690 46.280 1977.010 46.340 ;
      LAYER via ;
        RECT 800.960 376.080 801.220 376.340 ;
        RECT 805.100 376.080 805.360 376.340 ;
        RECT 800.960 46.280 801.220 46.540 ;
        RECT 1976.720 46.280 1976.980 46.540 ;
      LAYER met2 ;
        RECT 806.370 400.250 806.650 404.000 ;
        RECT 805.160 400.110 806.650 400.250 ;
        RECT 805.160 376.370 805.300 400.110 ;
        RECT 806.370 400.000 806.650 400.110 ;
        RECT 800.960 376.050 801.220 376.370 ;
        RECT 805.100 376.050 805.360 376.370 ;
        RECT 801.020 46.570 801.160 376.050 ;
        RECT 800.960 46.250 801.220 46.570 ;
        RECT 1976.720 46.250 1976.980 46.570 ;
        RECT 1976.780 2.400 1976.920 46.250 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.370 376.280 807.690 376.340 ;
        RECT 810.590 376.280 810.910 376.340 ;
        RECT 807.370 376.140 810.910 376.280 ;
        RECT 807.370 376.080 807.690 376.140 ;
        RECT 810.590 376.080 810.910 376.140 ;
        RECT 807.370 46.140 807.690 46.200 ;
        RECT 1994.630 46.140 1994.950 46.200 ;
        RECT 807.370 46.000 1994.950 46.140 ;
        RECT 807.370 45.940 807.690 46.000 ;
        RECT 1994.630 45.940 1994.950 46.000 ;
      LAYER via ;
        RECT 807.400 376.080 807.660 376.340 ;
        RECT 810.620 376.080 810.880 376.340 ;
        RECT 807.400 45.940 807.660 46.200 ;
        RECT 1994.660 45.940 1994.920 46.200 ;
      LAYER met2 ;
        RECT 811.890 400.250 812.170 404.000 ;
        RECT 810.680 400.110 812.170 400.250 ;
        RECT 810.680 376.370 810.820 400.110 ;
        RECT 811.890 400.000 812.170 400.110 ;
        RECT 807.400 376.050 807.660 376.370 ;
        RECT 810.620 376.050 810.880 376.370 ;
        RECT 807.460 46.230 807.600 376.050 ;
        RECT 807.400 45.910 807.660 46.230 ;
        RECT 1994.660 45.910 1994.920 46.230 ;
        RECT 1994.720 2.400 1994.860 45.910 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.270 375.940 814.590 376.000 ;
        RECT 816.110 375.940 816.430 376.000 ;
        RECT 814.270 375.800 816.430 375.940 ;
        RECT 814.270 375.740 814.590 375.800 ;
        RECT 816.110 375.740 816.430 375.800 ;
        RECT 814.270 45.800 814.590 45.860 ;
        RECT 2012.570 45.800 2012.890 45.860 ;
        RECT 814.270 45.660 2012.890 45.800 ;
        RECT 814.270 45.600 814.590 45.660 ;
        RECT 2012.570 45.600 2012.890 45.660 ;
      LAYER via ;
        RECT 814.300 375.740 814.560 376.000 ;
        RECT 816.140 375.740 816.400 376.000 ;
        RECT 814.300 45.600 814.560 45.860 ;
        RECT 2012.600 45.600 2012.860 45.860 ;
      LAYER met2 ;
        RECT 817.410 400.250 817.690 404.000 ;
        RECT 816.200 400.110 817.690 400.250 ;
        RECT 816.200 376.030 816.340 400.110 ;
        RECT 817.410 400.000 817.690 400.110 ;
        RECT 814.300 375.710 814.560 376.030 ;
        RECT 816.140 375.710 816.400 376.030 ;
        RECT 814.360 45.890 814.500 375.710 ;
        RECT 814.300 45.570 814.560 45.890 ;
        RECT 2012.600 45.570 2012.860 45.890 ;
        RECT 2012.660 2.400 2012.800 45.570 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.170 45.460 821.490 45.520 ;
        RECT 2030.050 45.460 2030.370 45.520 ;
        RECT 821.170 45.320 2030.370 45.460 ;
        RECT 821.170 45.260 821.490 45.320 ;
        RECT 2030.050 45.260 2030.370 45.320 ;
      LAYER via ;
        RECT 821.200 45.260 821.460 45.520 ;
        RECT 2030.080 45.260 2030.340 45.520 ;
      LAYER met2 ;
        RECT 822.930 400.250 823.210 404.000 ;
        RECT 822.640 400.110 823.210 400.250 ;
        RECT 822.640 390.050 822.780 400.110 ;
        RECT 822.930 400.000 823.210 400.110 ;
        RECT 821.260 389.910 822.780 390.050 ;
        RECT 821.260 45.550 821.400 389.910 ;
        RECT 821.200 45.230 821.460 45.550 ;
        RECT 2030.080 45.230 2030.340 45.550 ;
        RECT 2030.140 2.400 2030.280 45.230 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.870 387.160 428.190 387.220 ;
        RECT 429.710 387.160 430.030 387.220 ;
        RECT 427.870 387.020 430.030 387.160 ;
        RECT 427.870 386.960 428.190 387.020 ;
        RECT 429.710 386.960 430.030 387.020 ;
        RECT 427.870 26.760 428.190 26.820 ;
        RECT 753.090 26.760 753.410 26.820 ;
        RECT 427.870 26.620 753.410 26.760 ;
        RECT 427.870 26.560 428.190 26.620 ;
        RECT 753.090 26.560 753.410 26.620 ;
      LAYER via ;
        RECT 427.900 386.960 428.160 387.220 ;
        RECT 429.740 386.960 430.000 387.220 ;
        RECT 427.900 26.560 428.160 26.820 ;
        RECT 753.120 26.560 753.380 26.820 ;
      LAYER met2 ;
        RECT 431.010 400.250 431.290 404.000 ;
        RECT 429.800 400.110 431.290 400.250 ;
        RECT 429.800 387.250 429.940 400.110 ;
        RECT 431.010 400.000 431.290 400.110 ;
        RECT 427.900 386.930 428.160 387.250 ;
        RECT 429.740 386.930 430.000 387.250 ;
        RECT 427.960 26.850 428.100 386.930 ;
        RECT 427.900 26.530 428.160 26.850 ;
        RECT 753.120 26.530 753.380 26.850 ;
        RECT 753.180 2.400 753.320 26.530 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.070 45.120 828.390 45.180 ;
        RECT 2047.990 45.120 2048.310 45.180 ;
        RECT 828.070 44.980 2048.310 45.120 ;
        RECT 828.070 44.920 828.390 44.980 ;
        RECT 2047.990 44.920 2048.310 44.980 ;
      LAYER via ;
        RECT 828.100 44.920 828.360 45.180 ;
        RECT 2048.020 44.920 2048.280 45.180 ;
      LAYER met2 ;
        RECT 828.450 400.250 828.730 404.000 ;
        RECT 828.160 400.110 828.730 400.250 ;
        RECT 828.160 45.210 828.300 400.110 ;
        RECT 828.450 400.000 828.730 400.110 ;
        RECT 828.100 44.890 828.360 45.210 ;
        RECT 2048.020 44.890 2048.280 45.210 ;
        RECT 2048.080 2.400 2048.220 44.890 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.530 376.280 828.850 376.340 ;
        RECT 832.670 376.280 832.990 376.340 ;
        RECT 828.530 376.140 832.990 376.280 ;
        RECT 828.530 376.080 828.850 376.140 ;
        RECT 832.670 376.080 832.990 376.140 ;
        RECT 828.530 44.780 828.850 44.840 ;
        RECT 2065.470 44.780 2065.790 44.840 ;
        RECT 828.530 44.640 2065.790 44.780 ;
        RECT 828.530 44.580 828.850 44.640 ;
        RECT 2065.470 44.580 2065.790 44.640 ;
      LAYER via ;
        RECT 828.560 376.080 828.820 376.340 ;
        RECT 832.700 376.080 832.960 376.340 ;
        RECT 828.560 44.580 828.820 44.840 ;
        RECT 2065.500 44.580 2065.760 44.840 ;
      LAYER met2 ;
        RECT 833.970 400.250 834.250 404.000 ;
        RECT 832.760 400.110 834.250 400.250 ;
        RECT 832.760 376.370 832.900 400.110 ;
        RECT 833.970 400.000 834.250 400.110 ;
        RECT 828.560 376.050 828.820 376.370 ;
        RECT 832.700 376.050 832.960 376.370 ;
        RECT 828.620 44.870 828.760 376.050 ;
        RECT 828.560 44.550 828.820 44.870 ;
        RECT 2065.500 44.550 2065.760 44.870 ;
        RECT 2065.560 2.400 2065.700 44.550 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 834.970 375.940 835.290 376.000 ;
        RECT 837.730 375.940 838.050 376.000 ;
        RECT 834.970 375.800 838.050 375.940 ;
        RECT 834.970 375.740 835.290 375.800 ;
        RECT 837.730 375.740 838.050 375.800 ;
      LAYER via ;
        RECT 835.000 375.740 835.260 376.000 ;
        RECT 837.760 375.740 838.020 376.000 ;
      LAYER met2 ;
        RECT 839.030 400.250 839.310 404.000 ;
        RECT 837.820 400.110 839.310 400.250 ;
        RECT 837.820 376.030 837.960 400.110 ;
        RECT 839.030 400.000 839.310 400.110 ;
        RECT 835.000 375.710 835.260 376.030 ;
        RECT 837.760 375.710 838.020 376.030 ;
        RECT 835.060 45.405 835.200 375.710 ;
        RECT 834.990 45.035 835.270 45.405 ;
        RECT 2083.430 45.035 2083.710 45.405 ;
        RECT 2083.500 2.400 2083.640 45.035 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
      LAYER via2 ;
        RECT 834.990 45.080 835.270 45.360 ;
        RECT 2083.430 45.080 2083.710 45.360 ;
      LAYER met3 ;
        RECT 834.965 45.370 835.295 45.385 ;
        RECT 2083.405 45.370 2083.735 45.385 ;
        RECT 834.965 45.070 2083.735 45.370 ;
        RECT 834.965 45.055 835.295 45.070 ;
        RECT 2083.405 45.055 2083.735 45.070 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.550 400.250 844.830 404.000 ;
        RECT 843.340 400.110 844.830 400.250 ;
        RECT 843.340 389.370 843.480 400.110 ;
        RECT 844.550 400.000 844.830 400.110 ;
        RECT 841.960 389.230 843.480 389.370 ;
        RECT 841.960 44.725 842.100 389.230 ;
        RECT 841.890 44.355 842.170 44.725 ;
        RECT 2100.910 44.355 2101.190 44.725 ;
        RECT 2100.980 2.400 2101.120 44.355 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
      LAYER via2 ;
        RECT 841.890 44.400 842.170 44.680 ;
        RECT 2100.910 44.400 2101.190 44.680 ;
      LAYER met3 ;
        RECT 841.865 44.690 842.195 44.705 ;
        RECT 2100.885 44.690 2101.215 44.705 ;
        RECT 841.865 44.390 2101.215 44.690 ;
        RECT 841.865 44.375 842.195 44.390 ;
        RECT 2100.885 44.375 2101.215 44.390 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 849.230 116.520 849.550 116.580 ;
        RECT 2118.370 116.520 2118.690 116.580 ;
        RECT 849.230 116.380 2118.690 116.520 ;
        RECT 849.230 116.320 849.550 116.380 ;
        RECT 2118.370 116.320 2118.690 116.380 ;
      LAYER via ;
        RECT 849.260 116.320 849.520 116.580 ;
        RECT 2118.400 116.320 2118.660 116.580 ;
      LAYER met2 ;
        RECT 850.070 400.250 850.350 404.000 ;
        RECT 849.320 400.110 850.350 400.250 ;
        RECT 849.320 116.610 849.460 400.110 ;
        RECT 850.070 400.000 850.350 400.110 ;
        RECT 849.260 116.290 849.520 116.610 ;
        RECT 2118.400 116.290 2118.660 116.610 ;
        RECT 2118.460 14.690 2118.600 116.290 ;
        RECT 2118.460 14.550 2119.060 14.690 ;
        RECT 2118.920 2.400 2119.060 14.550 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 855.670 376.280 855.990 376.340 ;
        RECT 857.050 376.280 857.370 376.340 ;
        RECT 855.670 376.140 857.370 376.280 ;
        RECT 855.670 376.080 855.990 376.140 ;
        RECT 857.050 376.080 857.370 376.140 ;
        RECT 857.050 116.180 857.370 116.240 ;
        RECT 2132.170 116.180 2132.490 116.240 ;
        RECT 857.050 116.040 2132.490 116.180 ;
        RECT 857.050 115.980 857.370 116.040 ;
        RECT 2132.170 115.980 2132.490 116.040 ;
      LAYER via ;
        RECT 855.700 376.080 855.960 376.340 ;
        RECT 857.080 376.080 857.340 376.340 ;
        RECT 857.080 115.980 857.340 116.240 ;
        RECT 2132.200 115.980 2132.460 116.240 ;
      LAYER met2 ;
        RECT 855.590 400.180 855.870 404.000 ;
        RECT 855.590 400.000 855.900 400.180 ;
        RECT 855.760 376.370 855.900 400.000 ;
        RECT 855.700 376.050 855.960 376.370 ;
        RECT 857.080 376.050 857.340 376.370 ;
        RECT 857.140 116.270 857.280 376.050 ;
        RECT 857.080 115.950 857.340 116.270 ;
        RECT 2132.200 115.950 2132.460 116.270 ;
        RECT 2132.260 82.870 2132.400 115.950 ;
        RECT 2132.260 82.730 2134.240 82.870 ;
        RECT 2134.100 1.770 2134.240 82.730 ;
        RECT 2136.190 1.770 2136.750 2.400 ;
        RECT 2134.100 1.630 2136.750 1.770 ;
        RECT 2136.190 -4.800 2136.750 1.630 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.590 375.940 856.910 376.000 ;
        RECT 859.810 375.940 860.130 376.000 ;
        RECT 856.590 375.800 860.130 375.940 ;
        RECT 856.590 375.740 856.910 375.800 ;
        RECT 859.810 375.740 860.130 375.800 ;
        RECT 856.590 115.840 856.910 115.900 ;
        RECT 2152.870 115.840 2153.190 115.900 ;
        RECT 856.590 115.700 2153.190 115.840 ;
        RECT 856.590 115.640 856.910 115.700 ;
        RECT 2152.870 115.640 2153.190 115.700 ;
      LAYER via ;
        RECT 856.620 375.740 856.880 376.000 ;
        RECT 859.840 375.740 860.100 376.000 ;
        RECT 856.620 115.640 856.880 115.900 ;
        RECT 2152.900 115.640 2153.160 115.900 ;
      LAYER met2 ;
        RECT 861.110 400.250 861.390 404.000 ;
        RECT 859.900 400.110 861.390 400.250 ;
        RECT 859.900 376.030 860.040 400.110 ;
        RECT 861.110 400.000 861.390 400.110 ;
        RECT 856.620 375.710 856.880 376.030 ;
        RECT 859.840 375.710 860.100 376.030 ;
        RECT 856.680 115.930 856.820 375.710 ;
        RECT 856.620 115.610 856.880 115.930 ;
        RECT 2152.900 115.610 2153.160 115.930 ;
        RECT 2152.960 82.870 2153.100 115.610 ;
        RECT 2152.960 82.730 2154.480 82.870 ;
        RECT 2154.340 2.400 2154.480 82.730 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.950 115.500 864.270 115.560 ;
        RECT 2166.670 115.500 2166.990 115.560 ;
        RECT 863.950 115.360 2166.990 115.500 ;
        RECT 863.950 115.300 864.270 115.360 ;
        RECT 2166.670 115.300 2166.990 115.360 ;
      LAYER via ;
        RECT 863.980 115.300 864.240 115.560 ;
        RECT 2166.700 115.300 2166.960 115.560 ;
      LAYER met2 ;
        RECT 866.630 400.250 866.910 404.000 ;
        RECT 865.420 400.110 866.910 400.250 ;
        RECT 865.420 324.370 865.560 400.110 ;
        RECT 866.630 400.000 866.910 400.110 ;
        RECT 864.040 324.230 865.560 324.370 ;
        RECT 864.040 115.590 864.180 324.230 ;
        RECT 863.980 115.270 864.240 115.590 ;
        RECT 2166.700 115.270 2166.960 115.590 ;
        RECT 2166.760 82.870 2166.900 115.270 ;
        RECT 2166.760 82.730 2170.120 82.870 ;
        RECT 2169.980 1.770 2170.120 82.730 ;
        RECT 2172.070 1.770 2172.630 2.400 ;
        RECT 2169.980 1.630 2172.630 1.770 ;
        RECT 2172.070 -4.800 2172.630 1.630 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 870.850 115.160 871.170 115.220 ;
        RECT 2187.370 115.160 2187.690 115.220 ;
        RECT 870.850 115.020 2187.690 115.160 ;
        RECT 870.850 114.960 871.170 115.020 ;
        RECT 2187.370 114.960 2187.690 115.020 ;
      LAYER via ;
        RECT 870.880 114.960 871.140 115.220 ;
        RECT 2187.400 114.960 2187.660 115.220 ;
      LAYER met2 ;
        RECT 871.690 400.250 871.970 404.000 ;
        RECT 871.400 400.110 871.970 400.250 ;
        RECT 871.400 351.970 871.540 400.110 ;
        RECT 871.690 400.000 871.970 400.110 ;
        RECT 870.940 351.830 871.540 351.970 ;
        RECT 870.940 115.250 871.080 351.830 ;
        RECT 870.880 114.930 871.140 115.250 ;
        RECT 2187.400 114.930 2187.660 115.250 ;
        RECT 2187.460 1.770 2187.600 114.930 ;
        RECT 2189.550 1.770 2190.110 2.400 ;
        RECT 2187.460 1.630 2190.110 1.770 ;
        RECT 2189.550 -4.800 2190.110 1.630 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 877.290 50.220 877.610 50.280 ;
        RECT 2201.630 50.220 2201.950 50.280 ;
        RECT 877.290 50.080 2201.950 50.220 ;
        RECT 877.290 50.020 877.610 50.080 ;
        RECT 2201.630 50.020 2201.950 50.080 ;
        RECT 2201.630 16.560 2201.950 16.620 ;
        RECT 2207.610 16.560 2207.930 16.620 ;
        RECT 2201.630 16.420 2207.930 16.560 ;
        RECT 2201.630 16.360 2201.950 16.420 ;
        RECT 2207.610 16.360 2207.930 16.420 ;
      LAYER via ;
        RECT 877.320 50.020 877.580 50.280 ;
        RECT 2201.660 50.020 2201.920 50.280 ;
        RECT 2201.660 16.360 2201.920 16.620 ;
        RECT 2207.640 16.360 2207.900 16.620 ;
      LAYER met2 ;
        RECT 877.210 400.180 877.490 404.000 ;
        RECT 877.210 400.000 877.520 400.180 ;
        RECT 877.380 50.310 877.520 400.000 ;
        RECT 877.320 49.990 877.580 50.310 ;
        RECT 2201.660 49.990 2201.920 50.310 ;
        RECT 2201.720 16.650 2201.860 49.990 ;
        RECT 2201.660 16.330 2201.920 16.650 ;
        RECT 2207.640 16.330 2207.900 16.650 ;
        RECT 2207.700 2.400 2207.840 16.330 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.230 32.200 435.550 32.260 ;
        RECT 771.030 32.200 771.350 32.260 ;
        RECT 435.230 32.060 771.350 32.200 ;
        RECT 435.230 32.000 435.550 32.060 ;
        RECT 771.030 32.000 771.350 32.060 ;
      LAYER via ;
        RECT 435.260 32.000 435.520 32.260 ;
        RECT 771.060 32.000 771.320 32.260 ;
      LAYER met2 ;
        RECT 436.070 400.250 436.350 404.000 ;
        RECT 435.320 400.110 436.350 400.250 ;
        RECT 435.320 32.290 435.460 400.110 ;
        RECT 436.070 400.000 436.350 400.110 ;
        RECT 435.260 31.970 435.520 32.290 ;
        RECT 771.060 31.970 771.320 32.290 ;
        RECT 771.120 2.400 771.260 31.970 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.830 375.940 877.150 376.000 ;
        RECT 881.430 375.940 881.750 376.000 ;
        RECT 876.830 375.800 881.750 375.940 ;
        RECT 876.830 375.740 877.150 375.800 ;
        RECT 881.430 375.740 881.750 375.800 ;
        RECT 876.830 50.560 877.150 50.620 ;
        RECT 2225.090 50.560 2225.410 50.620 ;
        RECT 876.830 50.420 2225.410 50.560 ;
        RECT 876.830 50.360 877.150 50.420 ;
        RECT 2225.090 50.360 2225.410 50.420 ;
      LAYER via ;
        RECT 876.860 375.740 877.120 376.000 ;
        RECT 881.460 375.740 881.720 376.000 ;
        RECT 876.860 50.360 877.120 50.620 ;
        RECT 2225.120 50.360 2225.380 50.620 ;
      LAYER met2 ;
        RECT 882.730 400.250 883.010 404.000 ;
        RECT 881.520 400.110 883.010 400.250 ;
        RECT 881.520 376.030 881.660 400.110 ;
        RECT 882.730 400.000 883.010 400.110 ;
        RECT 876.860 375.710 877.120 376.030 ;
        RECT 881.460 375.710 881.720 376.030 ;
        RECT 876.920 50.650 877.060 375.710 ;
        RECT 876.860 50.330 877.120 50.650 ;
        RECT 2225.120 50.330 2225.380 50.650 ;
        RECT 2225.180 2.400 2225.320 50.330 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.730 375.940 884.050 376.000 ;
        RECT 886.950 375.940 887.270 376.000 ;
        RECT 883.730 375.800 887.270 375.940 ;
        RECT 883.730 375.740 884.050 375.800 ;
        RECT 886.950 375.740 887.270 375.800 ;
        RECT 883.730 50.900 884.050 50.960 ;
        RECT 2243.030 50.900 2243.350 50.960 ;
        RECT 883.730 50.760 2243.350 50.900 ;
        RECT 883.730 50.700 884.050 50.760 ;
        RECT 2243.030 50.700 2243.350 50.760 ;
      LAYER via ;
        RECT 883.760 375.740 884.020 376.000 ;
        RECT 886.980 375.740 887.240 376.000 ;
        RECT 883.760 50.700 884.020 50.960 ;
        RECT 2243.060 50.700 2243.320 50.960 ;
      LAYER met2 ;
        RECT 888.250 400.250 888.530 404.000 ;
        RECT 887.040 400.110 888.530 400.250 ;
        RECT 887.040 376.030 887.180 400.110 ;
        RECT 888.250 400.000 888.530 400.110 ;
        RECT 883.760 375.710 884.020 376.030 ;
        RECT 886.980 375.710 887.240 376.030 ;
        RECT 883.820 50.990 883.960 375.710 ;
        RECT 883.760 50.670 884.020 50.990 ;
        RECT 2243.060 50.670 2243.320 50.990 ;
        RECT 2243.120 2.400 2243.260 50.670 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.630 376.280 890.950 376.340 ;
        RECT 892.470 376.280 892.790 376.340 ;
        RECT 890.630 376.140 892.790 376.280 ;
        RECT 890.630 376.080 890.950 376.140 ;
        RECT 892.470 376.080 892.790 376.140 ;
        RECT 890.630 51.240 890.950 51.300 ;
        RECT 2258.210 51.240 2258.530 51.300 ;
        RECT 890.630 51.100 2258.530 51.240 ;
        RECT 890.630 51.040 890.950 51.100 ;
        RECT 2258.210 51.040 2258.530 51.100 ;
      LAYER via ;
        RECT 890.660 376.080 890.920 376.340 ;
        RECT 892.500 376.080 892.760 376.340 ;
        RECT 890.660 51.040 890.920 51.300 ;
        RECT 2258.240 51.040 2258.500 51.300 ;
      LAYER met2 ;
        RECT 893.770 400.250 894.050 404.000 ;
        RECT 892.560 400.110 894.050 400.250 ;
        RECT 892.560 376.370 892.700 400.110 ;
        RECT 893.770 400.000 894.050 400.110 ;
        RECT 890.660 376.050 890.920 376.370 ;
        RECT 892.500 376.050 892.760 376.370 ;
        RECT 890.720 51.330 890.860 376.050 ;
        RECT 890.660 51.010 890.920 51.330 ;
        RECT 2258.240 51.010 2258.500 51.330 ;
        RECT 2258.300 1.770 2258.440 51.010 ;
        RECT 2260.390 1.770 2260.950 2.400 ;
        RECT 2258.300 1.630 2260.950 1.770 ;
        RECT 2260.390 -4.800 2260.950 1.630 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.990 54.980 898.310 55.040 ;
        RECT 2278.450 54.980 2278.770 55.040 ;
        RECT 897.990 54.840 2278.770 54.980 ;
        RECT 897.990 54.780 898.310 54.840 ;
        RECT 2278.450 54.780 2278.770 54.840 ;
      LAYER via ;
        RECT 898.020 54.780 898.280 55.040 ;
        RECT 2278.480 54.780 2278.740 55.040 ;
      LAYER met2 ;
        RECT 899.290 400.250 899.570 404.000 ;
        RECT 898.080 400.110 899.570 400.250 ;
        RECT 898.080 55.070 898.220 400.110 ;
        RECT 899.290 400.000 899.570 400.110 ;
        RECT 898.020 54.750 898.280 55.070 ;
        RECT 2278.480 54.750 2278.740 55.070 ;
        RECT 2278.540 2.400 2278.680 54.750 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.890 54.640 905.210 54.700 ;
        RECT 2295.930 54.640 2296.250 54.700 ;
        RECT 904.890 54.500 2296.250 54.640 ;
        RECT 904.890 54.440 905.210 54.500 ;
        RECT 2295.930 54.440 2296.250 54.500 ;
      LAYER via ;
        RECT 904.920 54.440 905.180 54.700 ;
        RECT 2295.960 54.440 2296.220 54.700 ;
      LAYER met2 ;
        RECT 904.350 400.250 904.630 404.000 ;
        RECT 904.350 400.110 905.120 400.250 ;
        RECT 904.350 400.000 904.630 400.110 ;
        RECT 904.980 54.730 905.120 400.110 ;
        RECT 904.920 54.410 905.180 54.730 ;
        RECT 2295.960 54.410 2296.220 54.730 ;
        RECT 2296.020 2.400 2296.160 54.410 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 904.430 375.940 904.750 376.000 ;
        RECT 908.570 375.940 908.890 376.000 ;
        RECT 904.430 375.800 908.890 375.940 ;
        RECT 904.430 375.740 904.750 375.800 ;
        RECT 908.570 375.740 908.890 375.800 ;
        RECT 904.430 54.300 904.750 54.360 ;
        RECT 2311.570 54.300 2311.890 54.360 ;
        RECT 904.430 54.160 2311.890 54.300 ;
        RECT 904.430 54.100 904.750 54.160 ;
        RECT 2311.570 54.100 2311.890 54.160 ;
      LAYER via ;
        RECT 904.460 375.740 904.720 376.000 ;
        RECT 908.600 375.740 908.860 376.000 ;
        RECT 904.460 54.100 904.720 54.360 ;
        RECT 2311.600 54.100 2311.860 54.360 ;
      LAYER met2 ;
        RECT 909.870 400.250 910.150 404.000 ;
        RECT 908.660 400.110 910.150 400.250 ;
        RECT 908.660 376.030 908.800 400.110 ;
        RECT 909.870 400.000 910.150 400.110 ;
        RECT 904.460 375.710 904.720 376.030 ;
        RECT 908.600 375.710 908.860 376.030 ;
        RECT 904.520 54.390 904.660 375.710 ;
        RECT 904.460 54.070 904.720 54.390 ;
        RECT 2311.600 54.070 2311.860 54.390 ;
        RECT 2311.660 1.770 2311.800 54.070 ;
        RECT 2313.750 1.770 2314.310 2.400 ;
        RECT 2311.660 1.630 2314.310 1.770 ;
        RECT 2313.750 -4.800 2314.310 1.630 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.330 375.940 911.650 376.000 ;
        RECT 914.090 375.940 914.410 376.000 ;
        RECT 911.330 375.800 914.410 375.940 ;
        RECT 911.330 375.740 911.650 375.800 ;
        RECT 914.090 375.740 914.410 375.800 ;
        RECT 911.330 53.960 911.650 54.020 ;
        RECT 2329.050 53.960 2329.370 54.020 ;
        RECT 911.330 53.820 2329.370 53.960 ;
        RECT 911.330 53.760 911.650 53.820 ;
        RECT 2329.050 53.760 2329.370 53.820 ;
      LAYER via ;
        RECT 911.360 375.740 911.620 376.000 ;
        RECT 914.120 375.740 914.380 376.000 ;
        RECT 911.360 53.760 911.620 54.020 ;
        RECT 2329.080 53.760 2329.340 54.020 ;
      LAYER met2 ;
        RECT 915.390 400.250 915.670 404.000 ;
        RECT 914.180 400.110 915.670 400.250 ;
        RECT 914.180 376.030 914.320 400.110 ;
        RECT 915.390 400.000 915.670 400.110 ;
        RECT 911.360 375.710 911.620 376.030 ;
        RECT 914.120 375.710 914.380 376.030 ;
        RECT 911.420 54.050 911.560 375.710 ;
        RECT 911.360 53.730 911.620 54.050 ;
        RECT 2329.080 53.730 2329.340 54.050 ;
        RECT 2329.140 1.770 2329.280 53.730 ;
        RECT 2331.230 1.770 2331.790 2.400 ;
        RECT 2329.140 1.630 2331.790 1.770 ;
        RECT 2331.230 -4.800 2331.790 1.630 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.230 53.620 918.550 53.680 ;
        RECT 2349.290 53.620 2349.610 53.680 ;
        RECT 918.230 53.480 2349.610 53.620 ;
        RECT 918.230 53.420 918.550 53.480 ;
        RECT 2349.290 53.420 2349.610 53.480 ;
      LAYER via ;
        RECT 918.260 53.420 918.520 53.680 ;
        RECT 2349.320 53.420 2349.580 53.680 ;
      LAYER met2 ;
        RECT 920.910 400.250 921.190 404.000 ;
        RECT 919.700 400.110 921.190 400.250 ;
        RECT 919.700 351.970 919.840 400.110 ;
        RECT 920.910 400.000 921.190 400.110 ;
        RECT 918.320 351.830 919.840 351.970 ;
        RECT 918.320 53.710 918.460 351.830 ;
        RECT 918.260 53.390 918.520 53.710 ;
        RECT 2349.320 53.390 2349.580 53.710 ;
        RECT 2349.380 2.400 2349.520 53.390 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.590 53.280 925.910 53.340 ;
        RECT 2367.230 53.280 2367.550 53.340 ;
        RECT 925.590 53.140 2367.550 53.280 ;
        RECT 925.590 53.080 925.910 53.140 ;
        RECT 2367.230 53.080 2367.550 53.140 ;
      LAYER via ;
        RECT 925.620 53.080 925.880 53.340 ;
        RECT 2367.260 53.080 2367.520 53.340 ;
      LAYER met2 ;
        RECT 926.430 400.250 926.710 404.000 ;
        RECT 925.680 400.110 926.710 400.250 ;
        RECT 925.680 53.370 925.820 400.110 ;
        RECT 926.430 400.000 926.710 400.110 ;
        RECT 925.620 53.050 925.880 53.370 ;
        RECT 2367.260 53.050 2367.520 53.370 ;
        RECT 2367.320 2.400 2367.460 53.050 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.030 52.940 932.350 53.000 ;
        RECT 2382.410 52.940 2382.730 53.000 ;
        RECT 932.030 52.800 2382.730 52.940 ;
        RECT 932.030 52.740 932.350 52.800 ;
        RECT 2382.410 52.740 2382.730 52.800 ;
      LAYER via ;
        RECT 932.060 52.740 932.320 53.000 ;
        RECT 2382.440 52.740 2382.700 53.000 ;
      LAYER met2 ;
        RECT 931.950 400.180 932.230 404.000 ;
        RECT 931.950 400.000 932.260 400.180 ;
        RECT 932.120 53.030 932.260 400.000 ;
        RECT 932.060 52.710 932.320 53.030 ;
        RECT 2382.440 52.710 2382.700 53.030 ;
        RECT 2382.500 1.770 2382.640 52.710 ;
        RECT 2384.590 1.770 2385.150 2.400 ;
        RECT 2382.500 1.630 2385.150 1.770 ;
        RECT 2384.590 -4.800 2385.150 1.630 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 442.590 31.520 442.910 31.580 ;
        RECT 788.970 31.520 789.290 31.580 ;
        RECT 442.590 31.380 789.290 31.520 ;
        RECT 442.590 31.320 442.910 31.380 ;
        RECT 788.970 31.320 789.290 31.380 ;
      LAYER via ;
        RECT 442.620 31.320 442.880 31.580 ;
        RECT 789.000 31.320 789.260 31.580 ;
      LAYER met2 ;
        RECT 441.590 400.250 441.870 404.000 ;
        RECT 441.590 400.110 442.820 400.250 ;
        RECT 441.590 400.000 441.870 400.110 ;
        RECT 442.680 31.610 442.820 400.110 ;
        RECT 442.620 31.290 442.880 31.610 ;
        RECT 789.000 31.290 789.260 31.610 ;
        RECT 789.060 2.400 789.200 31.290 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.290 29.480 394.610 29.540 ;
        RECT 634.870 29.480 635.190 29.540 ;
        RECT 394.290 29.340 635.190 29.480 ;
        RECT 394.290 29.280 394.610 29.340 ;
        RECT 634.870 29.280 635.190 29.340 ;
      LAYER via ;
        RECT 394.320 29.280 394.580 29.540 ;
        RECT 634.900 29.280 635.160 29.540 ;
      LAYER met2 ;
        RECT 394.670 400.250 394.950 404.000 ;
        RECT 394.380 400.110 394.950 400.250 ;
        RECT 394.380 29.570 394.520 400.110 ;
        RECT 394.670 400.000 394.950 400.110 ;
        RECT 394.320 29.250 394.580 29.570 ;
        RECT 634.900 29.250 635.160 29.570 ;
        RECT 634.960 2.400 635.100 29.250 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.470 52.600 938.790 52.660 ;
        RECT 2408.630 52.600 2408.950 52.660 ;
        RECT 938.470 52.460 2408.950 52.600 ;
        RECT 938.470 52.400 938.790 52.460 ;
        RECT 2408.630 52.400 2408.950 52.460 ;
      LAYER via ;
        RECT 938.500 52.400 938.760 52.660 ;
        RECT 2408.660 52.400 2408.920 52.660 ;
      LAYER met2 ;
        RECT 938.850 400.250 939.130 404.000 ;
        RECT 938.560 400.110 939.130 400.250 ;
        RECT 938.560 52.690 938.700 400.110 ;
        RECT 938.850 400.000 939.130 400.110 ;
        RECT 938.500 52.370 938.760 52.690 ;
        RECT 2408.660 52.370 2408.920 52.690 ;
        RECT 2408.720 2.400 2408.860 52.370 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 938.930 386.480 939.250 386.540 ;
        RECT 943.070 386.480 943.390 386.540 ;
        RECT 938.930 386.340 943.390 386.480 ;
        RECT 938.930 386.280 939.250 386.340 ;
        RECT 943.070 386.280 943.390 386.340 ;
        RECT 938.930 52.260 939.250 52.320 ;
        RECT 2423.810 52.260 2424.130 52.320 ;
        RECT 938.930 52.120 2424.130 52.260 ;
        RECT 938.930 52.060 939.250 52.120 ;
        RECT 2423.810 52.060 2424.130 52.120 ;
      LAYER via ;
        RECT 938.960 386.280 939.220 386.540 ;
        RECT 943.100 386.280 943.360 386.540 ;
        RECT 938.960 52.060 939.220 52.320 ;
        RECT 2423.840 52.060 2424.100 52.320 ;
      LAYER met2 ;
        RECT 944.370 400.250 944.650 404.000 ;
        RECT 943.160 400.110 944.650 400.250 ;
        RECT 943.160 386.570 943.300 400.110 ;
        RECT 944.370 400.000 944.650 400.110 ;
        RECT 938.960 386.250 939.220 386.570 ;
        RECT 943.100 386.250 943.360 386.570 ;
        RECT 939.020 52.350 939.160 386.250 ;
        RECT 938.960 52.030 939.220 52.350 ;
        RECT 2423.840 52.030 2424.100 52.350 ;
        RECT 2423.900 1.770 2424.040 52.030 ;
        RECT 2425.990 1.770 2426.550 2.400 ;
        RECT 2423.900 1.630 2426.550 1.770 ;
        RECT 2425.990 -4.800 2426.550 1.630 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.370 386.480 945.690 386.540 ;
        RECT 948.590 386.480 948.910 386.540 ;
        RECT 945.370 386.340 948.910 386.480 ;
        RECT 945.370 386.280 945.690 386.340 ;
        RECT 948.590 386.280 948.910 386.340 ;
        RECT 945.370 51.920 945.690 51.980 ;
        RECT 2444.050 51.920 2444.370 51.980 ;
        RECT 945.370 51.780 2444.370 51.920 ;
        RECT 945.370 51.720 945.690 51.780 ;
        RECT 2444.050 51.720 2444.370 51.780 ;
      LAYER via ;
        RECT 945.400 386.280 945.660 386.540 ;
        RECT 948.620 386.280 948.880 386.540 ;
        RECT 945.400 51.720 945.660 51.980 ;
        RECT 2444.080 51.720 2444.340 51.980 ;
      LAYER met2 ;
        RECT 949.890 400.250 950.170 404.000 ;
        RECT 948.680 400.110 950.170 400.250 ;
        RECT 948.680 386.570 948.820 400.110 ;
        RECT 949.890 400.000 950.170 400.110 ;
        RECT 945.400 386.250 945.660 386.570 ;
        RECT 948.620 386.250 948.880 386.570 ;
        RECT 945.460 52.010 945.600 386.250 ;
        RECT 945.400 51.690 945.660 52.010 ;
        RECT 2444.080 51.690 2444.340 52.010 ;
        RECT 2444.140 2.400 2444.280 51.690 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.270 386.480 952.590 386.540 ;
        RECT 954.110 386.480 954.430 386.540 ;
        RECT 952.270 386.340 954.430 386.480 ;
        RECT 952.270 386.280 952.590 386.340 ;
        RECT 954.110 386.280 954.430 386.340 ;
      LAYER via ;
        RECT 952.300 386.280 952.560 386.540 ;
        RECT 954.140 386.280 954.400 386.540 ;
      LAYER met2 ;
        RECT 955.410 400.250 955.690 404.000 ;
        RECT 954.200 400.110 955.690 400.250 ;
        RECT 954.200 386.570 954.340 400.110 ;
        RECT 955.410 400.000 955.690 400.110 ;
        RECT 952.300 386.250 952.560 386.570 ;
        RECT 954.140 386.250 954.400 386.570 ;
        RECT 952.360 52.205 952.500 386.250 ;
        RECT 952.290 51.835 952.570 52.205 ;
        RECT 2461.550 51.835 2461.830 52.205 ;
        RECT 2461.620 2.400 2461.760 51.835 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
      LAYER via2 ;
        RECT 952.290 51.880 952.570 52.160 ;
        RECT 2461.550 51.880 2461.830 52.160 ;
      LAYER met3 ;
        RECT 952.265 52.170 952.595 52.185 ;
        RECT 2461.525 52.170 2461.855 52.185 ;
        RECT 952.265 51.870 2461.855 52.170 ;
        RECT 952.265 51.855 952.595 51.870 ;
        RECT 2461.525 51.855 2461.855 51.870 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.090 51.580 960.410 51.640 ;
        RECT 2477.170 51.580 2477.490 51.640 ;
        RECT 960.090 51.440 2477.490 51.580 ;
        RECT 960.090 51.380 960.410 51.440 ;
        RECT 2477.170 51.380 2477.490 51.440 ;
      LAYER via ;
        RECT 960.120 51.380 960.380 51.640 ;
        RECT 2477.200 51.380 2477.460 51.640 ;
      LAYER met2 ;
        RECT 960.930 400.250 961.210 404.000 ;
        RECT 960.180 400.110 961.210 400.250 ;
        RECT 960.180 51.670 960.320 400.110 ;
        RECT 960.930 400.000 961.210 400.110 ;
        RECT 960.120 51.350 960.380 51.670 ;
        RECT 2477.200 51.350 2477.460 51.670 ;
        RECT 2477.260 1.770 2477.400 51.350 ;
        RECT 2479.350 1.770 2479.910 2.400 ;
        RECT 2477.260 1.630 2479.910 1.770 ;
        RECT 2479.350 -4.800 2479.910 1.630 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.450 400.180 966.730 404.000 ;
        RECT 966.450 400.000 966.760 400.180 ;
        RECT 966.620 51.525 966.760 400.000 ;
        RECT 966.550 51.155 966.830 51.525 ;
        RECT 2494.670 51.155 2494.950 51.525 ;
        RECT 2494.740 1.770 2494.880 51.155 ;
        RECT 2496.830 1.770 2497.390 2.400 ;
        RECT 2494.740 1.630 2497.390 1.770 ;
        RECT 2496.830 -4.800 2497.390 1.630 ;
      LAYER via2 ;
        RECT 966.550 51.200 966.830 51.480 ;
        RECT 2494.670 51.200 2494.950 51.480 ;
      LAYER met3 ;
        RECT 966.525 51.490 966.855 51.505 ;
        RECT 2494.645 51.490 2494.975 51.505 ;
        RECT 966.525 51.190 2494.975 51.490 ;
        RECT 966.525 51.175 966.855 51.190 ;
        RECT 2494.645 51.175 2494.975 51.190 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 967.450 114.820 967.770 114.880 ;
        RECT 2511.670 114.820 2511.990 114.880 ;
        RECT 967.450 114.680 2511.990 114.820 ;
        RECT 967.450 114.620 967.770 114.680 ;
        RECT 2511.670 114.620 2511.990 114.680 ;
      LAYER via ;
        RECT 967.480 114.620 967.740 114.880 ;
        RECT 2511.700 114.620 2511.960 114.880 ;
      LAYER met2 ;
        RECT 971.510 400.250 971.790 404.000 ;
        RECT 970.300 400.110 971.790 400.250 ;
        RECT 970.300 324.370 970.440 400.110 ;
        RECT 971.510 400.000 971.790 400.110 ;
        RECT 967.540 324.230 970.440 324.370 ;
        RECT 967.540 114.910 967.680 324.230 ;
        RECT 967.480 114.590 967.740 114.910 ;
        RECT 2511.700 114.590 2511.960 114.910 ;
        RECT 2511.760 82.870 2511.900 114.590 ;
        RECT 2511.760 82.730 2515.120 82.870 ;
        RECT 2514.980 2.400 2515.120 82.730 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 974.350 114.480 974.670 114.540 ;
        RECT 2532.370 114.480 2532.690 114.540 ;
        RECT 974.350 114.340 2532.690 114.480 ;
        RECT 974.350 114.280 974.670 114.340 ;
        RECT 2532.370 114.280 2532.690 114.340 ;
      LAYER via ;
        RECT 974.380 114.280 974.640 114.540 ;
        RECT 2532.400 114.280 2532.660 114.540 ;
      LAYER met2 ;
        RECT 977.030 400.250 977.310 404.000 ;
        RECT 975.820 400.110 977.310 400.250 ;
        RECT 975.820 324.370 975.960 400.110 ;
        RECT 977.030 400.000 977.310 400.110 ;
        RECT 974.440 324.230 975.960 324.370 ;
        RECT 974.440 114.570 974.580 324.230 ;
        RECT 974.380 114.250 974.640 114.570 ;
        RECT 2532.400 114.250 2532.660 114.570 ;
        RECT 2532.460 2.400 2532.600 114.250 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 981.250 114.140 981.570 114.200 ;
        RECT 2546.170 114.140 2546.490 114.200 ;
        RECT 981.250 114.000 2546.490 114.140 ;
        RECT 981.250 113.940 981.570 114.000 ;
        RECT 2546.170 113.940 2546.490 114.000 ;
      LAYER via ;
        RECT 981.280 113.940 981.540 114.200 ;
        RECT 2546.200 113.940 2546.460 114.200 ;
      LAYER met2 ;
        RECT 982.550 400.250 982.830 404.000 ;
        RECT 981.340 400.110 982.830 400.250 ;
        RECT 981.340 114.230 981.480 400.110 ;
        RECT 982.550 400.000 982.830 400.110 ;
        RECT 981.280 113.910 981.540 114.230 ;
        RECT 2546.200 113.910 2546.460 114.230 ;
        RECT 2546.260 82.870 2546.400 113.910 ;
        RECT 2546.260 82.730 2548.240 82.870 ;
        RECT 2548.100 1.770 2548.240 82.730 ;
        RECT 2550.190 1.770 2550.750 2.400 ;
        RECT 2548.100 1.630 2550.750 1.770 ;
        RECT 2550.190 -4.800 2550.750 1.630 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.690 113.800 988.010 113.860 ;
        RECT 2566.870 113.800 2567.190 113.860 ;
        RECT 987.690 113.660 2567.190 113.800 ;
        RECT 987.690 113.600 988.010 113.660 ;
        RECT 2566.870 113.600 2567.190 113.660 ;
      LAYER via ;
        RECT 987.720 113.600 987.980 113.860 ;
        RECT 2566.900 113.600 2567.160 113.860 ;
      LAYER met2 ;
        RECT 988.070 400.250 988.350 404.000 ;
        RECT 987.780 400.110 988.350 400.250 ;
        RECT 987.780 113.890 987.920 400.110 ;
        RECT 988.070 400.000 988.350 400.110 ;
        RECT 987.720 113.570 987.980 113.890 ;
        RECT 2566.900 113.570 2567.160 113.890 ;
        RECT 2566.960 1.770 2567.100 113.570 ;
        RECT 2567.670 1.770 2568.230 2.400 ;
        RECT 2566.960 1.630 2568.230 1.770 ;
        RECT 2567.670 -4.800 2568.230 1.630 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.030 31.180 449.350 31.240 ;
        RECT 812.430 31.180 812.750 31.240 ;
        RECT 449.030 31.040 812.750 31.180 ;
        RECT 449.030 30.980 449.350 31.040 ;
        RECT 812.430 30.980 812.750 31.040 ;
      LAYER via ;
        RECT 449.060 30.980 449.320 31.240 ;
        RECT 812.460 30.980 812.720 31.240 ;
      LAYER met2 ;
        RECT 448.950 400.180 449.230 404.000 ;
        RECT 448.950 400.000 449.260 400.180 ;
        RECT 449.120 31.270 449.260 400.000 ;
        RECT 449.060 30.950 449.320 31.270 ;
        RECT 812.460 30.950 812.720 31.270 ;
        RECT 812.520 2.400 812.660 30.950 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.590 400.930 993.870 404.000 ;
        RECT 993.590 400.790 995.280 400.930 ;
        RECT 993.590 400.000 993.870 400.790 ;
        RECT 995.140 113.405 995.280 400.790 ;
        RECT 995.070 113.035 995.350 113.405 ;
        RECT 2580.690 113.035 2580.970 113.405 ;
        RECT 2580.760 82.870 2580.900 113.035 ;
        RECT 2580.760 82.730 2585.960 82.870 ;
        RECT 2585.820 2.400 2585.960 82.730 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
      LAYER via2 ;
        RECT 995.070 113.080 995.350 113.360 ;
        RECT 2580.690 113.080 2580.970 113.360 ;
      LAYER met3 ;
        RECT 995.045 113.370 995.375 113.385 ;
        RECT 2580.665 113.370 2580.995 113.385 ;
        RECT 995.045 113.070 2580.995 113.370 ;
        RECT 995.045 113.055 995.375 113.070 ;
        RECT 2580.665 113.055 2580.995 113.070 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.130 386.480 994.450 386.540 ;
        RECT 997.810 386.480 998.130 386.540 ;
        RECT 994.130 386.340 998.130 386.480 ;
        RECT 994.130 386.280 994.450 386.340 ;
        RECT 997.810 386.280 998.130 386.340 ;
        RECT 994.130 57.360 994.450 57.420 ;
        RECT 2601.370 57.360 2601.690 57.420 ;
        RECT 994.130 57.220 2601.690 57.360 ;
        RECT 994.130 57.160 994.450 57.220 ;
        RECT 2601.370 57.160 2601.690 57.220 ;
      LAYER via ;
        RECT 994.160 386.280 994.420 386.540 ;
        RECT 997.840 386.280 998.100 386.540 ;
        RECT 994.160 57.160 994.420 57.420 ;
        RECT 2601.400 57.160 2601.660 57.420 ;
      LAYER met2 ;
        RECT 999.110 400.250 999.390 404.000 ;
        RECT 997.900 400.110 999.390 400.250 ;
        RECT 997.900 386.570 998.040 400.110 ;
        RECT 999.110 400.000 999.390 400.110 ;
        RECT 994.160 386.250 994.420 386.570 ;
        RECT 997.840 386.250 998.100 386.570 ;
        RECT 994.220 57.450 994.360 386.250 ;
        RECT 994.160 57.130 994.420 57.450 ;
        RECT 2601.400 57.130 2601.660 57.450 ;
        RECT 2601.460 1.770 2601.600 57.130 ;
        RECT 2603.550 1.770 2604.110 2.400 ;
        RECT 2601.460 1.630 2604.110 1.770 ;
        RECT 2603.550 -4.800 2604.110 1.630 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.030 386.480 1001.350 386.540 ;
        RECT 1002.870 386.480 1003.190 386.540 ;
        RECT 1001.030 386.340 1003.190 386.480 ;
        RECT 1001.030 386.280 1001.350 386.340 ;
        RECT 1002.870 386.280 1003.190 386.340 ;
        RECT 1001.030 57.700 1001.350 57.760 ;
        RECT 2618.850 57.700 2619.170 57.760 ;
        RECT 1001.030 57.560 2619.170 57.700 ;
        RECT 1001.030 57.500 1001.350 57.560 ;
        RECT 2618.850 57.500 2619.170 57.560 ;
      LAYER via ;
        RECT 1001.060 386.280 1001.320 386.540 ;
        RECT 1002.900 386.280 1003.160 386.540 ;
        RECT 1001.060 57.500 1001.320 57.760 ;
        RECT 2618.880 57.500 2619.140 57.760 ;
      LAYER met2 ;
        RECT 1004.170 400.250 1004.450 404.000 ;
        RECT 1002.960 400.110 1004.450 400.250 ;
        RECT 1002.960 386.570 1003.100 400.110 ;
        RECT 1004.170 400.000 1004.450 400.110 ;
        RECT 1001.060 386.250 1001.320 386.570 ;
        RECT 1002.900 386.250 1003.160 386.570 ;
        RECT 1001.120 57.790 1001.260 386.250 ;
        RECT 1001.060 57.470 1001.320 57.790 ;
        RECT 2618.880 57.470 2619.140 57.790 ;
        RECT 2618.940 1.770 2619.080 57.470 ;
        RECT 2621.030 1.770 2621.590 2.400 ;
        RECT 2618.940 1.630 2621.590 1.770 ;
        RECT 2621.030 -4.800 2621.590 1.630 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1008.390 58.040 1008.710 58.100 ;
        RECT 2639.090 58.040 2639.410 58.100 ;
        RECT 1008.390 57.900 2639.410 58.040 ;
        RECT 1008.390 57.840 1008.710 57.900 ;
        RECT 2639.090 57.840 2639.410 57.900 ;
      LAYER via ;
        RECT 1008.420 57.840 1008.680 58.100 ;
        RECT 2639.120 57.840 2639.380 58.100 ;
      LAYER met2 ;
        RECT 1009.690 400.250 1009.970 404.000 ;
        RECT 1008.480 400.110 1009.970 400.250 ;
        RECT 1008.480 58.130 1008.620 400.110 ;
        RECT 1009.690 400.000 1009.970 400.110 ;
        RECT 1008.420 57.810 1008.680 58.130 ;
        RECT 2639.120 57.810 2639.380 58.130 ;
        RECT 2639.180 2.400 2639.320 57.810 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1014.830 58.380 1015.150 58.440 ;
        RECT 2657.030 58.380 2657.350 58.440 ;
        RECT 1014.830 58.240 2657.350 58.380 ;
        RECT 1014.830 58.180 1015.150 58.240 ;
        RECT 2657.030 58.180 2657.350 58.240 ;
      LAYER via ;
        RECT 1014.860 58.180 1015.120 58.440 ;
        RECT 2657.060 58.180 2657.320 58.440 ;
      LAYER met2 ;
        RECT 1015.210 400.250 1015.490 404.000 ;
        RECT 1014.920 400.110 1015.490 400.250 ;
        RECT 1014.920 58.470 1015.060 400.110 ;
        RECT 1015.210 400.000 1015.490 400.110 ;
        RECT 1014.860 58.150 1015.120 58.470 ;
        RECT 2657.060 58.150 2657.320 58.470 ;
        RECT 2657.120 16.730 2657.260 58.150 ;
        RECT 2656.660 16.590 2657.260 16.730 ;
        RECT 2656.660 2.400 2656.800 16.590 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1015.290 386.480 1015.610 386.540 ;
        RECT 1019.430 386.480 1019.750 386.540 ;
        RECT 1015.290 386.340 1019.750 386.480 ;
        RECT 1015.290 386.280 1015.610 386.340 ;
        RECT 1019.430 386.280 1019.750 386.340 ;
        RECT 1015.290 62.120 1015.610 62.180 ;
        RECT 2672.210 62.120 2672.530 62.180 ;
        RECT 1015.290 61.980 2672.530 62.120 ;
        RECT 1015.290 61.920 1015.610 61.980 ;
        RECT 2672.210 61.920 2672.530 61.980 ;
      LAYER via ;
        RECT 1015.320 386.280 1015.580 386.540 ;
        RECT 1019.460 386.280 1019.720 386.540 ;
        RECT 1015.320 61.920 1015.580 62.180 ;
        RECT 2672.240 61.920 2672.500 62.180 ;
      LAYER met2 ;
        RECT 1020.730 400.250 1021.010 404.000 ;
        RECT 1019.520 400.110 1021.010 400.250 ;
        RECT 1019.520 386.570 1019.660 400.110 ;
        RECT 1020.730 400.000 1021.010 400.110 ;
        RECT 1015.320 386.250 1015.580 386.570 ;
        RECT 1019.460 386.250 1019.720 386.570 ;
        RECT 1015.380 62.210 1015.520 386.250 ;
        RECT 1015.320 61.890 1015.580 62.210 ;
        RECT 2672.240 61.890 2672.500 62.210 ;
        RECT 2672.300 1.770 2672.440 61.890 ;
        RECT 2674.390 1.770 2674.950 2.400 ;
        RECT 2672.300 1.630 2674.950 1.770 ;
        RECT 2674.390 -4.800 2674.950 1.630 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1021.730 385.800 1022.050 385.860 ;
        RECT 1024.950 385.800 1025.270 385.860 ;
        RECT 1021.730 385.660 1025.270 385.800 ;
        RECT 1021.730 385.600 1022.050 385.660 ;
        RECT 1024.950 385.600 1025.270 385.660 ;
        RECT 1021.730 61.780 1022.050 61.840 ;
        RECT 2691.070 61.780 2691.390 61.840 ;
        RECT 1021.730 61.640 2691.390 61.780 ;
        RECT 1021.730 61.580 1022.050 61.640 ;
        RECT 2691.070 61.580 2691.390 61.640 ;
      LAYER via ;
        RECT 1021.760 385.600 1022.020 385.860 ;
        RECT 1024.980 385.600 1025.240 385.860 ;
        RECT 1021.760 61.580 1022.020 61.840 ;
        RECT 2691.100 61.580 2691.360 61.840 ;
      LAYER met2 ;
        RECT 1026.250 400.250 1026.530 404.000 ;
        RECT 1025.040 400.110 1026.530 400.250 ;
        RECT 1025.040 385.890 1025.180 400.110 ;
        RECT 1026.250 400.000 1026.530 400.110 ;
        RECT 1021.760 385.570 1022.020 385.890 ;
        RECT 1024.980 385.570 1025.240 385.890 ;
        RECT 1021.820 61.870 1021.960 385.570 ;
        RECT 1021.760 61.550 1022.020 61.870 ;
        RECT 2691.100 61.550 2691.360 61.870 ;
        RECT 2691.160 1.770 2691.300 61.550 ;
        RECT 2691.870 1.770 2692.430 2.400 ;
        RECT 2691.160 1.630 2692.430 1.770 ;
        RECT 2691.870 -4.800 2692.430 1.630 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1028.630 61.440 1028.950 61.500 ;
        RECT 2709.930 61.440 2710.250 61.500 ;
        RECT 1028.630 61.300 2710.250 61.440 ;
        RECT 1028.630 61.240 1028.950 61.300 ;
        RECT 2709.930 61.240 2710.250 61.300 ;
      LAYER via ;
        RECT 1028.660 61.240 1028.920 61.500 ;
        RECT 2709.960 61.240 2710.220 61.500 ;
      LAYER met2 ;
        RECT 1031.770 400.250 1032.050 404.000 ;
        RECT 1030.560 400.110 1032.050 400.250 ;
        RECT 1030.560 387.330 1030.700 400.110 ;
        RECT 1031.770 400.000 1032.050 400.110 ;
        RECT 1028.720 387.190 1030.700 387.330 ;
        RECT 1028.720 61.530 1028.860 387.190 ;
        RECT 1028.660 61.210 1028.920 61.530 ;
        RECT 2709.960 61.210 2710.220 61.530 ;
        RECT 2710.020 2.400 2710.160 61.210 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.990 61.100 1036.310 61.160 ;
        RECT 2727.410 61.100 2727.730 61.160 ;
        RECT 1035.990 60.960 2727.730 61.100 ;
        RECT 1035.990 60.900 1036.310 60.960 ;
        RECT 2727.410 60.900 2727.730 60.960 ;
      LAYER via ;
        RECT 1036.020 60.900 1036.280 61.160 ;
        RECT 2727.440 60.900 2727.700 61.160 ;
      LAYER met2 ;
        RECT 1036.830 400.250 1037.110 404.000 ;
        RECT 1036.080 400.110 1037.110 400.250 ;
        RECT 1036.080 61.190 1036.220 400.110 ;
        RECT 1036.830 400.000 1037.110 400.110 ;
        RECT 1036.020 60.870 1036.280 61.190 ;
        RECT 2727.440 60.870 2727.700 61.190 ;
        RECT 2727.500 2.400 2727.640 60.870 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.890 60.760 1043.210 60.820 ;
        RECT 2743.050 60.760 2743.370 60.820 ;
        RECT 1042.890 60.620 2743.370 60.760 ;
        RECT 1042.890 60.560 1043.210 60.620 ;
        RECT 2743.050 60.560 2743.370 60.620 ;
      LAYER via ;
        RECT 1042.920 60.560 1043.180 60.820 ;
        RECT 2743.080 60.560 2743.340 60.820 ;
      LAYER met2 ;
        RECT 1042.350 400.250 1042.630 404.000 ;
        RECT 1042.350 400.110 1043.120 400.250 ;
        RECT 1042.350 400.000 1042.630 400.110 ;
        RECT 1042.980 60.850 1043.120 400.110 ;
        RECT 1042.920 60.530 1043.180 60.850 ;
        RECT 2743.080 60.530 2743.340 60.850 ;
        RECT 2743.140 1.770 2743.280 60.530 ;
        RECT 2745.230 1.770 2745.790 2.400 ;
        RECT 2743.140 1.630 2745.790 1.770 ;
        RECT 2745.230 -4.800 2745.790 1.630 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 448.570 376.280 448.890 376.340 ;
        RECT 453.170 376.280 453.490 376.340 ;
        RECT 448.570 376.140 453.490 376.280 ;
        RECT 448.570 376.080 448.890 376.140 ;
        RECT 453.170 376.080 453.490 376.140 ;
        RECT 448.570 29.140 448.890 29.200 ;
        RECT 620.610 29.140 620.930 29.200 ;
        RECT 448.570 29.000 620.930 29.140 ;
        RECT 448.570 28.940 448.890 29.000 ;
        RECT 620.610 28.940 620.930 29.000 ;
        RECT 620.610 19.280 620.930 19.340 ;
        RECT 830.370 19.280 830.690 19.340 ;
        RECT 620.610 19.140 830.690 19.280 ;
        RECT 620.610 19.080 620.930 19.140 ;
        RECT 830.370 19.080 830.690 19.140 ;
      LAYER via ;
        RECT 448.600 376.080 448.860 376.340 ;
        RECT 453.200 376.080 453.460 376.340 ;
        RECT 448.600 28.940 448.860 29.200 ;
        RECT 620.640 28.940 620.900 29.200 ;
        RECT 620.640 19.080 620.900 19.340 ;
        RECT 830.400 19.080 830.660 19.340 ;
      LAYER met2 ;
        RECT 454.470 400.250 454.750 404.000 ;
        RECT 453.260 400.110 454.750 400.250 ;
        RECT 453.260 376.370 453.400 400.110 ;
        RECT 454.470 400.000 454.750 400.110 ;
        RECT 448.600 376.050 448.860 376.370 ;
        RECT 453.200 376.050 453.460 376.370 ;
        RECT 448.660 29.230 448.800 376.050 ;
        RECT 448.600 28.910 448.860 29.230 ;
        RECT 620.640 28.910 620.900 29.230 ;
        RECT 620.700 19.370 620.840 28.910 ;
        RECT 620.640 19.050 620.900 19.370 ;
        RECT 830.400 19.050 830.660 19.370 ;
        RECT 830.460 2.400 830.600 19.050 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1042.430 375.940 1042.750 376.000 ;
        RECT 1046.570 375.940 1046.890 376.000 ;
        RECT 1042.430 375.800 1046.890 375.940 ;
        RECT 1042.430 375.740 1042.750 375.800 ;
        RECT 1046.570 375.740 1046.890 375.800 ;
        RECT 1042.430 60.420 1042.750 60.480 ;
        RECT 2763.290 60.420 2763.610 60.480 ;
        RECT 1042.430 60.280 2763.610 60.420 ;
        RECT 1042.430 60.220 1042.750 60.280 ;
        RECT 2763.290 60.220 2763.610 60.280 ;
      LAYER via ;
        RECT 1042.460 375.740 1042.720 376.000 ;
        RECT 1046.600 375.740 1046.860 376.000 ;
        RECT 1042.460 60.220 1042.720 60.480 ;
        RECT 2763.320 60.220 2763.580 60.480 ;
      LAYER met2 ;
        RECT 1047.870 400.250 1048.150 404.000 ;
        RECT 1046.660 400.110 1048.150 400.250 ;
        RECT 1046.660 376.030 1046.800 400.110 ;
        RECT 1047.870 400.000 1048.150 400.110 ;
        RECT 1042.460 375.710 1042.720 376.030 ;
        RECT 1046.600 375.710 1046.860 376.030 ;
        RECT 1042.520 60.510 1042.660 375.710 ;
        RECT 1042.460 60.190 1042.720 60.510 ;
        RECT 2763.320 60.190 2763.580 60.510 ;
        RECT 2763.380 2.400 2763.520 60.190 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1048.870 376.280 1049.190 376.340 ;
        RECT 1052.090 376.280 1052.410 376.340 ;
        RECT 1048.870 376.140 1052.410 376.280 ;
        RECT 1048.870 376.080 1049.190 376.140 ;
        RECT 1052.090 376.080 1052.410 376.140 ;
        RECT 1048.870 60.080 1049.190 60.140 ;
        RECT 2781.230 60.080 2781.550 60.140 ;
        RECT 1048.870 59.940 2781.550 60.080 ;
        RECT 1048.870 59.880 1049.190 59.940 ;
        RECT 2781.230 59.880 2781.550 59.940 ;
      LAYER via ;
        RECT 1048.900 376.080 1049.160 376.340 ;
        RECT 1052.120 376.080 1052.380 376.340 ;
        RECT 1048.900 59.880 1049.160 60.140 ;
        RECT 2781.260 59.880 2781.520 60.140 ;
      LAYER met2 ;
        RECT 1053.390 400.250 1053.670 404.000 ;
        RECT 1052.180 400.110 1053.670 400.250 ;
        RECT 1052.180 376.370 1052.320 400.110 ;
        RECT 1053.390 400.000 1053.670 400.110 ;
        RECT 1048.900 376.050 1049.160 376.370 ;
        RECT 1052.120 376.050 1052.380 376.370 ;
        RECT 1048.960 60.170 1049.100 376.050 ;
        RECT 1048.900 59.850 1049.160 60.170 ;
        RECT 2781.260 59.850 2781.520 60.170 ;
        RECT 2781.320 16.730 2781.460 59.850 ;
        RECT 2780.860 16.590 2781.460 16.730 ;
        RECT 2780.860 2.400 2781.000 16.590 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1055.770 375.940 1056.090 376.000 ;
        RECT 1057.610 375.940 1057.930 376.000 ;
        RECT 1055.770 375.800 1057.930 375.940 ;
        RECT 1055.770 375.740 1056.090 375.800 ;
        RECT 1057.610 375.740 1057.930 375.800 ;
        RECT 1055.770 59.740 1056.090 59.800 ;
        RECT 2796.410 59.740 2796.730 59.800 ;
        RECT 1055.770 59.600 2796.730 59.740 ;
        RECT 1055.770 59.540 1056.090 59.600 ;
        RECT 2796.410 59.540 2796.730 59.600 ;
      LAYER via ;
        RECT 1055.800 375.740 1056.060 376.000 ;
        RECT 1057.640 375.740 1057.900 376.000 ;
        RECT 1055.800 59.540 1056.060 59.800 ;
        RECT 2796.440 59.540 2796.700 59.800 ;
      LAYER met2 ;
        RECT 1058.910 400.250 1059.190 404.000 ;
        RECT 1057.700 400.110 1059.190 400.250 ;
        RECT 1057.700 376.030 1057.840 400.110 ;
        RECT 1058.910 400.000 1059.190 400.110 ;
        RECT 1055.800 375.710 1056.060 376.030 ;
        RECT 1057.640 375.710 1057.900 376.030 ;
        RECT 1055.860 59.830 1056.000 375.710 ;
        RECT 1055.800 59.510 1056.060 59.830 ;
        RECT 2796.440 59.510 2796.700 59.830 ;
        RECT 2796.500 1.770 2796.640 59.510 ;
        RECT 2798.590 1.770 2799.150 2.400 ;
        RECT 2796.500 1.630 2799.150 1.770 ;
        RECT 2798.590 -4.800 2799.150 1.630 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1062.670 376.280 1062.990 376.340 ;
        RECT 1064.050 376.280 1064.370 376.340 ;
        RECT 1062.670 376.140 1064.370 376.280 ;
        RECT 1062.670 376.080 1062.990 376.140 ;
        RECT 1064.050 376.080 1064.370 376.140 ;
        RECT 1062.670 59.400 1062.990 59.460 ;
        RECT 2815.270 59.400 2815.590 59.460 ;
        RECT 1062.670 59.260 2815.590 59.400 ;
        RECT 1062.670 59.200 1062.990 59.260 ;
        RECT 2815.270 59.200 2815.590 59.260 ;
      LAYER via ;
        RECT 1062.700 376.080 1062.960 376.340 ;
        RECT 1064.080 376.080 1064.340 376.340 ;
        RECT 1062.700 59.200 1062.960 59.460 ;
        RECT 2815.300 59.200 2815.560 59.460 ;
      LAYER met2 ;
        RECT 1064.430 400.250 1064.710 404.000 ;
        RECT 1064.140 400.110 1064.710 400.250 ;
        RECT 1064.140 376.370 1064.280 400.110 ;
        RECT 1064.430 400.000 1064.710 400.110 ;
        RECT 1062.700 376.050 1062.960 376.370 ;
        RECT 1064.080 376.050 1064.340 376.370 ;
        RECT 1062.760 59.490 1062.900 376.050 ;
        RECT 1062.700 59.170 1062.960 59.490 ;
        RECT 2815.300 59.170 2815.560 59.490 ;
        RECT 2815.360 1.770 2815.500 59.170 ;
        RECT 2816.070 1.770 2816.630 2.400 ;
        RECT 2815.360 1.630 2816.630 1.770 ;
        RECT 2816.070 -4.800 2816.630 1.630 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.030 376.280 1070.350 376.340 ;
        RECT 1070.950 376.280 1071.270 376.340 ;
        RECT 1070.030 376.140 1071.270 376.280 ;
        RECT 1070.030 376.080 1070.350 376.140 ;
        RECT 1070.950 376.080 1071.270 376.140 ;
      LAYER via ;
        RECT 1070.060 376.080 1070.320 376.340 ;
        RECT 1070.980 376.080 1071.240 376.340 ;
      LAYER met2 ;
        RECT 1069.490 400.250 1069.770 404.000 ;
        RECT 1069.490 400.110 1070.260 400.250 ;
        RECT 1069.490 400.000 1069.770 400.110 ;
        RECT 1070.120 376.370 1070.260 400.110 ;
        RECT 1070.060 376.050 1070.320 376.370 ;
        RECT 1070.980 376.050 1071.240 376.370 ;
        RECT 1071.040 59.005 1071.180 376.050 ;
        RECT 1070.970 58.635 1071.250 59.005 ;
        RECT 2834.150 58.635 2834.430 59.005 ;
        RECT 2834.220 2.400 2834.360 58.635 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
      LAYER via2 ;
        RECT 1070.970 58.680 1071.250 58.960 ;
        RECT 2834.150 58.680 2834.430 58.960 ;
      LAYER met3 ;
        RECT 1070.945 58.970 1071.275 58.985 ;
        RECT 2834.125 58.970 2834.455 58.985 ;
        RECT 1070.945 58.670 2834.455 58.970 ;
        RECT 1070.945 58.655 1071.275 58.670 ;
        RECT 2834.125 58.655 2834.455 58.670 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.030 375.600 1070.350 375.660 ;
        RECT 1073.710 375.600 1074.030 375.660 ;
        RECT 1070.030 375.460 1074.030 375.600 ;
        RECT 1070.030 375.400 1070.350 375.460 ;
        RECT 1073.710 375.400 1074.030 375.460 ;
      LAYER via ;
        RECT 1070.060 375.400 1070.320 375.660 ;
        RECT 1073.740 375.400 1074.000 375.660 ;
      LAYER met2 ;
        RECT 1075.010 400.250 1075.290 404.000 ;
        RECT 1073.800 400.110 1075.290 400.250 ;
        RECT 1073.800 375.690 1073.940 400.110 ;
        RECT 1075.010 400.000 1075.290 400.110 ;
        RECT 1070.060 375.370 1070.320 375.690 ;
        RECT 1073.740 375.370 1074.000 375.690 ;
        RECT 1070.120 58.325 1070.260 375.370 ;
        RECT 1070.050 57.955 1070.330 58.325 ;
        RECT 2851.630 57.955 2851.910 58.325 ;
        RECT 2851.700 2.400 2851.840 57.955 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
      LAYER via2 ;
        RECT 1070.050 58.000 1070.330 58.280 ;
        RECT 2851.630 58.000 2851.910 58.280 ;
      LAYER met3 ;
        RECT 1070.025 58.290 1070.355 58.305 ;
        RECT 2851.605 58.290 2851.935 58.305 ;
        RECT 1070.025 57.990 2851.935 58.290 ;
        RECT 1070.025 57.975 1070.355 57.990 ;
        RECT 2851.605 57.975 2851.935 57.990 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.930 375.940 1077.250 376.000 ;
        RECT 1079.230 375.940 1079.550 376.000 ;
        RECT 1076.930 375.800 1079.550 375.940 ;
        RECT 1076.930 375.740 1077.250 375.800 ;
        RECT 1079.230 375.740 1079.550 375.800 ;
        RECT 1076.930 59.060 1077.250 59.120 ;
        RECT 2867.250 59.060 2867.570 59.120 ;
        RECT 1076.930 58.920 2867.570 59.060 ;
        RECT 1076.930 58.860 1077.250 58.920 ;
        RECT 2867.250 58.860 2867.570 58.920 ;
      LAYER via ;
        RECT 1076.960 375.740 1077.220 376.000 ;
        RECT 1079.260 375.740 1079.520 376.000 ;
        RECT 1076.960 58.860 1077.220 59.120 ;
        RECT 2867.280 58.860 2867.540 59.120 ;
      LAYER met2 ;
        RECT 1080.530 400.250 1080.810 404.000 ;
        RECT 1079.320 400.110 1080.810 400.250 ;
        RECT 1079.320 376.030 1079.460 400.110 ;
        RECT 1080.530 400.000 1080.810 400.110 ;
        RECT 1076.960 375.710 1077.220 376.030 ;
        RECT 1079.260 375.710 1079.520 376.030 ;
        RECT 1077.020 59.150 1077.160 375.710 ;
        RECT 1076.960 58.830 1077.220 59.150 ;
        RECT 2867.280 58.830 2867.540 59.150 ;
        RECT 2867.340 1.770 2867.480 58.830 ;
        RECT 2869.430 1.770 2869.990 2.400 ;
        RECT 2867.340 1.630 2869.990 1.770 ;
        RECT 2869.430 -4.800 2869.990 1.630 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.750 400.080 1085.070 400.140 ;
        RECT 1083.920 399.940 1085.070 400.080 ;
        RECT 1083.920 399.120 1084.060 399.940 ;
        RECT 1084.750 399.880 1085.070 399.940 ;
        RECT 1083.830 398.860 1084.150 399.120 ;
        RECT 1083.830 30.840 1084.150 30.900 ;
        RECT 2887.030 30.840 2887.350 30.900 ;
        RECT 1083.830 30.700 2887.350 30.840 ;
        RECT 1083.830 30.640 1084.150 30.700 ;
        RECT 2887.030 30.640 2887.350 30.700 ;
      LAYER via ;
        RECT 1084.780 399.880 1085.040 400.140 ;
        RECT 1083.860 398.860 1084.120 399.120 ;
        RECT 1083.860 30.640 1084.120 30.900 ;
        RECT 2887.060 30.640 2887.320 30.900 ;
      LAYER met2 ;
        RECT 1086.050 400.250 1086.330 404.000 ;
        RECT 1084.840 400.170 1086.330 400.250 ;
        RECT 1084.780 400.110 1086.330 400.170 ;
        RECT 1084.780 399.850 1085.040 400.110 ;
        RECT 1086.050 400.000 1086.330 400.110 ;
        RECT 1083.860 398.830 1084.120 399.150 ;
        RECT 1083.920 30.930 1084.060 398.830 ;
        RECT 1083.860 30.610 1084.120 30.930 ;
        RECT 2887.060 30.610 2887.320 30.930 ;
        RECT 2887.120 2.400 2887.260 30.610 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.470 378.320 455.790 378.380 ;
        RECT 458.690 378.320 459.010 378.380 ;
        RECT 455.470 378.180 459.010 378.320 ;
        RECT 455.470 378.120 455.790 378.180 ;
        RECT 458.690 378.120 459.010 378.180 ;
        RECT 455.470 28.800 455.790 28.860 ;
        RECT 607.270 28.800 607.590 28.860 ;
        RECT 455.470 28.660 607.590 28.800 ;
        RECT 455.470 28.600 455.790 28.660 ;
        RECT 607.270 28.600 607.590 28.660 ;
        RECT 607.270 18.940 607.590 19.000 ;
        RECT 847.850 18.940 848.170 19.000 ;
        RECT 607.270 18.800 848.170 18.940 ;
        RECT 607.270 18.740 607.590 18.800 ;
        RECT 847.850 18.740 848.170 18.800 ;
      LAYER via ;
        RECT 455.500 378.120 455.760 378.380 ;
        RECT 458.720 378.120 458.980 378.380 ;
        RECT 455.500 28.600 455.760 28.860 ;
        RECT 607.300 28.600 607.560 28.860 ;
        RECT 607.300 18.740 607.560 19.000 ;
        RECT 847.880 18.740 848.140 19.000 ;
      LAYER met2 ;
        RECT 459.990 400.250 460.270 404.000 ;
        RECT 458.780 400.110 460.270 400.250 ;
        RECT 458.780 378.410 458.920 400.110 ;
        RECT 459.990 400.000 460.270 400.110 ;
        RECT 455.500 378.090 455.760 378.410 ;
        RECT 458.720 378.090 458.980 378.410 ;
        RECT 455.560 28.890 455.700 378.090 ;
        RECT 455.500 28.570 455.760 28.890 ;
        RECT 607.300 28.570 607.560 28.890 ;
        RECT 607.360 19.030 607.500 28.570 ;
        RECT 607.300 18.710 607.560 19.030 ;
        RECT 847.880 18.710 848.140 19.030 ;
        RECT 847.940 2.400 848.080 18.710 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.830 40.360 463.150 40.420 ;
        RECT 656.030 40.360 656.350 40.420 ;
        RECT 462.830 40.220 656.350 40.360 ;
        RECT 462.830 40.160 463.150 40.220 ;
        RECT 656.030 40.160 656.350 40.220 ;
        RECT 656.030 20.300 656.350 20.360 ;
        RECT 865.790 20.300 866.110 20.360 ;
        RECT 656.030 20.160 866.110 20.300 ;
        RECT 656.030 20.100 656.350 20.160 ;
        RECT 865.790 20.100 866.110 20.160 ;
      LAYER via ;
        RECT 462.860 40.160 463.120 40.420 ;
        RECT 656.060 40.160 656.320 40.420 ;
        RECT 656.060 20.100 656.320 20.360 ;
        RECT 865.820 20.100 866.080 20.360 ;
      LAYER met2 ;
        RECT 465.510 400.250 465.790 404.000 ;
        RECT 464.300 400.110 465.790 400.250 ;
        RECT 464.300 399.570 464.440 400.110 ;
        RECT 465.510 400.000 465.790 400.110 ;
        RECT 462.920 399.430 464.440 399.570 ;
        RECT 462.920 40.450 463.060 399.430 ;
        RECT 462.860 40.130 463.120 40.450 ;
        RECT 656.060 40.130 656.320 40.450 ;
        RECT 656.120 20.390 656.260 40.130 ;
        RECT 656.060 20.070 656.320 20.390 ;
        RECT 865.820 20.070 866.080 20.390 ;
        RECT 865.880 2.400 866.020 20.070 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.270 52.600 469.590 52.660 ;
        RECT 884.650 52.600 884.970 52.660 ;
        RECT 469.270 52.460 884.970 52.600 ;
        RECT 469.270 52.400 469.590 52.460 ;
        RECT 884.650 52.400 884.970 52.460 ;
      LAYER via ;
        RECT 469.300 52.400 469.560 52.660 ;
        RECT 884.680 52.400 884.940 52.660 ;
      LAYER met2 ;
        RECT 470.570 400.250 470.850 404.000 ;
        RECT 469.360 400.110 470.850 400.250 ;
        RECT 469.360 52.690 469.500 400.110 ;
        RECT 470.570 400.000 470.850 400.110 ;
        RECT 469.300 52.370 469.560 52.690 ;
        RECT 884.680 52.370 884.940 52.690 ;
        RECT 884.740 9.930 884.880 52.370 ;
        RECT 883.360 9.790 884.880 9.930 ;
        RECT 883.360 2.400 883.500 9.790 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.170 393.280 476.490 393.340 ;
        RECT 637.630 393.280 637.950 393.340 ;
        RECT 476.170 393.140 637.950 393.280 ;
        RECT 476.170 393.080 476.490 393.140 ;
        RECT 637.630 393.080 637.950 393.140 ;
        RECT 638.090 22.680 638.410 22.740 ;
        RECT 901.210 22.680 901.530 22.740 ;
        RECT 638.090 22.540 901.530 22.680 ;
        RECT 638.090 22.480 638.410 22.540 ;
        RECT 901.210 22.480 901.530 22.540 ;
      LAYER via ;
        RECT 476.200 393.080 476.460 393.340 ;
        RECT 637.660 393.080 637.920 393.340 ;
        RECT 638.120 22.480 638.380 22.740 ;
        RECT 901.240 22.480 901.500 22.740 ;
      LAYER met2 ;
        RECT 476.090 400.180 476.370 404.000 ;
        RECT 476.090 400.000 476.400 400.180 ;
        RECT 476.260 393.370 476.400 400.000 ;
        RECT 476.200 393.050 476.460 393.370 ;
        RECT 637.660 393.050 637.920 393.370 ;
        RECT 637.720 351.970 637.860 393.050 ;
        RECT 637.720 351.830 638.320 351.970 ;
        RECT 638.180 22.770 638.320 351.830 ;
        RECT 638.120 22.450 638.380 22.770 ;
        RECT 901.240 22.450 901.500 22.770 ;
        RECT 901.300 2.400 901.440 22.450 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 481.690 392.600 482.010 392.660 ;
        RECT 658.790 392.600 659.110 392.660 ;
        RECT 481.690 392.460 659.110 392.600 ;
        RECT 481.690 392.400 482.010 392.460 ;
        RECT 658.790 392.400 659.110 392.460 ;
        RECT 658.790 22.340 659.110 22.400 ;
        RECT 918.690 22.340 919.010 22.400 ;
        RECT 658.790 22.200 919.010 22.340 ;
        RECT 658.790 22.140 659.110 22.200 ;
        RECT 918.690 22.140 919.010 22.200 ;
      LAYER via ;
        RECT 481.720 392.400 481.980 392.660 ;
        RECT 658.820 392.400 659.080 392.660 ;
        RECT 658.820 22.140 659.080 22.400 ;
        RECT 918.720 22.140 918.980 22.400 ;
      LAYER met2 ;
        RECT 481.610 400.180 481.890 404.000 ;
        RECT 481.610 400.000 481.920 400.180 ;
        RECT 481.780 392.690 481.920 400.000 ;
        RECT 481.720 392.370 481.980 392.690 ;
        RECT 658.820 392.370 659.080 392.690 ;
        RECT 658.880 22.430 659.020 392.370 ;
        RECT 658.820 22.110 659.080 22.430 ;
        RECT 918.720 22.110 918.980 22.430 ;
        RECT 918.780 2.400 918.920 22.110 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 541.490 392.940 541.810 393.000 ;
        RECT 617.390 392.940 617.710 393.000 ;
        RECT 541.490 392.800 617.710 392.940 ;
        RECT 541.490 392.740 541.810 392.800 ;
        RECT 617.390 392.740 617.710 392.800 ;
        RECT 487.210 390.560 487.530 390.620 ;
        RECT 541.490 390.560 541.810 390.620 ;
        RECT 487.210 390.420 541.810 390.560 ;
        RECT 487.210 390.360 487.530 390.420 ;
        RECT 541.490 390.360 541.810 390.420 ;
        RECT 617.390 389.540 617.710 389.600 ;
        RECT 666.150 389.540 666.470 389.600 ;
        RECT 617.390 389.400 666.470 389.540 ;
        RECT 617.390 389.340 617.710 389.400 ;
        RECT 666.150 389.340 666.470 389.400 ;
        RECT 665.690 23.020 666.010 23.080 ;
        RECT 936.630 23.020 936.950 23.080 ;
        RECT 665.690 22.880 936.950 23.020 ;
        RECT 665.690 22.820 666.010 22.880 ;
        RECT 936.630 22.820 936.950 22.880 ;
      LAYER via ;
        RECT 541.520 392.740 541.780 393.000 ;
        RECT 617.420 392.740 617.680 393.000 ;
        RECT 487.240 390.360 487.500 390.620 ;
        RECT 541.520 390.360 541.780 390.620 ;
        RECT 617.420 389.340 617.680 389.600 ;
        RECT 666.180 389.340 666.440 389.600 ;
        RECT 665.720 22.820 665.980 23.080 ;
        RECT 936.660 22.820 936.920 23.080 ;
      LAYER met2 ;
        RECT 487.130 400.180 487.410 404.000 ;
        RECT 487.130 400.000 487.440 400.180 ;
        RECT 487.300 390.650 487.440 400.000 ;
        RECT 541.520 392.710 541.780 393.030 ;
        RECT 617.420 392.710 617.680 393.030 ;
        RECT 541.580 390.650 541.720 392.710 ;
        RECT 487.240 390.330 487.500 390.650 ;
        RECT 541.520 390.330 541.780 390.650 ;
        RECT 617.480 389.630 617.620 392.710 ;
        RECT 617.420 389.310 617.680 389.630 ;
        RECT 666.180 389.310 666.440 389.630 ;
        RECT 666.240 324.370 666.380 389.310 ;
        RECT 665.780 324.230 666.380 324.370 ;
        RECT 665.780 23.110 665.920 324.230 ;
        RECT 665.720 22.790 665.980 23.110 ;
        RECT 936.660 22.790 936.920 23.110 ;
        RECT 936.720 2.400 936.860 22.790 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 492.270 392.260 492.590 392.320 ;
        RECT 693.290 392.260 693.610 392.320 ;
        RECT 492.270 392.120 693.610 392.260 ;
        RECT 492.270 392.060 492.590 392.120 ;
        RECT 693.290 392.060 693.610 392.120 ;
        RECT 693.290 23.360 693.610 23.420 ;
        RECT 954.110 23.360 954.430 23.420 ;
        RECT 693.290 23.220 954.430 23.360 ;
        RECT 693.290 23.160 693.610 23.220 ;
        RECT 954.110 23.160 954.430 23.220 ;
      LAYER via ;
        RECT 492.300 392.060 492.560 392.320 ;
        RECT 693.320 392.060 693.580 392.320 ;
        RECT 693.320 23.160 693.580 23.420 ;
        RECT 954.140 23.160 954.400 23.420 ;
      LAYER met2 ;
        RECT 492.650 400.250 492.930 404.000 ;
        RECT 492.360 400.110 492.930 400.250 ;
        RECT 492.360 392.350 492.500 400.110 ;
        RECT 492.650 400.000 492.930 400.110 ;
        RECT 492.300 392.030 492.560 392.350 ;
        RECT 693.320 392.030 693.580 392.350 ;
        RECT 693.380 23.450 693.520 392.030 ;
        RECT 693.320 23.130 693.580 23.450 ;
        RECT 954.140 23.130 954.400 23.450 ;
        RECT 954.200 2.400 954.340 23.130 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 498.250 391.580 498.570 391.640 ;
        RECT 713.990 391.580 714.310 391.640 ;
        RECT 498.250 391.440 714.310 391.580 ;
        RECT 498.250 391.380 498.570 391.440 ;
        RECT 713.990 391.380 714.310 391.440 ;
        RECT 713.990 23.700 714.310 23.760 ;
        RECT 972.050 23.700 972.370 23.760 ;
        RECT 713.990 23.560 972.370 23.700 ;
        RECT 713.990 23.500 714.310 23.560 ;
        RECT 972.050 23.500 972.370 23.560 ;
      LAYER via ;
        RECT 498.280 391.380 498.540 391.640 ;
        RECT 714.020 391.380 714.280 391.640 ;
        RECT 714.020 23.500 714.280 23.760 ;
        RECT 972.080 23.500 972.340 23.760 ;
      LAYER met2 ;
        RECT 498.170 400.180 498.450 404.000 ;
        RECT 498.170 400.000 498.480 400.180 ;
        RECT 498.340 391.670 498.480 400.000 ;
        RECT 498.280 391.350 498.540 391.670 ;
        RECT 714.020 391.350 714.280 391.670 ;
        RECT 714.080 23.790 714.220 391.350 ;
        RECT 714.020 23.470 714.280 23.790 ;
        RECT 972.080 23.470 972.340 23.790 ;
        RECT 972.140 2.400 972.280 23.470 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 400.730 39.340 401.050 39.400 ;
        RECT 652.810 39.340 653.130 39.400 ;
        RECT 400.730 39.200 653.130 39.340 ;
        RECT 400.730 39.140 401.050 39.200 ;
        RECT 652.810 39.140 653.130 39.200 ;
      LAYER via ;
        RECT 400.760 39.140 401.020 39.400 ;
        RECT 652.840 39.140 653.100 39.400 ;
      LAYER met2 ;
        RECT 400.190 400.250 400.470 404.000 ;
        RECT 400.190 400.110 400.960 400.250 ;
        RECT 400.190 400.000 400.470 400.110 ;
        RECT 400.820 39.430 400.960 400.110 ;
        RECT 400.760 39.110 401.020 39.430 ;
        RECT 652.840 39.110 653.100 39.430 ;
        RECT 652.900 2.400 653.040 39.110 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.330 386.140 497.650 386.200 ;
        RECT 501.930 386.140 502.250 386.200 ;
        RECT 497.330 386.000 502.250 386.140 ;
        RECT 497.330 385.940 497.650 386.000 ;
        RECT 501.930 385.940 502.250 386.000 ;
        RECT 497.330 49.880 497.650 49.940 ;
        RECT 989.530 49.880 989.850 49.940 ;
        RECT 497.330 49.740 989.850 49.880 ;
        RECT 497.330 49.680 497.650 49.740 ;
        RECT 989.530 49.680 989.850 49.740 ;
      LAYER via ;
        RECT 497.360 385.940 497.620 386.200 ;
        RECT 501.960 385.940 502.220 386.200 ;
        RECT 497.360 49.680 497.620 49.940 ;
        RECT 989.560 49.680 989.820 49.940 ;
      LAYER met2 ;
        RECT 503.230 400.250 503.510 404.000 ;
        RECT 502.020 400.110 503.510 400.250 ;
        RECT 502.020 386.230 502.160 400.110 ;
        RECT 503.230 400.000 503.510 400.110 ;
        RECT 497.360 385.910 497.620 386.230 ;
        RECT 501.960 385.910 502.220 386.230 ;
        RECT 497.420 49.970 497.560 385.910 ;
        RECT 497.360 49.650 497.620 49.970 ;
        RECT 989.560 49.650 989.820 49.970 ;
        RECT 989.620 2.400 989.760 49.650 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.230 386.140 504.550 386.200 ;
        RECT 507.450 386.140 507.770 386.200 ;
        RECT 504.230 386.000 507.770 386.140 ;
        RECT 504.230 385.940 504.550 386.000 ;
        RECT 507.450 385.940 507.770 386.000 ;
        RECT 504.230 59.740 504.550 59.800 ;
        RECT 1009.310 59.740 1009.630 59.800 ;
        RECT 504.230 59.600 1009.630 59.740 ;
        RECT 504.230 59.540 504.550 59.600 ;
        RECT 1009.310 59.540 1009.630 59.600 ;
        RECT 1007.470 20.980 1007.790 21.040 ;
        RECT 1009.310 20.980 1009.630 21.040 ;
        RECT 1007.470 20.840 1009.630 20.980 ;
        RECT 1007.470 20.780 1007.790 20.840 ;
        RECT 1009.310 20.780 1009.630 20.840 ;
      LAYER via ;
        RECT 504.260 385.940 504.520 386.200 ;
        RECT 507.480 385.940 507.740 386.200 ;
        RECT 504.260 59.540 504.520 59.800 ;
        RECT 1009.340 59.540 1009.600 59.800 ;
        RECT 1007.500 20.780 1007.760 21.040 ;
        RECT 1009.340 20.780 1009.600 21.040 ;
      LAYER met2 ;
        RECT 508.750 400.250 509.030 404.000 ;
        RECT 507.540 400.110 509.030 400.250 ;
        RECT 507.540 386.230 507.680 400.110 ;
        RECT 508.750 400.000 509.030 400.110 ;
        RECT 504.260 385.910 504.520 386.230 ;
        RECT 507.480 385.910 507.740 386.230 ;
        RECT 504.320 59.830 504.460 385.910 ;
        RECT 504.260 59.510 504.520 59.830 ;
        RECT 1009.340 59.510 1009.600 59.830 ;
        RECT 1009.400 21.070 1009.540 59.510 ;
        RECT 1007.500 20.750 1007.760 21.070 ;
        RECT 1009.340 20.750 1009.600 21.070 ;
        RECT 1007.560 2.400 1007.700 20.750 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 514.350 391.920 514.670 391.980 ;
        RECT 720.890 391.920 721.210 391.980 ;
        RECT 514.350 391.780 721.210 391.920 ;
        RECT 514.350 391.720 514.670 391.780 ;
        RECT 720.890 391.720 721.210 391.780 ;
        RECT 720.890 22.000 721.210 22.060 ;
        RECT 1025.410 22.000 1025.730 22.060 ;
        RECT 720.890 21.860 1025.730 22.000 ;
        RECT 720.890 21.800 721.210 21.860 ;
        RECT 1025.410 21.800 1025.730 21.860 ;
      LAYER via ;
        RECT 514.380 391.720 514.640 391.980 ;
        RECT 720.920 391.720 721.180 391.980 ;
        RECT 720.920 21.800 721.180 22.060 ;
        RECT 1025.440 21.800 1025.700 22.060 ;
      LAYER met2 ;
        RECT 514.270 400.180 514.550 404.000 ;
        RECT 514.270 400.000 514.580 400.180 ;
        RECT 514.440 392.010 514.580 400.000 ;
        RECT 514.380 391.690 514.640 392.010 ;
        RECT 720.920 391.690 721.180 392.010 ;
        RECT 720.980 22.090 721.120 391.690 ;
        RECT 720.920 21.770 721.180 22.090 ;
        RECT 1025.440 21.770 1025.700 22.090 ;
        RECT 1025.500 2.400 1025.640 21.770 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 568.630 390.900 568.950 390.960 ;
        RECT 749.410 390.900 749.730 390.960 ;
        RECT 568.630 390.760 749.730 390.900 ;
        RECT 568.630 390.700 568.950 390.760 ;
        RECT 749.410 390.700 749.730 390.760 ;
        RECT 519.870 388.180 520.190 388.240 ;
        RECT 568.630 388.180 568.950 388.240 ;
        RECT 519.870 388.040 568.950 388.180 ;
        RECT 519.870 387.980 520.190 388.040 ;
        RECT 568.630 387.980 568.950 388.040 ;
        RECT 748.490 21.660 748.810 21.720 ;
        RECT 1042.890 21.660 1043.210 21.720 ;
        RECT 748.490 21.520 1043.210 21.660 ;
        RECT 748.490 21.460 748.810 21.520 ;
        RECT 1042.890 21.460 1043.210 21.520 ;
      LAYER via ;
        RECT 568.660 390.700 568.920 390.960 ;
        RECT 749.440 390.700 749.700 390.960 ;
        RECT 519.900 387.980 520.160 388.240 ;
        RECT 568.660 387.980 568.920 388.240 ;
        RECT 748.520 21.460 748.780 21.720 ;
        RECT 1042.920 21.460 1043.180 21.720 ;
      LAYER met2 ;
        RECT 519.790 400.180 520.070 404.000 ;
        RECT 519.790 400.000 520.100 400.180 ;
        RECT 519.960 388.270 520.100 400.000 ;
        RECT 568.660 390.670 568.920 390.990 ;
        RECT 749.440 390.670 749.700 390.990 ;
        RECT 568.720 388.270 568.860 390.670 ;
        RECT 519.900 387.950 520.160 388.270 ;
        RECT 568.660 387.950 568.920 388.270 ;
        RECT 749.500 324.370 749.640 390.670 ;
        RECT 748.580 324.230 749.640 324.370 ;
        RECT 748.580 21.750 748.720 324.230 ;
        RECT 748.520 21.430 748.780 21.750 ;
        RECT 1042.920 21.430 1043.180 21.750 ;
        RECT 1042.980 2.400 1043.120 21.430 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 525.390 387.840 525.710 387.900 ;
        RECT 610.490 387.840 610.810 387.900 ;
        RECT 525.390 387.700 610.810 387.840 ;
        RECT 525.390 387.640 525.710 387.700 ;
        RECT 610.490 387.640 610.810 387.700 ;
        RECT 610.950 30.840 611.270 30.900 ;
        RECT 1060.830 30.840 1061.150 30.900 ;
        RECT 610.950 30.700 1061.150 30.840 ;
        RECT 610.950 30.640 611.270 30.700 ;
        RECT 1060.830 30.640 1061.150 30.700 ;
      LAYER via ;
        RECT 525.420 387.640 525.680 387.900 ;
        RECT 610.520 387.640 610.780 387.900 ;
        RECT 610.980 30.640 611.240 30.900 ;
        RECT 1060.860 30.640 1061.120 30.900 ;
      LAYER met2 ;
        RECT 525.310 400.180 525.590 404.000 ;
        RECT 525.310 400.000 525.620 400.180 ;
        RECT 525.480 387.930 525.620 400.000 ;
        RECT 525.420 387.610 525.680 387.930 ;
        RECT 610.520 387.610 610.780 387.930 ;
        RECT 610.580 375.770 610.720 387.610 ;
        RECT 610.580 375.630 611.180 375.770 ;
        RECT 611.040 30.930 611.180 375.630 ;
        RECT 610.980 30.610 611.240 30.930 ;
        RECT 1060.860 30.610 1061.120 30.930 ;
        RECT 1060.920 2.400 1061.060 30.610 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.930 385.800 525.250 385.860 ;
        RECT 529.530 385.800 529.850 385.860 ;
        RECT 524.930 385.660 529.850 385.800 ;
        RECT 524.930 385.600 525.250 385.660 ;
        RECT 529.530 385.600 529.850 385.660 ;
        RECT 524.930 56.680 525.250 56.740 ;
        RECT 1076.930 56.680 1077.250 56.740 ;
        RECT 524.930 56.540 1077.250 56.680 ;
        RECT 524.930 56.480 525.250 56.540 ;
        RECT 1076.930 56.480 1077.250 56.540 ;
      LAYER via ;
        RECT 524.960 385.600 525.220 385.860 ;
        RECT 529.560 385.600 529.820 385.860 ;
        RECT 524.960 56.480 525.220 56.740 ;
        RECT 1076.960 56.480 1077.220 56.740 ;
      LAYER met2 ;
        RECT 530.830 400.250 531.110 404.000 ;
        RECT 529.620 400.110 531.110 400.250 ;
        RECT 529.620 385.890 529.760 400.110 ;
        RECT 530.830 400.000 531.110 400.110 ;
        RECT 524.960 385.570 525.220 385.890 ;
        RECT 529.560 385.570 529.820 385.890 ;
        RECT 525.020 56.770 525.160 385.570 ;
        RECT 524.960 56.450 525.220 56.770 ;
        RECT 1076.960 56.450 1077.220 56.770 ;
        RECT 1077.020 1.770 1077.160 56.450 ;
        RECT 1078.190 1.770 1078.750 2.400 ;
        RECT 1077.020 1.630 1078.750 1.770 ;
        RECT 1078.190 -4.800 1078.750 1.630 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.370 387.160 531.690 387.220 ;
        RECT 534.590 387.160 534.910 387.220 ;
        RECT 531.370 387.020 534.910 387.160 ;
        RECT 531.370 386.960 531.690 387.020 ;
        RECT 534.590 386.960 534.910 387.020 ;
        RECT 531.370 57.020 531.690 57.080 ;
        RECT 1090.270 57.020 1090.590 57.080 ;
        RECT 531.370 56.880 1090.590 57.020 ;
        RECT 531.370 56.820 531.690 56.880 ;
        RECT 1090.270 56.820 1090.590 56.880 ;
        RECT 1090.270 17.240 1090.590 17.300 ;
        RECT 1096.250 17.240 1096.570 17.300 ;
        RECT 1090.270 17.100 1096.570 17.240 ;
        RECT 1090.270 17.040 1090.590 17.100 ;
        RECT 1096.250 17.040 1096.570 17.100 ;
      LAYER via ;
        RECT 531.400 386.960 531.660 387.220 ;
        RECT 534.620 386.960 534.880 387.220 ;
        RECT 531.400 56.820 531.660 57.080 ;
        RECT 1090.300 56.820 1090.560 57.080 ;
        RECT 1090.300 17.040 1090.560 17.300 ;
        RECT 1096.280 17.040 1096.540 17.300 ;
      LAYER met2 ;
        RECT 535.890 400.250 536.170 404.000 ;
        RECT 534.680 400.110 536.170 400.250 ;
        RECT 534.680 387.250 534.820 400.110 ;
        RECT 535.890 400.000 536.170 400.110 ;
        RECT 531.400 386.930 531.660 387.250 ;
        RECT 534.620 386.930 534.880 387.250 ;
        RECT 531.460 57.110 531.600 386.930 ;
        RECT 531.400 56.790 531.660 57.110 ;
        RECT 1090.300 56.790 1090.560 57.110 ;
        RECT 1090.360 17.330 1090.500 56.790 ;
        RECT 1090.300 17.010 1090.560 17.330 ;
        RECT 1096.280 17.010 1096.540 17.330 ;
        RECT 1096.340 2.400 1096.480 17.010 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.730 105.300 539.050 105.360 ;
        RECT 1110.970 105.300 1111.290 105.360 ;
        RECT 538.730 105.160 1111.290 105.300 ;
        RECT 538.730 105.100 539.050 105.160 ;
        RECT 1110.970 105.100 1111.290 105.160 ;
      LAYER via ;
        RECT 538.760 105.100 539.020 105.360 ;
        RECT 1111.000 105.100 1111.260 105.360 ;
      LAYER met2 ;
        RECT 541.410 400.250 541.690 404.000 ;
        RECT 540.200 400.110 541.690 400.250 ;
        RECT 540.200 324.370 540.340 400.110 ;
        RECT 541.410 400.000 541.690 400.110 ;
        RECT 538.820 324.230 540.340 324.370 ;
        RECT 538.820 105.390 538.960 324.230 ;
        RECT 538.760 105.070 539.020 105.390 ;
        RECT 1111.000 105.070 1111.260 105.390 ;
        RECT 1111.060 82.870 1111.200 105.070 ;
        RECT 1111.060 82.730 1113.960 82.870 ;
        RECT 1113.820 2.400 1113.960 82.730 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.550 112.100 546.870 112.160 ;
        RECT 1131.670 112.100 1131.990 112.160 ;
        RECT 546.550 111.960 1131.990 112.100 ;
        RECT 546.550 111.900 546.870 111.960 ;
        RECT 1131.670 111.900 1131.990 111.960 ;
      LAYER via ;
        RECT 546.580 111.900 546.840 112.160 ;
        RECT 1131.700 111.900 1131.960 112.160 ;
      LAYER met2 ;
        RECT 546.930 400.250 547.210 404.000 ;
        RECT 546.640 400.110 547.210 400.250 ;
        RECT 546.640 112.190 546.780 400.110 ;
        RECT 546.930 400.000 547.210 400.110 ;
        RECT 546.580 111.870 546.840 112.190 ;
        RECT 1131.700 111.870 1131.960 112.190 ;
        RECT 1131.760 2.400 1131.900 111.870 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.990 112.440 553.310 112.500 ;
        RECT 1145.470 112.440 1145.790 112.500 ;
        RECT 552.990 112.300 1145.790 112.440 ;
        RECT 552.990 112.240 553.310 112.300 ;
        RECT 1145.470 112.240 1145.790 112.300 ;
      LAYER via ;
        RECT 553.020 112.240 553.280 112.500 ;
        RECT 1145.500 112.240 1145.760 112.500 ;
      LAYER met2 ;
        RECT 552.450 400.250 552.730 404.000 ;
        RECT 552.450 400.110 553.220 400.250 ;
        RECT 552.450 400.000 552.730 400.110 ;
        RECT 553.080 112.530 553.220 400.110 ;
        RECT 553.020 112.210 553.280 112.530 ;
        RECT 1145.500 112.210 1145.760 112.530 ;
        RECT 1145.560 82.870 1145.700 112.210 ;
        RECT 1145.560 82.730 1147.080 82.870 ;
        RECT 1146.940 1.770 1147.080 82.730 ;
        RECT 1149.030 1.770 1149.590 2.400 ;
        RECT 1146.940 1.630 1149.590 1.770 ;
        RECT 1149.030 -4.800 1149.590 1.630 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 401.190 39.000 401.510 39.060 ;
        RECT 670.750 39.000 671.070 39.060 ;
        RECT 401.190 38.860 671.070 39.000 ;
        RECT 401.190 38.800 401.510 38.860 ;
        RECT 670.750 38.800 671.070 38.860 ;
      LAYER via ;
        RECT 401.220 38.800 401.480 39.060 ;
        RECT 670.780 38.800 671.040 39.060 ;
      LAYER met2 ;
        RECT 405.250 400.250 405.530 404.000 ;
        RECT 404.040 400.110 405.530 400.250 ;
        RECT 404.040 386.470 404.180 400.110 ;
        RECT 405.250 400.000 405.530 400.110 ;
        RECT 401.280 386.330 404.180 386.470 ;
        RECT 401.280 39.090 401.420 386.330 ;
        RECT 401.220 38.770 401.480 39.090 ;
        RECT 670.780 38.770 671.040 39.090 ;
        RECT 670.840 2.400 670.980 38.770 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 553.450 112.780 553.770 112.840 ;
        RECT 1166.170 112.780 1166.490 112.840 ;
        RECT 553.450 112.640 1166.490 112.780 ;
        RECT 553.450 112.580 553.770 112.640 ;
        RECT 1166.170 112.580 1166.490 112.640 ;
      LAYER via ;
        RECT 553.480 112.580 553.740 112.840 ;
        RECT 1166.200 112.580 1166.460 112.840 ;
      LAYER met2 ;
        RECT 557.970 400.250 558.250 404.000 ;
        RECT 556.760 400.110 558.250 400.250 ;
        RECT 556.760 324.370 556.900 400.110 ;
        RECT 557.970 400.000 558.250 400.110 ;
        RECT 553.540 324.230 556.900 324.370 ;
        RECT 553.540 112.870 553.680 324.230 ;
        RECT 553.480 112.550 553.740 112.870 ;
        RECT 1166.200 112.550 1166.460 112.870 ;
        RECT 1166.260 82.870 1166.400 112.550 ;
        RECT 1166.260 82.730 1167.320 82.870 ;
        RECT 1167.180 2.400 1167.320 82.730 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.430 376.280 559.750 376.340 ;
        RECT 562.190 376.280 562.510 376.340 ;
        RECT 559.430 376.140 562.510 376.280 ;
        RECT 559.430 376.080 559.750 376.140 ;
        RECT 562.190 376.080 562.510 376.140 ;
        RECT 559.430 63.820 559.750 63.880 ;
        RECT 1182.730 63.820 1183.050 63.880 ;
        RECT 559.430 63.680 1183.050 63.820 ;
        RECT 559.430 63.620 559.750 63.680 ;
        RECT 1182.730 63.620 1183.050 63.680 ;
      LAYER via ;
        RECT 559.460 376.080 559.720 376.340 ;
        RECT 562.220 376.080 562.480 376.340 ;
        RECT 559.460 63.620 559.720 63.880 ;
        RECT 1182.760 63.620 1183.020 63.880 ;
      LAYER met2 ;
        RECT 563.490 400.250 563.770 404.000 ;
        RECT 562.280 400.110 563.770 400.250 ;
        RECT 562.280 376.370 562.420 400.110 ;
        RECT 563.490 400.000 563.770 400.110 ;
        RECT 559.460 376.050 559.720 376.370 ;
        RECT 562.220 376.050 562.480 376.370 ;
        RECT 559.520 63.910 559.660 376.050 ;
        RECT 559.460 63.590 559.720 63.910 ;
        RECT 1182.760 63.590 1183.020 63.910 ;
        RECT 1182.820 1.770 1182.960 63.590 ;
        RECT 1184.910 1.770 1185.470 2.400 ;
        RECT 1182.820 1.630 1185.470 1.770 ;
        RECT 1184.910 -4.800 1185.470 1.630 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.790 64.160 567.110 64.220 ;
        RECT 1200.670 64.160 1200.990 64.220 ;
        RECT 566.790 64.020 1200.990 64.160 ;
        RECT 566.790 63.960 567.110 64.020 ;
        RECT 1200.670 63.960 1200.990 64.020 ;
      LAYER via ;
        RECT 566.820 63.960 567.080 64.220 ;
        RECT 1200.700 63.960 1200.960 64.220 ;
      LAYER met2 ;
        RECT 568.550 400.250 568.830 404.000 ;
        RECT 567.800 400.110 568.830 400.250 ;
        RECT 567.800 351.970 567.940 400.110 ;
        RECT 568.550 400.000 568.830 400.110 ;
        RECT 566.880 351.830 567.940 351.970 ;
        RECT 566.880 64.250 567.020 351.830 ;
        RECT 566.820 63.930 567.080 64.250 ;
        RECT 1200.700 63.930 1200.960 64.250 ;
        RECT 1200.760 1.770 1200.900 63.930 ;
        RECT 1202.390 1.770 1202.950 2.400 ;
        RECT 1200.760 1.630 1202.950 1.770 ;
        RECT 1202.390 -4.800 1202.950 1.630 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.230 64.500 573.550 64.560 ;
        RECT 1214.470 64.500 1214.790 64.560 ;
        RECT 573.230 64.360 1214.790 64.500 ;
        RECT 573.230 64.300 573.550 64.360 ;
        RECT 1214.470 64.300 1214.790 64.360 ;
        RECT 1214.470 15.200 1214.790 15.260 ;
        RECT 1220.450 15.200 1220.770 15.260 ;
        RECT 1214.470 15.060 1220.770 15.200 ;
        RECT 1214.470 15.000 1214.790 15.060 ;
        RECT 1220.450 15.000 1220.770 15.060 ;
      LAYER via ;
        RECT 573.260 64.300 573.520 64.560 ;
        RECT 1214.500 64.300 1214.760 64.560 ;
        RECT 1214.500 15.000 1214.760 15.260 ;
        RECT 1220.480 15.000 1220.740 15.260 ;
      LAYER met2 ;
        RECT 574.070 400.250 574.350 404.000 ;
        RECT 573.320 400.110 574.350 400.250 ;
        RECT 573.320 64.590 573.460 400.110 ;
        RECT 574.070 400.000 574.350 400.110 ;
        RECT 573.260 64.270 573.520 64.590 ;
        RECT 1214.500 64.270 1214.760 64.590 ;
        RECT 1214.560 15.290 1214.700 64.270 ;
        RECT 1214.500 14.970 1214.760 15.290 ;
        RECT 1220.480 14.970 1220.740 15.290 ;
        RECT 1220.540 2.400 1220.680 14.970 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.590 64.840 580.910 64.900 ;
        RECT 1237.930 64.840 1238.250 64.900 ;
        RECT 580.590 64.700 1238.250 64.840 ;
        RECT 580.590 64.640 580.910 64.700 ;
        RECT 1237.930 64.640 1238.250 64.700 ;
      LAYER via ;
        RECT 580.620 64.640 580.880 64.900 ;
        RECT 1237.960 64.640 1238.220 64.900 ;
      LAYER met2 ;
        RECT 579.590 400.250 579.870 404.000 ;
        RECT 579.590 400.110 580.820 400.250 ;
        RECT 579.590 400.000 579.870 400.110 ;
        RECT 580.680 64.930 580.820 400.110 ;
        RECT 580.620 64.610 580.880 64.930 ;
        RECT 1237.960 64.610 1238.220 64.930 ;
        RECT 1238.020 2.400 1238.160 64.610 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 580.130 376.280 580.450 376.340 ;
        RECT 583.810 376.280 584.130 376.340 ;
        RECT 580.130 376.140 584.130 376.280 ;
        RECT 580.130 376.080 580.450 376.140 ;
        RECT 583.810 376.080 584.130 376.140 ;
        RECT 580.130 65.180 580.450 65.240 ;
        RECT 1256.330 65.180 1256.650 65.240 ;
        RECT 580.130 65.040 1256.650 65.180 ;
        RECT 580.130 64.980 580.450 65.040 ;
        RECT 1256.330 64.980 1256.650 65.040 ;
      LAYER via ;
        RECT 580.160 376.080 580.420 376.340 ;
        RECT 583.840 376.080 584.100 376.340 ;
        RECT 580.160 64.980 580.420 65.240 ;
        RECT 1256.360 64.980 1256.620 65.240 ;
      LAYER met2 ;
        RECT 585.110 400.250 585.390 404.000 ;
        RECT 583.900 400.110 585.390 400.250 ;
        RECT 583.900 376.370 584.040 400.110 ;
        RECT 585.110 400.000 585.390 400.110 ;
        RECT 580.160 376.050 580.420 376.370 ;
        RECT 583.840 376.050 584.100 376.370 ;
        RECT 580.220 65.270 580.360 376.050 ;
        RECT 580.160 64.950 580.420 65.270 ;
        RECT 1256.360 64.950 1256.620 65.270 ;
        RECT 1256.420 17.410 1256.560 64.950 ;
        RECT 1255.960 17.270 1256.560 17.410 ;
        RECT 1255.960 2.400 1256.100 17.270 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.030 375.940 587.350 376.000 ;
        RECT 589.330 375.940 589.650 376.000 ;
        RECT 587.030 375.800 589.650 375.940 ;
        RECT 587.030 375.740 587.350 375.800 ;
        RECT 589.330 375.740 589.650 375.800 ;
        RECT 587.030 68.920 587.350 68.980 ;
        RECT 1271.050 68.920 1271.370 68.980 ;
        RECT 587.030 68.780 1271.370 68.920 ;
        RECT 587.030 68.720 587.350 68.780 ;
        RECT 1271.050 68.720 1271.370 68.780 ;
      LAYER via ;
        RECT 587.060 375.740 587.320 376.000 ;
        RECT 589.360 375.740 589.620 376.000 ;
        RECT 587.060 68.720 587.320 68.980 ;
        RECT 1271.080 68.720 1271.340 68.980 ;
      LAYER met2 ;
        RECT 590.630 400.250 590.910 404.000 ;
        RECT 589.420 400.110 590.910 400.250 ;
        RECT 589.420 376.030 589.560 400.110 ;
        RECT 590.630 400.000 590.910 400.110 ;
        RECT 587.060 375.710 587.320 376.030 ;
        RECT 589.360 375.710 589.620 376.030 ;
        RECT 587.120 69.010 587.260 375.710 ;
        RECT 587.060 68.690 587.320 69.010 ;
        RECT 1271.080 68.690 1271.340 69.010 ;
        RECT 1271.140 1.770 1271.280 68.690 ;
        RECT 1273.230 1.770 1273.790 2.400 ;
        RECT 1271.140 1.630 1273.790 1.770 ;
        RECT 1273.230 -4.800 1273.790 1.630 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.390 68.580 594.710 68.640 ;
        RECT 1291.290 68.580 1291.610 68.640 ;
        RECT 594.390 68.440 1291.610 68.580 ;
        RECT 594.390 68.380 594.710 68.440 ;
        RECT 1291.290 68.380 1291.610 68.440 ;
      LAYER via ;
        RECT 594.420 68.380 594.680 68.640 ;
        RECT 1291.320 68.380 1291.580 68.640 ;
      LAYER met2 ;
        RECT 596.150 400.250 596.430 404.000 ;
        RECT 594.940 400.110 596.430 400.250 ;
        RECT 594.940 351.970 595.080 400.110 ;
        RECT 596.150 400.000 596.430 400.110 ;
        RECT 594.480 351.830 595.080 351.970 ;
        RECT 594.480 68.670 594.620 351.830 ;
        RECT 594.420 68.350 594.680 68.670 ;
        RECT 1291.320 68.350 1291.580 68.670 ;
        RECT 1291.380 2.400 1291.520 68.350 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.830 68.240 601.150 68.300 ;
        RECT 1308.770 68.240 1309.090 68.300 ;
        RECT 600.830 68.100 1309.090 68.240 ;
        RECT 600.830 68.040 601.150 68.100 ;
        RECT 1308.770 68.040 1309.090 68.100 ;
      LAYER via ;
        RECT 600.860 68.040 601.120 68.300 ;
        RECT 1308.800 68.040 1309.060 68.300 ;
      LAYER met2 ;
        RECT 601.210 400.250 601.490 404.000 ;
        RECT 600.920 400.110 601.490 400.250 ;
        RECT 600.920 68.330 601.060 400.110 ;
        RECT 601.210 400.000 601.490 400.110 ;
        RECT 600.860 68.010 601.120 68.330 ;
        RECT 1308.800 68.010 1309.060 68.330 ;
        RECT 1308.860 2.400 1309.000 68.010 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.290 376.280 601.610 376.340 ;
        RECT 605.430 376.280 605.750 376.340 ;
        RECT 601.290 376.140 605.750 376.280 ;
        RECT 601.290 376.080 601.610 376.140 ;
        RECT 605.430 376.080 605.750 376.140 ;
        RECT 601.290 67.900 601.610 67.960 ;
        RECT 1324.870 67.900 1325.190 67.960 ;
        RECT 601.290 67.760 1325.190 67.900 ;
        RECT 601.290 67.700 601.610 67.760 ;
        RECT 1324.870 67.700 1325.190 67.760 ;
      LAYER via ;
        RECT 601.320 376.080 601.580 376.340 ;
        RECT 605.460 376.080 605.720 376.340 ;
        RECT 601.320 67.700 601.580 67.960 ;
        RECT 1324.900 67.700 1325.160 67.960 ;
      LAYER met2 ;
        RECT 606.730 400.250 607.010 404.000 ;
        RECT 605.520 400.110 607.010 400.250 ;
        RECT 605.520 376.370 605.660 400.110 ;
        RECT 606.730 400.000 607.010 400.110 ;
        RECT 601.320 376.050 601.580 376.370 ;
        RECT 605.460 376.050 605.720 376.370 ;
        RECT 601.380 67.990 601.520 376.050 ;
        RECT 601.320 67.670 601.580 67.990 ;
        RECT 1324.900 67.670 1325.160 67.990 ;
        RECT 1324.960 1.770 1325.100 67.670 ;
        RECT 1326.590 1.770 1327.150 2.400 ;
        RECT 1324.960 1.630 1327.150 1.770 ;
        RECT 1326.590 -4.800 1327.150 1.630 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.550 38.320 408.870 38.380 ;
        RECT 688.230 38.320 688.550 38.380 ;
        RECT 408.550 38.180 688.550 38.320 ;
        RECT 408.550 38.120 408.870 38.180 ;
        RECT 688.230 38.120 688.550 38.180 ;
      LAYER via ;
        RECT 408.580 38.120 408.840 38.380 ;
        RECT 688.260 38.120 688.520 38.380 ;
      LAYER met2 ;
        RECT 410.770 400.250 411.050 404.000 ;
        RECT 409.560 400.110 411.050 400.250 ;
        RECT 409.560 324.370 409.700 400.110 ;
        RECT 410.770 400.000 411.050 400.110 ;
        RECT 408.640 324.230 409.700 324.370 ;
        RECT 408.640 38.410 408.780 324.230 ;
        RECT 408.580 38.090 408.840 38.410 ;
        RECT 688.260 38.090 688.520 38.410 ;
        RECT 688.320 2.400 688.460 38.090 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.270 376.280 607.590 376.340 ;
        RECT 610.950 376.280 611.270 376.340 ;
        RECT 607.270 376.140 611.270 376.280 ;
        RECT 607.270 376.080 607.590 376.140 ;
        RECT 610.950 376.080 611.270 376.140 ;
        RECT 607.270 67.560 607.590 67.620 ;
        RECT 1341.890 67.560 1342.210 67.620 ;
        RECT 607.270 67.420 1342.210 67.560 ;
        RECT 607.270 67.360 607.590 67.420 ;
        RECT 1341.890 67.360 1342.210 67.420 ;
      LAYER via ;
        RECT 607.300 376.080 607.560 376.340 ;
        RECT 610.980 376.080 611.240 376.340 ;
        RECT 607.300 67.360 607.560 67.620 ;
        RECT 1341.920 67.360 1342.180 67.620 ;
      LAYER met2 ;
        RECT 612.250 400.250 612.530 404.000 ;
        RECT 611.040 400.110 612.530 400.250 ;
        RECT 611.040 376.370 611.180 400.110 ;
        RECT 612.250 400.000 612.530 400.110 ;
        RECT 607.300 376.050 607.560 376.370 ;
        RECT 610.980 376.050 611.240 376.370 ;
        RECT 607.360 67.650 607.500 376.050 ;
        RECT 607.300 67.330 607.560 67.650 ;
        RECT 1341.920 67.330 1342.180 67.650 ;
        RECT 1341.980 1.770 1342.120 67.330 ;
        RECT 1344.070 1.770 1344.630 2.400 ;
        RECT 1341.980 1.630 1344.630 1.770 ;
        RECT 1344.070 -4.800 1344.630 1.630 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.170 375.940 614.490 376.000 ;
        RECT 616.470 375.940 616.790 376.000 ;
        RECT 614.170 375.800 616.790 375.940 ;
        RECT 614.170 375.740 614.490 375.800 ;
        RECT 616.470 375.740 616.790 375.800 ;
        RECT 614.170 67.220 614.490 67.280 ;
        RECT 1362.130 67.220 1362.450 67.280 ;
        RECT 614.170 67.080 1362.450 67.220 ;
        RECT 614.170 67.020 614.490 67.080 ;
        RECT 1362.130 67.020 1362.450 67.080 ;
      LAYER via ;
        RECT 614.200 375.740 614.460 376.000 ;
        RECT 616.500 375.740 616.760 376.000 ;
        RECT 614.200 67.020 614.460 67.280 ;
        RECT 1362.160 67.020 1362.420 67.280 ;
      LAYER met2 ;
        RECT 617.770 400.250 618.050 404.000 ;
        RECT 616.560 400.110 618.050 400.250 ;
        RECT 616.560 376.030 616.700 400.110 ;
        RECT 617.770 400.000 618.050 400.110 ;
        RECT 614.200 375.710 614.460 376.030 ;
        RECT 616.500 375.710 616.760 376.030 ;
        RECT 614.260 67.310 614.400 375.710 ;
        RECT 614.200 66.990 614.460 67.310 ;
        RECT 1362.160 66.990 1362.420 67.310 ;
        RECT 1362.220 2.400 1362.360 66.990 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.070 376.280 621.390 376.340 ;
        RECT 622.450 376.280 622.770 376.340 ;
        RECT 621.070 376.140 622.770 376.280 ;
        RECT 621.070 376.080 621.390 376.140 ;
        RECT 622.450 376.080 622.770 376.140 ;
        RECT 621.070 66.880 621.390 66.940 ;
        RECT 1380.530 66.880 1380.850 66.940 ;
        RECT 621.070 66.740 1380.850 66.880 ;
        RECT 621.070 66.680 621.390 66.740 ;
        RECT 1380.530 66.680 1380.850 66.740 ;
      LAYER via ;
        RECT 621.100 376.080 621.360 376.340 ;
        RECT 622.480 376.080 622.740 376.340 ;
        RECT 621.100 66.680 621.360 66.940 ;
        RECT 1380.560 66.680 1380.820 66.940 ;
      LAYER met2 ;
        RECT 623.290 400.250 623.570 404.000 ;
        RECT 622.540 400.110 623.570 400.250 ;
        RECT 622.540 376.370 622.680 400.110 ;
        RECT 623.290 400.000 623.570 400.110 ;
        RECT 621.100 376.050 621.360 376.370 ;
        RECT 622.480 376.050 622.740 376.370 ;
        RECT 621.160 66.970 621.300 376.050 ;
        RECT 621.100 66.650 621.360 66.970 ;
        RECT 1380.560 66.650 1380.820 66.970 ;
        RECT 1380.620 17.410 1380.760 66.650 ;
        RECT 1380.160 17.270 1380.760 17.410 ;
        RECT 1380.160 2.400 1380.300 17.270 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 627.970 66.540 628.290 66.600 ;
        RECT 1395.250 66.540 1395.570 66.600 ;
        RECT 627.970 66.400 1395.570 66.540 ;
        RECT 627.970 66.340 628.290 66.400 ;
        RECT 1395.250 66.340 1395.570 66.400 ;
      LAYER via ;
        RECT 628.000 66.340 628.260 66.600 ;
        RECT 1395.280 66.340 1395.540 66.600 ;
      LAYER met2 ;
        RECT 628.810 400.250 629.090 404.000 ;
        RECT 628.060 400.110 629.090 400.250 ;
        RECT 628.060 66.630 628.200 400.110 ;
        RECT 628.810 400.000 629.090 400.110 ;
        RECT 628.000 66.310 628.260 66.630 ;
        RECT 1395.280 66.310 1395.540 66.630 ;
        RECT 1395.340 1.770 1395.480 66.310 ;
        RECT 1397.430 1.770 1397.990 2.400 ;
        RECT 1395.340 1.630 1397.990 1.770 ;
        RECT 1397.430 -4.800 1397.990 1.630 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.430 376.280 628.750 376.340 ;
        RECT 633.030 376.280 633.350 376.340 ;
        RECT 628.430 376.140 633.350 376.280 ;
        RECT 628.430 376.080 628.750 376.140 ;
        RECT 633.030 376.080 633.350 376.140 ;
        RECT 628.430 66.200 628.750 66.260 ;
        RECT 1415.490 66.200 1415.810 66.260 ;
        RECT 628.430 66.060 1415.810 66.200 ;
        RECT 628.430 66.000 628.750 66.060 ;
        RECT 1415.490 66.000 1415.810 66.060 ;
      LAYER via ;
        RECT 628.460 376.080 628.720 376.340 ;
        RECT 633.060 376.080 633.320 376.340 ;
        RECT 628.460 66.000 628.720 66.260 ;
        RECT 1415.520 66.000 1415.780 66.260 ;
      LAYER met2 ;
        RECT 633.870 400.250 634.150 404.000 ;
        RECT 633.120 400.110 634.150 400.250 ;
        RECT 633.120 376.370 633.260 400.110 ;
        RECT 633.870 400.000 634.150 400.110 ;
        RECT 628.460 376.050 628.720 376.370 ;
        RECT 633.060 376.050 633.320 376.370 ;
        RECT 628.520 66.290 628.660 376.050 ;
        RECT 628.460 65.970 628.720 66.290 ;
        RECT 1415.520 65.970 1415.780 66.290 ;
        RECT 1415.580 2.400 1415.720 65.970 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.330 376.280 635.650 376.340 ;
        RECT 638.090 376.280 638.410 376.340 ;
        RECT 635.330 376.140 638.410 376.280 ;
        RECT 635.330 376.080 635.650 376.140 ;
        RECT 638.090 376.080 638.410 376.140 ;
        RECT 635.330 65.860 635.650 65.920 ;
        RECT 1432.970 65.860 1433.290 65.920 ;
        RECT 635.330 65.720 1433.290 65.860 ;
        RECT 635.330 65.660 635.650 65.720 ;
        RECT 1432.970 65.660 1433.290 65.720 ;
      LAYER via ;
        RECT 635.360 376.080 635.620 376.340 ;
        RECT 638.120 376.080 638.380 376.340 ;
        RECT 635.360 65.660 635.620 65.920 ;
        RECT 1433.000 65.660 1433.260 65.920 ;
      LAYER met2 ;
        RECT 639.390 400.250 639.670 404.000 ;
        RECT 638.180 400.110 639.670 400.250 ;
        RECT 638.180 376.370 638.320 400.110 ;
        RECT 639.390 400.000 639.670 400.110 ;
        RECT 635.360 376.050 635.620 376.370 ;
        RECT 638.120 376.050 638.380 376.370 ;
        RECT 635.420 65.950 635.560 376.050 ;
        RECT 635.360 65.630 635.620 65.950 ;
        RECT 1433.000 65.630 1433.260 65.950 ;
        RECT 1433.060 2.400 1433.200 65.630 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.230 65.520 642.550 65.580 ;
        RECT 1449.070 65.520 1449.390 65.580 ;
        RECT 642.230 65.380 1449.390 65.520 ;
        RECT 642.230 65.320 642.550 65.380 ;
        RECT 1449.070 65.320 1449.390 65.380 ;
      LAYER via ;
        RECT 642.260 65.320 642.520 65.580 ;
        RECT 1449.100 65.320 1449.360 65.580 ;
      LAYER met2 ;
        RECT 644.910 400.250 645.190 404.000 ;
        RECT 643.700 400.110 645.190 400.250 ;
        RECT 643.700 386.480 643.840 400.110 ;
        RECT 644.910 400.000 645.190 400.110 ;
        RECT 642.320 386.340 643.840 386.480 ;
        RECT 642.320 65.610 642.460 386.340 ;
        RECT 642.260 65.290 642.520 65.610 ;
        RECT 1449.100 65.290 1449.360 65.610 ;
        RECT 1449.160 1.770 1449.300 65.290 ;
        RECT 1450.790 1.770 1451.350 2.400 ;
        RECT 1449.160 1.630 1451.350 1.770 ;
        RECT 1450.790 -4.800 1451.350 1.630 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.430 400.250 650.710 404.000 ;
        RECT 649.680 400.110 650.710 400.250 ;
        RECT 649.680 65.125 649.820 400.110 ;
        RECT 650.430 400.000 650.710 400.110 ;
        RECT 649.610 64.755 649.890 65.125 ;
        RECT 1466.110 64.755 1466.390 65.125 ;
        RECT 1466.180 1.770 1466.320 64.755 ;
        RECT 1468.270 1.770 1468.830 2.400 ;
        RECT 1466.180 1.630 1468.830 1.770 ;
        RECT 1468.270 -4.800 1468.830 1.630 ;
      LAYER via2 ;
        RECT 649.610 64.800 649.890 65.080 ;
        RECT 1466.110 64.800 1466.390 65.080 ;
      LAYER met3 ;
        RECT 649.585 65.090 649.915 65.105 ;
        RECT 1466.085 65.090 1466.415 65.105 ;
        RECT 649.585 64.790 1466.415 65.090 ;
        RECT 649.585 64.775 649.915 64.790 ;
        RECT 1466.085 64.775 1466.415 64.790 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 655.570 386.480 655.890 386.540 ;
        RECT 656.950 386.480 657.270 386.540 ;
        RECT 655.570 386.340 657.270 386.480 ;
        RECT 655.570 386.280 655.890 386.340 ;
        RECT 656.950 386.280 657.270 386.340 ;
        RECT 656.950 113.120 657.270 113.180 ;
        RECT 1483.570 113.120 1483.890 113.180 ;
        RECT 656.950 112.980 1483.890 113.120 ;
        RECT 656.950 112.920 657.270 112.980 ;
        RECT 1483.570 112.920 1483.890 112.980 ;
      LAYER via ;
        RECT 655.600 386.280 655.860 386.540 ;
        RECT 656.980 386.280 657.240 386.540 ;
        RECT 656.980 112.920 657.240 113.180 ;
        RECT 1483.600 112.920 1483.860 113.180 ;
      LAYER met2 ;
        RECT 655.950 400.250 656.230 404.000 ;
        RECT 655.660 400.110 656.230 400.250 ;
        RECT 655.660 386.570 655.800 400.110 ;
        RECT 655.950 400.000 656.230 400.110 ;
        RECT 655.600 386.250 655.860 386.570 ;
        RECT 656.980 386.250 657.240 386.570 ;
        RECT 657.040 113.210 657.180 386.250 ;
        RECT 656.980 112.890 657.240 113.210 ;
        RECT 1483.600 112.890 1483.860 113.210 ;
        RECT 1483.660 82.870 1483.800 112.890 ;
        RECT 1483.660 82.730 1486.560 82.870 ;
        RECT 1486.420 2.400 1486.560 82.730 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.490 386.140 656.810 386.200 ;
        RECT 660.170 386.140 660.490 386.200 ;
        RECT 656.490 386.000 660.490 386.140 ;
        RECT 656.490 385.940 656.810 386.000 ;
        RECT 660.170 385.940 660.490 386.000 ;
        RECT 656.490 113.460 656.810 113.520 ;
        RECT 1497.370 113.460 1497.690 113.520 ;
        RECT 656.490 113.320 1497.690 113.460 ;
        RECT 656.490 113.260 656.810 113.320 ;
        RECT 1497.370 113.260 1497.690 113.320 ;
        RECT 1497.370 15.200 1497.690 15.260 ;
        RECT 1503.810 15.200 1504.130 15.260 ;
        RECT 1497.370 15.060 1504.130 15.200 ;
        RECT 1497.370 15.000 1497.690 15.060 ;
        RECT 1503.810 15.000 1504.130 15.060 ;
      LAYER via ;
        RECT 656.520 385.940 656.780 386.200 ;
        RECT 660.200 385.940 660.460 386.200 ;
        RECT 656.520 113.260 656.780 113.520 ;
        RECT 1497.400 113.260 1497.660 113.520 ;
        RECT 1497.400 15.000 1497.660 15.260 ;
        RECT 1503.840 15.000 1504.100 15.260 ;
      LAYER met2 ;
        RECT 661.470 400.250 661.750 404.000 ;
        RECT 660.260 400.110 661.750 400.250 ;
        RECT 660.260 386.230 660.400 400.110 ;
        RECT 661.470 400.000 661.750 400.110 ;
        RECT 656.520 385.910 656.780 386.230 ;
        RECT 660.200 385.910 660.460 386.230 ;
        RECT 656.580 113.550 656.720 385.910 ;
        RECT 656.520 113.230 656.780 113.550 ;
        RECT 1497.400 113.230 1497.660 113.550 ;
        RECT 1497.460 15.290 1497.600 113.230 ;
        RECT 1497.400 14.970 1497.660 15.290 ;
        RECT 1503.840 14.970 1504.100 15.290 ;
        RECT 1503.900 2.400 1504.040 14.970 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 415.450 37.980 415.770 38.040 ;
        RECT 706.170 37.980 706.490 38.040 ;
        RECT 415.450 37.840 706.490 37.980 ;
        RECT 415.450 37.780 415.770 37.840 ;
        RECT 706.170 37.780 706.490 37.840 ;
      LAYER via ;
        RECT 415.480 37.780 415.740 38.040 ;
        RECT 706.200 37.780 706.460 38.040 ;
      LAYER met2 ;
        RECT 416.290 400.250 416.570 404.000 ;
        RECT 415.540 400.110 416.570 400.250 ;
        RECT 415.540 38.070 415.680 400.110 ;
        RECT 416.290 400.000 416.570 400.110 ;
        RECT 415.480 37.750 415.740 38.070 ;
        RECT 706.200 37.750 706.460 38.070 ;
        RECT 706.260 2.400 706.400 37.750 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.850 118.900 664.170 118.960 ;
        RECT 1518.070 118.900 1518.390 118.960 ;
        RECT 663.850 118.760 1518.390 118.900 ;
        RECT 663.850 118.700 664.170 118.760 ;
        RECT 1518.070 118.700 1518.390 118.760 ;
      LAYER via ;
        RECT 663.880 118.700 664.140 118.960 ;
        RECT 1518.100 118.700 1518.360 118.960 ;
      LAYER met2 ;
        RECT 666.990 400.250 667.270 404.000 ;
        RECT 665.780 400.110 667.270 400.250 ;
        RECT 665.780 386.650 665.920 400.110 ;
        RECT 666.990 400.000 667.270 400.110 ;
        RECT 663.940 386.510 665.920 386.650 ;
        RECT 663.940 118.990 664.080 386.510 ;
        RECT 663.880 118.670 664.140 118.990 ;
        RECT 1518.100 118.670 1518.360 118.990 ;
        RECT 1518.160 82.870 1518.300 118.670 ;
        RECT 1518.160 82.730 1519.680 82.870 ;
        RECT 1519.540 1.770 1519.680 82.730 ;
        RECT 1521.630 1.770 1522.190 2.400 ;
        RECT 1519.540 1.630 1522.190 1.770 ;
        RECT 1521.630 -4.800 1522.190 1.630 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.750 119.240 671.070 119.300 ;
        RECT 1538.770 119.240 1539.090 119.300 ;
        RECT 670.750 119.100 1539.090 119.240 ;
        RECT 670.750 119.040 671.070 119.100 ;
        RECT 1538.770 119.040 1539.090 119.100 ;
      LAYER via ;
        RECT 670.780 119.040 671.040 119.300 ;
        RECT 1538.800 119.040 1539.060 119.300 ;
      LAYER met2 ;
        RECT 672.050 400.250 672.330 404.000 ;
        RECT 670.840 400.110 672.330 400.250 ;
        RECT 670.840 119.330 670.980 400.110 ;
        RECT 672.050 400.000 672.330 400.110 ;
        RECT 670.780 119.010 671.040 119.330 ;
        RECT 1538.800 119.010 1539.060 119.330 ;
        RECT 1538.860 17.410 1539.000 119.010 ;
        RECT 1538.860 17.270 1539.920 17.410 ;
        RECT 1539.780 2.400 1539.920 17.270 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 677.190 119.580 677.510 119.640 ;
        RECT 1552.570 119.580 1552.890 119.640 ;
        RECT 677.190 119.440 1552.890 119.580 ;
        RECT 677.190 119.380 677.510 119.440 ;
        RECT 1552.570 119.380 1552.890 119.440 ;
      LAYER via ;
        RECT 677.220 119.380 677.480 119.640 ;
        RECT 1552.600 119.380 1552.860 119.640 ;
      LAYER met2 ;
        RECT 677.570 400.180 677.850 404.000 ;
        RECT 677.570 400.000 677.880 400.180 ;
        RECT 677.740 373.050 677.880 400.000 ;
        RECT 677.280 372.910 677.880 373.050 ;
        RECT 677.280 119.670 677.420 372.910 ;
        RECT 677.220 119.350 677.480 119.670 ;
        RECT 1552.600 119.350 1552.860 119.670 ;
        RECT 1552.660 82.870 1552.800 119.350 ;
        RECT 1552.660 82.730 1557.400 82.870 ;
        RECT 1557.260 2.400 1557.400 82.730 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 683.630 70.620 683.950 70.680 ;
        RECT 1573.270 70.620 1573.590 70.680 ;
        RECT 683.630 70.480 1573.590 70.620 ;
        RECT 683.630 70.420 683.950 70.480 ;
        RECT 1573.270 70.420 1573.590 70.480 ;
      LAYER via ;
        RECT 683.660 70.420 683.920 70.680 ;
        RECT 1573.300 70.420 1573.560 70.680 ;
      LAYER met2 ;
        RECT 683.090 400.250 683.370 404.000 ;
        RECT 683.090 400.110 683.860 400.250 ;
        RECT 683.090 400.000 683.370 400.110 ;
        RECT 683.720 70.710 683.860 400.110 ;
        RECT 683.660 70.390 683.920 70.710 ;
        RECT 1573.300 70.390 1573.560 70.710 ;
        RECT 1573.360 1.770 1573.500 70.390 ;
        RECT 1574.990 1.770 1575.550 2.400 ;
        RECT 1573.360 1.630 1575.550 1.770 ;
        RECT 1574.990 -4.800 1575.550 1.630 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 684.090 386.480 684.410 386.540 ;
        RECT 687.310 386.480 687.630 386.540 ;
        RECT 684.090 386.340 687.630 386.480 ;
        RECT 684.090 386.280 684.410 386.340 ;
        RECT 687.310 386.280 687.630 386.340 ;
        RECT 684.090 70.960 684.410 71.020 ;
        RECT 1590.290 70.960 1590.610 71.020 ;
        RECT 684.090 70.820 1590.610 70.960 ;
        RECT 684.090 70.760 684.410 70.820 ;
        RECT 1590.290 70.760 1590.610 70.820 ;
      LAYER via ;
        RECT 684.120 386.280 684.380 386.540 ;
        RECT 687.340 386.280 687.600 386.540 ;
        RECT 684.120 70.760 684.380 71.020 ;
        RECT 1590.320 70.760 1590.580 71.020 ;
      LAYER met2 ;
        RECT 688.610 400.250 688.890 404.000 ;
        RECT 687.400 400.110 688.890 400.250 ;
        RECT 687.400 386.570 687.540 400.110 ;
        RECT 688.610 400.000 688.890 400.110 ;
        RECT 684.120 386.250 684.380 386.570 ;
        RECT 687.340 386.250 687.600 386.570 ;
        RECT 684.180 71.050 684.320 386.250 ;
        RECT 684.120 70.730 684.380 71.050 ;
        RECT 1590.320 70.730 1590.580 71.050 ;
        RECT 1590.380 1.770 1590.520 70.730 ;
        RECT 1592.470 1.770 1593.030 2.400 ;
        RECT 1590.380 1.630 1593.030 1.770 ;
        RECT 1592.470 -4.800 1593.030 1.630 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.530 386.820 690.850 386.880 ;
        RECT 692.830 386.820 693.150 386.880 ;
        RECT 690.530 386.680 693.150 386.820 ;
        RECT 690.530 386.620 690.850 386.680 ;
        RECT 692.830 386.620 693.150 386.680 ;
        RECT 690.530 71.300 690.850 71.360 ;
        RECT 1610.530 71.300 1610.850 71.360 ;
        RECT 690.530 71.160 1610.850 71.300 ;
        RECT 690.530 71.100 690.850 71.160 ;
        RECT 1610.530 71.100 1610.850 71.160 ;
      LAYER via ;
        RECT 690.560 386.620 690.820 386.880 ;
        RECT 692.860 386.620 693.120 386.880 ;
        RECT 690.560 71.100 690.820 71.360 ;
        RECT 1610.560 71.100 1610.820 71.360 ;
      LAYER met2 ;
        RECT 694.130 400.250 694.410 404.000 ;
        RECT 692.920 400.110 694.410 400.250 ;
        RECT 692.920 386.910 693.060 400.110 ;
        RECT 694.130 400.000 694.410 400.110 ;
        RECT 690.560 386.590 690.820 386.910 ;
        RECT 692.860 386.590 693.120 386.910 ;
        RECT 690.620 71.390 690.760 386.590 ;
        RECT 690.560 71.070 690.820 71.390 ;
        RECT 1610.560 71.070 1610.820 71.390 ;
        RECT 1610.620 2.400 1610.760 71.070 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 697.890 71.640 698.210 71.700 ;
        RECT 1621.570 71.640 1621.890 71.700 ;
        RECT 697.890 71.500 1621.890 71.640 ;
        RECT 697.890 71.440 698.210 71.500 ;
        RECT 1621.570 71.440 1621.890 71.500 ;
        RECT 1621.570 15.200 1621.890 15.260 ;
        RECT 1628.010 15.200 1628.330 15.260 ;
        RECT 1621.570 15.060 1628.330 15.200 ;
        RECT 1621.570 15.000 1621.890 15.060 ;
        RECT 1628.010 15.000 1628.330 15.060 ;
      LAYER via ;
        RECT 697.920 71.440 698.180 71.700 ;
        RECT 1621.600 71.440 1621.860 71.700 ;
        RECT 1621.600 15.000 1621.860 15.260 ;
        RECT 1628.040 15.000 1628.300 15.260 ;
      LAYER met2 ;
        RECT 699.650 400.250 699.930 404.000 ;
        RECT 698.440 400.110 699.930 400.250 ;
        RECT 698.440 386.650 698.580 400.110 ;
        RECT 699.650 400.000 699.930 400.110 ;
        RECT 697.980 386.510 698.580 386.650 ;
        RECT 697.980 71.730 698.120 386.510 ;
        RECT 697.920 71.410 698.180 71.730 ;
        RECT 1621.600 71.410 1621.860 71.730 ;
        RECT 1621.660 15.290 1621.800 71.410 ;
        RECT 1621.600 14.970 1621.860 15.290 ;
        RECT 1628.040 14.970 1628.300 15.290 ;
        RECT 1628.100 2.400 1628.240 14.970 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.330 71.980 704.650 72.040 ;
        RECT 1643.650 71.980 1643.970 72.040 ;
        RECT 704.330 71.840 1643.970 71.980 ;
        RECT 704.330 71.780 704.650 71.840 ;
        RECT 1643.650 71.780 1643.970 71.840 ;
      LAYER via ;
        RECT 704.360 71.780 704.620 72.040 ;
        RECT 1643.680 71.780 1643.940 72.040 ;
      LAYER met2 ;
        RECT 704.710 400.250 704.990 404.000 ;
        RECT 704.420 400.110 704.990 400.250 ;
        RECT 704.420 72.070 704.560 400.110 ;
        RECT 704.710 400.000 704.990 400.110 ;
        RECT 704.360 71.750 704.620 72.070 ;
        RECT 1643.680 71.750 1643.940 72.070 ;
        RECT 1643.740 1.770 1643.880 71.750 ;
        RECT 1645.830 1.770 1646.390 2.400 ;
        RECT 1643.740 1.630 1646.390 1.770 ;
        RECT 1645.830 -4.800 1646.390 1.630 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 704.790 386.480 705.110 386.540 ;
        RECT 708.930 386.480 709.250 386.540 ;
        RECT 704.790 386.340 709.250 386.480 ;
        RECT 704.790 386.280 705.110 386.340 ;
        RECT 708.930 386.280 709.250 386.340 ;
        RECT 704.790 75.720 705.110 75.780 ;
        RECT 1663.430 75.720 1663.750 75.780 ;
        RECT 704.790 75.580 1663.750 75.720 ;
        RECT 704.790 75.520 705.110 75.580 ;
        RECT 1663.430 75.520 1663.750 75.580 ;
      LAYER via ;
        RECT 704.820 386.280 705.080 386.540 ;
        RECT 708.960 386.280 709.220 386.540 ;
        RECT 704.820 75.520 705.080 75.780 ;
        RECT 1663.460 75.520 1663.720 75.780 ;
      LAYER met2 ;
        RECT 710.230 400.250 710.510 404.000 ;
        RECT 709.020 400.110 710.510 400.250 ;
        RECT 709.020 386.570 709.160 400.110 ;
        RECT 710.230 400.000 710.510 400.110 ;
        RECT 704.820 386.250 705.080 386.570 ;
        RECT 708.960 386.250 709.220 386.570 ;
        RECT 704.880 75.810 705.020 386.250 ;
        RECT 704.820 75.490 705.080 75.810 ;
        RECT 1663.460 75.490 1663.720 75.810 ;
        RECT 1663.520 2.400 1663.660 75.490 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.230 386.140 711.550 386.200 ;
        RECT 714.450 386.140 714.770 386.200 ;
        RECT 711.230 386.000 714.770 386.140 ;
        RECT 711.230 385.940 711.550 386.000 ;
        RECT 714.450 385.940 714.770 386.000 ;
        RECT 711.230 75.380 711.550 75.440 ;
        RECT 1681.370 75.380 1681.690 75.440 ;
        RECT 711.230 75.240 1681.690 75.380 ;
        RECT 711.230 75.180 711.550 75.240 ;
        RECT 1681.370 75.180 1681.690 75.240 ;
      LAYER via ;
        RECT 711.260 385.940 711.520 386.200 ;
        RECT 714.480 385.940 714.740 386.200 ;
        RECT 711.260 75.180 711.520 75.440 ;
        RECT 1681.400 75.180 1681.660 75.440 ;
      LAYER met2 ;
        RECT 715.750 400.250 716.030 404.000 ;
        RECT 714.540 400.110 716.030 400.250 ;
        RECT 714.540 386.230 714.680 400.110 ;
        RECT 715.750 400.000 716.030 400.110 ;
        RECT 711.260 385.910 711.520 386.230 ;
        RECT 714.480 385.910 714.740 386.230 ;
        RECT 711.320 75.470 711.460 385.910 ;
        RECT 711.260 75.150 711.520 75.470 ;
        RECT 1681.400 75.150 1681.660 75.470 ;
        RECT 1681.460 2.400 1681.600 75.150 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.890 35.940 422.210 36.000 ;
        RECT 723.650 35.940 723.970 36.000 ;
        RECT 421.890 35.800 723.970 35.940 ;
        RECT 421.890 35.740 422.210 35.800 ;
        RECT 723.650 35.740 723.970 35.800 ;
      LAYER via ;
        RECT 421.920 35.740 422.180 36.000 ;
        RECT 723.680 35.740 723.940 36.000 ;
      LAYER met2 ;
        RECT 421.810 400.180 422.090 404.000 ;
        RECT 421.810 400.000 422.120 400.180 ;
        RECT 421.980 36.030 422.120 400.000 ;
        RECT 421.920 35.710 422.180 36.030 ;
        RECT 723.680 35.710 723.940 36.030 ;
        RECT 723.740 2.400 723.880 35.710 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.130 385.800 718.450 385.860 ;
        RECT 719.970 385.800 720.290 385.860 ;
        RECT 718.130 385.660 720.290 385.800 ;
        RECT 718.130 385.600 718.450 385.660 ;
        RECT 719.970 385.600 720.290 385.660 ;
        RECT 718.130 75.040 718.450 75.100 ;
        RECT 1697.470 75.040 1697.790 75.100 ;
        RECT 718.130 74.900 1697.790 75.040 ;
        RECT 718.130 74.840 718.450 74.900 ;
        RECT 1697.470 74.840 1697.790 74.900 ;
      LAYER via ;
        RECT 718.160 385.600 718.420 385.860 ;
        RECT 720.000 385.600 720.260 385.860 ;
        RECT 718.160 74.840 718.420 75.100 ;
        RECT 1697.500 74.840 1697.760 75.100 ;
      LAYER met2 ;
        RECT 721.270 400.250 721.550 404.000 ;
        RECT 720.060 400.110 721.550 400.250 ;
        RECT 720.060 385.890 720.200 400.110 ;
        RECT 721.270 400.000 721.550 400.110 ;
        RECT 718.160 385.570 718.420 385.890 ;
        RECT 720.000 385.570 720.260 385.890 ;
        RECT 718.220 75.130 718.360 385.570 ;
        RECT 718.160 74.810 718.420 75.130 ;
        RECT 1697.500 74.810 1697.760 75.130 ;
        RECT 1697.560 1.770 1697.700 74.810 ;
        RECT 1699.190 1.770 1699.750 2.400 ;
        RECT 1697.560 1.630 1699.750 1.770 ;
        RECT 1699.190 -4.800 1699.750 1.630 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.030 74.700 725.350 74.760 ;
        RECT 1714.490 74.700 1714.810 74.760 ;
        RECT 725.030 74.560 1714.810 74.700 ;
        RECT 725.030 74.500 725.350 74.560 ;
        RECT 1714.490 74.500 1714.810 74.560 ;
      LAYER via ;
        RECT 725.060 74.500 725.320 74.760 ;
        RECT 1714.520 74.500 1714.780 74.760 ;
      LAYER met2 ;
        RECT 726.790 400.250 727.070 404.000 ;
        RECT 725.580 400.110 727.070 400.250 ;
        RECT 725.580 386.480 725.720 400.110 ;
        RECT 726.790 400.000 727.070 400.110 ;
        RECT 725.120 386.340 725.720 386.480 ;
        RECT 725.120 74.790 725.260 386.340 ;
        RECT 725.060 74.470 725.320 74.790 ;
        RECT 1714.520 74.470 1714.780 74.790 ;
        RECT 1714.580 1.770 1714.720 74.470 ;
        RECT 1716.670 1.770 1717.230 2.400 ;
        RECT 1714.580 1.630 1717.230 1.770 ;
        RECT 1716.670 -4.800 1717.230 1.630 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.930 74.360 732.250 74.420 ;
        RECT 1734.730 74.360 1735.050 74.420 ;
        RECT 731.930 74.220 1735.050 74.360 ;
        RECT 731.930 74.160 732.250 74.220 ;
        RECT 1734.730 74.160 1735.050 74.220 ;
      LAYER via ;
        RECT 731.960 74.160 732.220 74.420 ;
        RECT 1734.760 74.160 1735.020 74.420 ;
      LAYER met2 ;
        RECT 732.310 400.250 732.590 404.000 ;
        RECT 732.020 400.110 732.590 400.250 ;
        RECT 732.020 74.450 732.160 400.110 ;
        RECT 732.310 400.000 732.590 400.110 ;
        RECT 731.960 74.130 732.220 74.450 ;
        RECT 1734.760 74.130 1735.020 74.450 ;
        RECT 1734.820 2.400 1734.960 74.130 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 731.470 386.140 731.790 386.200 ;
        RECT 736.070 386.140 736.390 386.200 ;
        RECT 731.470 386.000 736.390 386.140 ;
        RECT 731.470 385.940 731.790 386.000 ;
        RECT 736.070 385.940 736.390 386.000 ;
        RECT 731.470 74.020 731.790 74.080 ;
        RECT 1746.230 74.020 1746.550 74.080 ;
        RECT 731.470 73.880 1746.550 74.020 ;
        RECT 731.470 73.820 731.790 73.880 ;
        RECT 1746.230 73.820 1746.550 73.880 ;
        RECT 1746.230 15.200 1746.550 15.260 ;
        RECT 1752.210 15.200 1752.530 15.260 ;
        RECT 1746.230 15.060 1752.530 15.200 ;
        RECT 1746.230 15.000 1746.550 15.060 ;
        RECT 1752.210 15.000 1752.530 15.060 ;
      LAYER via ;
        RECT 731.500 385.940 731.760 386.200 ;
        RECT 736.100 385.940 736.360 386.200 ;
        RECT 731.500 73.820 731.760 74.080 ;
        RECT 1746.260 73.820 1746.520 74.080 ;
        RECT 1746.260 15.000 1746.520 15.260 ;
        RECT 1752.240 15.000 1752.500 15.260 ;
      LAYER met2 ;
        RECT 737.370 400.250 737.650 404.000 ;
        RECT 736.160 400.110 737.650 400.250 ;
        RECT 736.160 386.230 736.300 400.110 ;
        RECT 737.370 400.000 737.650 400.110 ;
        RECT 731.500 385.910 731.760 386.230 ;
        RECT 736.100 385.910 736.360 386.230 ;
        RECT 731.560 74.110 731.700 385.910 ;
        RECT 731.500 73.790 731.760 74.110 ;
        RECT 1746.260 73.790 1746.520 74.110 ;
        RECT 1746.320 15.290 1746.460 73.790 ;
        RECT 1746.260 14.970 1746.520 15.290 ;
        RECT 1752.240 14.970 1752.500 15.290 ;
        RECT 1752.300 2.400 1752.440 14.970 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 738.370 386.140 738.690 386.200 ;
        RECT 741.590 386.140 741.910 386.200 ;
        RECT 738.370 386.000 741.910 386.140 ;
        RECT 738.370 385.940 738.690 386.000 ;
        RECT 741.590 385.940 741.910 386.000 ;
        RECT 738.370 73.680 738.690 73.740 ;
        RECT 1767.850 73.680 1768.170 73.740 ;
        RECT 738.370 73.540 1768.170 73.680 ;
        RECT 738.370 73.480 738.690 73.540 ;
        RECT 1767.850 73.480 1768.170 73.540 ;
      LAYER via ;
        RECT 738.400 385.940 738.660 386.200 ;
        RECT 741.620 385.940 741.880 386.200 ;
        RECT 738.400 73.480 738.660 73.740 ;
        RECT 1767.880 73.480 1768.140 73.740 ;
      LAYER met2 ;
        RECT 742.890 400.250 743.170 404.000 ;
        RECT 741.680 400.110 743.170 400.250 ;
        RECT 741.680 386.230 741.820 400.110 ;
        RECT 742.890 400.000 743.170 400.110 ;
        RECT 738.400 385.910 738.660 386.230 ;
        RECT 741.620 385.910 741.880 386.230 ;
        RECT 738.460 73.770 738.600 385.910 ;
        RECT 738.400 73.450 738.660 73.770 ;
        RECT 1767.880 73.450 1768.140 73.770 ;
        RECT 1767.940 1.770 1768.080 73.450 ;
        RECT 1770.030 1.770 1770.590 2.400 ;
        RECT 1767.940 1.630 1770.590 1.770 ;
        RECT 1770.030 -4.800 1770.590 1.630 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 745.270 387.160 745.590 387.220 ;
        RECT 747.110 387.160 747.430 387.220 ;
        RECT 745.270 387.020 747.430 387.160 ;
        RECT 745.270 386.960 745.590 387.020 ;
        RECT 747.110 386.960 747.430 387.020 ;
        RECT 745.270 73.340 745.590 73.400 ;
        RECT 1787.630 73.340 1787.950 73.400 ;
        RECT 745.270 73.200 1787.950 73.340 ;
        RECT 745.270 73.140 745.590 73.200 ;
        RECT 1787.630 73.140 1787.950 73.200 ;
      LAYER via ;
        RECT 745.300 386.960 745.560 387.220 ;
        RECT 747.140 386.960 747.400 387.220 ;
        RECT 745.300 73.140 745.560 73.400 ;
        RECT 1787.660 73.140 1787.920 73.400 ;
      LAYER met2 ;
        RECT 748.410 400.250 748.690 404.000 ;
        RECT 747.200 400.110 748.690 400.250 ;
        RECT 747.200 387.250 747.340 400.110 ;
        RECT 748.410 400.000 748.690 400.110 ;
        RECT 745.300 386.930 745.560 387.250 ;
        RECT 747.140 386.930 747.400 387.250 ;
        RECT 745.360 73.430 745.500 386.930 ;
        RECT 745.300 73.110 745.560 73.430 ;
        RECT 1787.660 73.110 1787.920 73.430 ;
        RECT 1787.720 2.400 1787.860 73.110 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.630 73.000 752.950 73.060 ;
        RECT 1805.570 73.000 1805.890 73.060 ;
        RECT 752.630 72.860 1805.890 73.000 ;
        RECT 752.630 72.800 752.950 72.860 ;
        RECT 1805.570 72.800 1805.890 72.860 ;
      LAYER via ;
        RECT 752.660 72.800 752.920 73.060 ;
        RECT 1805.600 72.800 1805.860 73.060 ;
      LAYER met2 ;
        RECT 753.930 400.930 754.210 404.000 ;
        RECT 752.720 400.790 754.210 400.930 ;
        RECT 752.720 73.090 752.860 400.790 ;
        RECT 753.930 400.000 754.210 400.790 ;
        RECT 752.660 72.770 752.920 73.090 ;
        RECT 1805.600 72.770 1805.860 73.090 ;
        RECT 1805.660 2.400 1805.800 72.770 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.990 72.660 760.310 72.720 ;
        RECT 1823.050 72.660 1823.370 72.720 ;
        RECT 759.990 72.520 1823.370 72.660 ;
        RECT 759.990 72.460 760.310 72.520 ;
        RECT 1823.050 72.460 1823.370 72.520 ;
      LAYER via ;
        RECT 760.020 72.460 760.280 72.720 ;
        RECT 1823.080 72.460 1823.340 72.720 ;
      LAYER met2 ;
        RECT 759.450 400.250 759.730 404.000 ;
        RECT 759.450 400.110 760.220 400.250 ;
        RECT 759.450 400.000 759.730 400.110 ;
        RECT 760.080 72.750 760.220 400.110 ;
        RECT 760.020 72.430 760.280 72.750 ;
        RECT 1823.080 72.430 1823.340 72.750 ;
        RECT 1823.140 2.400 1823.280 72.430 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 759.530 386.140 759.850 386.200 ;
        RECT 763.670 386.140 763.990 386.200 ;
        RECT 759.530 386.000 763.990 386.140 ;
        RECT 759.530 385.940 759.850 386.000 ;
        RECT 763.670 385.940 763.990 386.000 ;
        RECT 759.530 72.320 759.850 72.380 ;
        RECT 1838.690 72.320 1839.010 72.380 ;
        RECT 759.530 72.180 1839.010 72.320 ;
        RECT 759.530 72.120 759.850 72.180 ;
        RECT 1838.690 72.120 1839.010 72.180 ;
      LAYER via ;
        RECT 759.560 385.940 759.820 386.200 ;
        RECT 763.700 385.940 763.960 386.200 ;
        RECT 759.560 72.120 759.820 72.380 ;
        RECT 1838.720 72.120 1838.980 72.380 ;
      LAYER met2 ;
        RECT 764.970 400.250 765.250 404.000 ;
        RECT 763.760 400.110 765.250 400.250 ;
        RECT 763.760 386.230 763.900 400.110 ;
        RECT 764.970 400.000 765.250 400.110 ;
        RECT 759.560 385.910 759.820 386.230 ;
        RECT 763.700 385.910 763.960 386.230 ;
        RECT 759.620 72.410 759.760 385.910 ;
        RECT 759.560 72.090 759.820 72.410 ;
        RECT 1838.720 72.090 1838.980 72.410 ;
        RECT 1838.780 1.770 1838.920 72.090 ;
        RECT 1840.870 1.770 1841.430 2.400 ;
        RECT 1838.780 1.630 1841.430 1.770 ;
        RECT 1840.870 -4.800 1841.430 1.630 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.030 400.250 770.310 404.000 ;
        RECT 768.820 400.110 770.310 400.250 ;
        RECT 768.820 385.970 768.960 400.110 ;
        RECT 770.030 400.000 770.310 400.110 ;
        RECT 766.520 385.830 768.960 385.970 ;
        RECT 766.520 72.605 766.660 385.830 ;
        RECT 766.450 72.235 766.730 72.605 ;
        RECT 1856.190 72.235 1856.470 72.605 ;
        RECT 1856.260 1.770 1856.400 72.235 ;
        RECT 1858.350 1.770 1858.910 2.400 ;
        RECT 1856.260 1.630 1858.910 1.770 ;
        RECT 1858.350 -4.800 1858.910 1.630 ;
      LAYER via2 ;
        RECT 766.450 72.280 766.730 72.560 ;
        RECT 1856.190 72.280 1856.470 72.560 ;
      LAYER met3 ;
        RECT 766.425 72.570 766.755 72.585 ;
        RECT 1856.165 72.570 1856.495 72.585 ;
        RECT 766.425 72.270 1856.495 72.570 ;
        RECT 766.425 72.255 766.755 72.270 ;
        RECT 1856.165 72.255 1856.495 72.270 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 422.350 46.140 422.670 46.200 ;
        RECT 741.590 46.140 741.910 46.200 ;
        RECT 422.350 46.000 741.910 46.140 ;
        RECT 422.350 45.940 422.670 46.000 ;
        RECT 741.590 45.940 741.910 46.000 ;
      LAYER via ;
        RECT 422.380 45.940 422.640 46.200 ;
        RECT 741.620 45.940 741.880 46.200 ;
      LAYER met2 ;
        RECT 427.330 400.250 427.610 404.000 ;
        RECT 426.120 400.110 427.610 400.250 ;
        RECT 426.120 324.370 426.260 400.110 ;
        RECT 427.330 400.000 427.610 400.110 ;
        RECT 422.440 324.230 426.260 324.370 ;
        RECT 422.440 46.230 422.580 324.230 ;
        RECT 422.380 45.910 422.640 46.230 ;
        RECT 741.620 45.910 741.880 46.230 ;
        RECT 741.680 2.400 741.820 45.910 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 773.790 119.920 774.110 119.980 ;
        RECT 1869.970 119.920 1870.290 119.980 ;
        RECT 773.790 119.780 1870.290 119.920 ;
        RECT 773.790 119.720 774.110 119.780 ;
        RECT 1869.970 119.720 1870.290 119.780 ;
        RECT 1869.970 15.200 1870.290 15.260 ;
        RECT 1876.410 15.200 1876.730 15.260 ;
        RECT 1869.970 15.060 1876.730 15.200 ;
        RECT 1869.970 15.000 1870.290 15.060 ;
        RECT 1876.410 15.000 1876.730 15.060 ;
      LAYER via ;
        RECT 773.820 119.720 774.080 119.980 ;
        RECT 1870.000 119.720 1870.260 119.980 ;
        RECT 1870.000 15.000 1870.260 15.260 ;
        RECT 1876.440 15.000 1876.700 15.260 ;
      LAYER met2 ;
        RECT 775.550 400.250 775.830 404.000 ;
        RECT 774.340 400.110 775.830 400.250 ;
        RECT 774.340 324.370 774.480 400.110 ;
        RECT 775.550 400.000 775.830 400.110 ;
        RECT 773.880 324.230 774.480 324.370 ;
        RECT 773.880 120.010 774.020 324.230 ;
        RECT 773.820 119.690 774.080 120.010 ;
        RECT 1870.000 119.690 1870.260 120.010 ;
        RECT 1870.060 15.290 1870.200 119.690 ;
        RECT 1870.000 14.970 1870.260 15.290 ;
        RECT 1876.440 14.970 1876.700 15.290 ;
        RECT 1876.500 2.400 1876.640 14.970 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.230 120.260 780.550 120.320 ;
        RECT 1890.670 120.260 1890.990 120.320 ;
        RECT 780.230 120.120 1890.990 120.260 ;
        RECT 780.230 120.060 780.550 120.120 ;
        RECT 1890.670 120.060 1890.990 120.120 ;
      LAYER via ;
        RECT 780.260 120.060 780.520 120.320 ;
        RECT 1890.700 120.060 1890.960 120.320 ;
      LAYER met2 ;
        RECT 781.070 400.250 781.350 404.000 ;
        RECT 780.320 400.110 781.350 400.250 ;
        RECT 780.320 120.350 780.460 400.110 ;
        RECT 781.070 400.000 781.350 400.110 ;
        RECT 780.260 120.030 780.520 120.350 ;
        RECT 1890.700 120.030 1890.960 120.350 ;
        RECT 1890.760 82.870 1890.900 120.030 ;
        RECT 1890.760 82.730 1892.280 82.870 ;
        RECT 1892.140 1.770 1892.280 82.730 ;
        RECT 1894.230 1.770 1894.790 2.400 ;
        RECT 1892.140 1.630 1894.790 1.770 ;
        RECT 1894.230 -4.800 1894.790 1.630 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.130 124.000 787.450 124.060 ;
        RECT 1911.830 124.000 1912.150 124.060 ;
        RECT 787.130 123.860 1912.150 124.000 ;
        RECT 787.130 123.800 787.450 123.860 ;
        RECT 1911.830 123.800 1912.150 123.860 ;
      LAYER via ;
        RECT 787.160 123.800 787.420 124.060 ;
        RECT 1911.860 123.800 1912.120 124.060 ;
      LAYER met2 ;
        RECT 786.590 400.250 786.870 404.000 ;
        RECT 786.590 400.110 787.360 400.250 ;
        RECT 786.590 400.000 786.870 400.110 ;
        RECT 787.220 124.090 787.360 400.110 ;
        RECT 787.160 123.770 787.420 124.090 ;
        RECT 1911.860 123.770 1912.120 124.090 ;
        RECT 1911.920 2.400 1912.060 123.770 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 787.590 123.660 787.910 123.720 ;
        RECT 1925.170 123.660 1925.490 123.720 ;
        RECT 787.590 123.520 1925.490 123.660 ;
        RECT 787.590 123.460 787.910 123.520 ;
        RECT 1925.170 123.460 1925.490 123.520 ;
      LAYER via ;
        RECT 787.620 123.460 787.880 123.720 ;
        RECT 1925.200 123.460 1925.460 123.720 ;
      LAYER met2 ;
        RECT 792.110 400.250 792.390 404.000 ;
        RECT 790.900 400.110 792.390 400.250 ;
        RECT 790.900 324.370 791.040 400.110 ;
        RECT 792.110 400.000 792.390 400.110 ;
        RECT 787.680 324.230 791.040 324.370 ;
        RECT 787.680 123.750 787.820 324.230 ;
        RECT 787.620 123.430 787.880 123.750 ;
        RECT 1925.200 123.430 1925.460 123.750 ;
        RECT 1925.260 82.870 1925.400 123.430 ;
        RECT 1925.260 82.730 1930.000 82.870 ;
        RECT 1929.860 2.400 1930.000 82.730 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.030 376.280 794.350 376.340 ;
        RECT 796.330 376.280 796.650 376.340 ;
        RECT 794.030 376.140 796.650 376.280 ;
        RECT 794.030 376.080 794.350 376.140 ;
        RECT 796.330 376.080 796.650 376.140 ;
        RECT 794.030 123.320 794.350 123.380 ;
        RECT 1945.870 123.320 1946.190 123.380 ;
        RECT 794.030 123.180 1946.190 123.320 ;
        RECT 794.030 123.120 794.350 123.180 ;
        RECT 1945.870 123.120 1946.190 123.180 ;
      LAYER via ;
        RECT 794.060 376.080 794.320 376.340 ;
        RECT 796.360 376.080 796.620 376.340 ;
        RECT 794.060 123.120 794.320 123.380 ;
        RECT 1945.900 123.120 1946.160 123.380 ;
      LAYER met2 ;
        RECT 797.630 400.250 797.910 404.000 ;
        RECT 796.420 400.110 797.910 400.250 ;
        RECT 796.420 376.370 796.560 400.110 ;
        RECT 797.630 400.000 797.910 400.110 ;
        RECT 794.060 376.050 794.320 376.370 ;
        RECT 796.360 376.050 796.620 376.370 ;
        RECT 794.120 123.410 794.260 376.050 ;
        RECT 794.060 123.090 794.320 123.410 ;
        RECT 1945.900 123.090 1946.160 123.410 ;
        RECT 1945.960 82.870 1946.100 123.090 ;
        RECT 1945.960 82.730 1947.480 82.870 ;
        RECT 1947.340 2.400 1947.480 82.730 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 801.390 78.100 801.710 78.160 ;
        RECT 1962.890 78.100 1963.210 78.160 ;
        RECT 801.390 77.960 1963.210 78.100 ;
        RECT 801.390 77.900 801.710 77.960 ;
        RECT 1962.890 77.900 1963.210 77.960 ;
      LAYER via ;
        RECT 801.420 77.900 801.680 78.160 ;
        RECT 1962.920 77.900 1963.180 78.160 ;
      LAYER met2 ;
        RECT 802.690 400.250 802.970 404.000 ;
        RECT 801.480 400.110 802.970 400.250 ;
        RECT 801.480 78.190 801.620 400.110 ;
        RECT 802.690 400.000 802.970 400.110 ;
        RECT 801.420 77.870 801.680 78.190 ;
        RECT 1962.920 77.870 1963.180 78.190 ;
        RECT 1962.980 1.770 1963.120 77.870 ;
        RECT 1965.070 1.770 1965.630 2.400 ;
        RECT 1962.980 1.630 1965.630 1.770 ;
        RECT 1965.070 -4.800 1965.630 1.630 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 808.290 78.440 808.610 78.500 ;
        RECT 1980.370 78.440 1980.690 78.500 ;
        RECT 808.290 78.300 1980.690 78.440 ;
        RECT 808.290 78.240 808.610 78.300 ;
        RECT 1980.370 78.240 1980.690 78.300 ;
      LAYER via ;
        RECT 808.320 78.240 808.580 78.500 ;
        RECT 1980.400 78.240 1980.660 78.500 ;
      LAYER met2 ;
        RECT 808.210 400.180 808.490 404.000 ;
        RECT 808.210 400.000 808.520 400.180 ;
        RECT 808.380 78.530 808.520 400.000 ;
        RECT 808.320 78.210 808.580 78.530 ;
        RECT 1980.400 78.210 1980.660 78.530 ;
        RECT 1980.460 1.770 1980.600 78.210 ;
        RECT 1982.550 1.770 1983.110 2.400 ;
        RECT 1980.460 1.630 1983.110 1.770 ;
        RECT 1982.550 -4.800 1983.110 1.630 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 807.830 375.940 808.150 376.000 ;
        RECT 812.430 375.940 812.750 376.000 ;
        RECT 807.830 375.800 812.750 375.940 ;
        RECT 807.830 375.740 808.150 375.800 ;
        RECT 812.430 375.740 812.750 375.800 ;
        RECT 807.830 78.780 808.150 78.840 ;
        RECT 1994.170 78.780 1994.490 78.840 ;
        RECT 807.830 78.640 1994.490 78.780 ;
        RECT 807.830 78.580 808.150 78.640 ;
        RECT 1994.170 78.580 1994.490 78.640 ;
        RECT 1994.170 15.200 1994.490 15.260 ;
        RECT 2000.610 15.200 2000.930 15.260 ;
        RECT 1994.170 15.060 2000.930 15.200 ;
        RECT 1994.170 15.000 1994.490 15.060 ;
        RECT 2000.610 15.000 2000.930 15.060 ;
      LAYER via ;
        RECT 807.860 375.740 808.120 376.000 ;
        RECT 812.460 375.740 812.720 376.000 ;
        RECT 807.860 78.580 808.120 78.840 ;
        RECT 1994.200 78.580 1994.460 78.840 ;
        RECT 1994.200 15.000 1994.460 15.260 ;
        RECT 2000.640 15.000 2000.900 15.260 ;
      LAYER met2 ;
        RECT 813.730 400.250 814.010 404.000 ;
        RECT 812.520 400.110 814.010 400.250 ;
        RECT 812.520 376.030 812.660 400.110 ;
        RECT 813.730 400.000 814.010 400.110 ;
        RECT 807.860 375.710 808.120 376.030 ;
        RECT 812.460 375.710 812.720 376.030 ;
        RECT 807.920 78.870 808.060 375.710 ;
        RECT 807.860 78.550 808.120 78.870 ;
        RECT 1994.200 78.550 1994.460 78.870 ;
        RECT 1994.260 15.290 1994.400 78.550 ;
        RECT 1994.200 14.970 1994.460 15.290 ;
        RECT 2000.640 14.970 2000.900 15.290 ;
        RECT 2000.700 2.400 2000.840 14.970 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 814.730 376.280 815.050 376.340 ;
        RECT 817.950 376.280 818.270 376.340 ;
        RECT 814.730 376.140 818.270 376.280 ;
        RECT 814.730 376.080 815.050 376.140 ;
        RECT 817.950 376.080 818.270 376.140 ;
        RECT 814.730 79.120 815.050 79.180 ;
        RECT 2018.090 79.120 2018.410 79.180 ;
        RECT 814.730 78.980 2018.410 79.120 ;
        RECT 814.730 78.920 815.050 78.980 ;
        RECT 2018.090 78.920 2018.410 78.980 ;
      LAYER via ;
        RECT 814.760 376.080 815.020 376.340 ;
        RECT 817.980 376.080 818.240 376.340 ;
        RECT 814.760 78.920 815.020 79.180 ;
        RECT 2018.120 78.920 2018.380 79.180 ;
      LAYER met2 ;
        RECT 819.250 400.250 819.530 404.000 ;
        RECT 818.040 400.110 819.530 400.250 ;
        RECT 818.040 376.370 818.180 400.110 ;
        RECT 819.250 400.000 819.530 400.110 ;
        RECT 814.760 376.050 815.020 376.370 ;
        RECT 817.980 376.050 818.240 376.370 ;
        RECT 814.820 79.210 814.960 376.050 ;
        RECT 814.760 78.890 815.020 79.210 ;
        RECT 2018.120 78.890 2018.380 79.210 ;
        RECT 2018.180 2.400 2018.320 78.890 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.630 82.860 821.950 82.920 ;
        RECT 2036.030 82.860 2036.350 82.920 ;
        RECT 821.630 82.720 2036.350 82.860 ;
        RECT 821.630 82.660 821.950 82.720 ;
        RECT 2036.030 82.660 2036.350 82.720 ;
      LAYER via ;
        RECT 821.660 82.660 821.920 82.920 ;
        RECT 2036.060 82.660 2036.320 82.920 ;
      LAYER met2 ;
        RECT 824.770 400.250 825.050 404.000 ;
        RECT 823.560 400.110 825.050 400.250 ;
        RECT 823.560 351.970 823.700 400.110 ;
        RECT 824.770 400.000 825.050 400.110 ;
        RECT 821.720 351.830 823.700 351.970 ;
        RECT 821.720 82.950 821.860 351.830 ;
        RECT 821.660 82.630 821.920 82.950 ;
        RECT 2036.060 82.630 2036.320 82.950 ;
        RECT 2036.120 2.400 2036.260 82.630 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.790 45.800 429.110 45.860 ;
        RECT 759.070 45.800 759.390 45.860 ;
        RECT 428.790 45.660 759.390 45.800 ;
        RECT 428.790 45.600 429.110 45.660 ;
        RECT 759.070 45.600 759.390 45.660 ;
      LAYER via ;
        RECT 428.820 45.600 429.080 45.860 ;
        RECT 759.100 45.600 759.360 45.860 ;
      LAYER met2 ;
        RECT 432.850 400.250 433.130 404.000 ;
        RECT 431.640 400.110 433.130 400.250 ;
        RECT 431.640 386.650 431.780 400.110 ;
        RECT 432.850 400.000 433.130 400.110 ;
        RECT 428.880 386.510 431.780 386.650 ;
        RECT 428.880 45.890 429.020 386.510 ;
        RECT 428.820 45.570 429.080 45.890 ;
        RECT 759.100 45.570 759.360 45.890 ;
        RECT 759.160 2.400 759.300 45.570 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 828.990 82.520 829.310 82.580 ;
        RECT 2053.970 82.520 2054.290 82.580 ;
        RECT 828.990 82.380 2054.290 82.520 ;
        RECT 828.990 82.320 829.310 82.380 ;
        RECT 2053.970 82.320 2054.290 82.380 ;
      LAYER via ;
        RECT 829.020 82.320 829.280 82.580 ;
        RECT 2054.000 82.320 2054.260 82.580 ;
      LAYER met2 ;
        RECT 830.290 400.250 830.570 404.000 ;
        RECT 829.080 400.110 830.570 400.250 ;
        RECT 829.080 82.610 829.220 400.110 ;
        RECT 830.290 400.000 830.570 400.110 ;
        RECT 829.020 82.290 829.280 82.610 ;
        RECT 2054.000 82.290 2054.260 82.610 ;
        RECT 2054.060 2.400 2054.200 82.290 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.430 82.180 835.750 82.240 ;
        RECT 2071.450 82.180 2071.770 82.240 ;
        RECT 835.430 82.040 2071.770 82.180 ;
        RECT 835.430 81.980 835.750 82.040 ;
        RECT 2071.450 81.980 2071.770 82.040 ;
      LAYER via ;
        RECT 835.460 81.980 835.720 82.240 ;
        RECT 2071.480 81.980 2071.740 82.240 ;
      LAYER met2 ;
        RECT 835.350 400.180 835.630 404.000 ;
        RECT 835.350 400.000 835.660 400.180 ;
        RECT 835.520 82.270 835.660 400.000 ;
        RECT 835.460 81.950 835.720 82.270 ;
        RECT 2071.480 81.950 2071.740 82.270 ;
        RECT 2071.540 2.400 2071.680 81.950 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 835.890 376.280 836.210 376.340 ;
        RECT 839.570 376.280 839.890 376.340 ;
        RECT 835.890 376.140 839.890 376.280 ;
        RECT 835.890 376.080 836.210 376.140 ;
        RECT 839.570 376.080 839.890 376.140 ;
        RECT 835.890 81.840 836.210 81.900 ;
        RECT 2087.090 81.840 2087.410 81.900 ;
        RECT 835.890 81.700 2087.410 81.840 ;
        RECT 835.890 81.640 836.210 81.700 ;
        RECT 2087.090 81.640 2087.410 81.700 ;
      LAYER via ;
        RECT 835.920 376.080 836.180 376.340 ;
        RECT 839.600 376.080 839.860 376.340 ;
        RECT 835.920 81.640 836.180 81.900 ;
        RECT 2087.120 81.640 2087.380 81.900 ;
      LAYER met2 ;
        RECT 840.870 400.250 841.150 404.000 ;
        RECT 839.660 400.110 841.150 400.250 ;
        RECT 839.660 376.370 839.800 400.110 ;
        RECT 840.870 400.000 841.150 400.110 ;
        RECT 835.920 376.050 836.180 376.370 ;
        RECT 839.600 376.050 839.860 376.370 ;
        RECT 835.980 81.930 836.120 376.050 ;
        RECT 835.920 81.610 836.180 81.930 ;
        RECT 2087.120 81.610 2087.380 81.930 ;
        RECT 2087.180 1.770 2087.320 81.610 ;
        RECT 2089.270 1.770 2089.830 2.400 ;
        RECT 2087.180 1.630 2089.830 1.770 ;
        RECT 2089.270 -4.800 2089.830 1.630 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.330 81.500 842.650 81.560 ;
        RECT 2104.570 81.500 2104.890 81.560 ;
        RECT 842.330 81.360 2104.890 81.500 ;
        RECT 842.330 81.300 842.650 81.360 ;
        RECT 2104.570 81.300 2104.890 81.360 ;
      LAYER via ;
        RECT 842.360 81.300 842.620 81.560 ;
        RECT 2104.600 81.300 2104.860 81.560 ;
      LAYER met2 ;
        RECT 846.390 400.250 846.670 404.000 ;
        RECT 845.180 400.110 846.670 400.250 ;
        RECT 845.180 351.970 845.320 400.110 ;
        RECT 846.390 400.000 846.670 400.110 ;
        RECT 842.420 351.830 845.320 351.970 ;
        RECT 842.420 81.590 842.560 351.830 ;
        RECT 842.360 81.270 842.620 81.590 ;
        RECT 2104.600 81.270 2104.860 81.590 ;
        RECT 2104.660 1.770 2104.800 81.270 ;
        RECT 2106.750 1.770 2107.310 2.400 ;
        RECT 2104.660 1.630 2107.310 1.770 ;
        RECT 2106.750 -4.800 2107.310 1.630 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 848.770 376.280 849.090 376.340 ;
        RECT 850.610 376.280 850.930 376.340 ;
        RECT 848.770 376.140 850.930 376.280 ;
        RECT 848.770 376.080 849.090 376.140 ;
        RECT 850.610 376.080 850.930 376.140 ;
        RECT 848.770 81.160 849.090 81.220 ;
        RECT 2118.830 81.160 2119.150 81.220 ;
        RECT 848.770 81.020 2119.150 81.160 ;
        RECT 848.770 80.960 849.090 81.020 ;
        RECT 2118.830 80.960 2119.150 81.020 ;
        RECT 2118.830 15.540 2119.150 15.600 ;
        RECT 2124.810 15.540 2125.130 15.600 ;
        RECT 2118.830 15.400 2125.130 15.540 ;
        RECT 2118.830 15.340 2119.150 15.400 ;
        RECT 2124.810 15.340 2125.130 15.400 ;
      LAYER via ;
        RECT 848.800 376.080 849.060 376.340 ;
        RECT 850.640 376.080 850.900 376.340 ;
        RECT 848.800 80.960 849.060 81.220 ;
        RECT 2118.860 80.960 2119.120 81.220 ;
        RECT 2118.860 15.340 2119.120 15.600 ;
        RECT 2124.840 15.340 2125.100 15.600 ;
      LAYER met2 ;
        RECT 851.910 400.250 852.190 404.000 ;
        RECT 850.700 400.110 852.190 400.250 ;
        RECT 850.700 376.370 850.840 400.110 ;
        RECT 851.910 400.000 852.190 400.110 ;
        RECT 848.800 376.050 849.060 376.370 ;
        RECT 850.640 376.050 850.900 376.370 ;
        RECT 848.860 81.250 849.000 376.050 ;
        RECT 848.800 80.930 849.060 81.250 ;
        RECT 2118.860 80.930 2119.120 81.250 ;
        RECT 2118.920 15.630 2119.060 80.930 ;
        RECT 2118.860 15.310 2119.120 15.630 ;
        RECT 2124.840 15.310 2125.100 15.630 ;
        RECT 2124.900 2.400 2125.040 15.310 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 856.130 80.820 856.450 80.880 ;
        RECT 2142.290 80.820 2142.610 80.880 ;
        RECT 856.130 80.680 2142.610 80.820 ;
        RECT 856.130 80.620 856.450 80.680 ;
        RECT 2142.290 80.620 2142.610 80.680 ;
      LAYER via ;
        RECT 856.160 80.620 856.420 80.880 ;
        RECT 2142.320 80.620 2142.580 80.880 ;
      LAYER met2 ;
        RECT 857.430 400.250 857.710 404.000 ;
        RECT 856.220 400.110 857.710 400.250 ;
        RECT 856.220 80.910 856.360 400.110 ;
        RECT 857.430 400.000 857.710 400.110 ;
        RECT 856.160 80.590 856.420 80.910 ;
        RECT 2142.320 80.590 2142.580 80.910 ;
        RECT 2142.380 2.400 2142.520 80.590 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.490 80.480 863.810 80.540 ;
        RECT 2160.230 80.480 2160.550 80.540 ;
        RECT 863.490 80.340 2160.550 80.480 ;
        RECT 863.490 80.280 863.810 80.340 ;
        RECT 2160.230 80.280 2160.550 80.340 ;
      LAYER via ;
        RECT 863.520 80.280 863.780 80.540 ;
        RECT 2160.260 80.280 2160.520 80.540 ;
      LAYER met2 ;
        RECT 862.950 400.250 863.230 404.000 ;
        RECT 862.660 400.110 863.230 400.250 ;
        RECT 862.660 398.890 862.800 400.110 ;
        RECT 862.950 400.000 863.230 400.110 ;
        RECT 862.660 398.750 863.260 398.890 ;
        RECT 863.120 377.130 863.260 398.750 ;
        RECT 863.120 376.990 863.720 377.130 ;
        RECT 863.580 80.570 863.720 376.990 ;
        RECT 863.520 80.250 863.780 80.570 ;
        RECT 2160.260 80.250 2160.520 80.570 ;
        RECT 2160.320 2.400 2160.460 80.250 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 863.030 376.280 863.350 376.340 ;
        RECT 867.170 376.280 867.490 376.340 ;
        RECT 863.030 376.140 867.490 376.280 ;
        RECT 863.030 376.080 863.350 376.140 ;
        RECT 867.170 376.080 867.490 376.140 ;
        RECT 863.030 80.140 863.350 80.200 ;
        RECT 2175.410 80.140 2175.730 80.200 ;
        RECT 863.030 80.000 2175.730 80.140 ;
        RECT 863.030 79.940 863.350 80.000 ;
        RECT 2175.410 79.940 2175.730 80.000 ;
      LAYER via ;
        RECT 863.060 376.080 863.320 376.340 ;
        RECT 867.200 376.080 867.460 376.340 ;
        RECT 863.060 79.940 863.320 80.200 ;
        RECT 2175.440 79.940 2175.700 80.200 ;
      LAYER met2 ;
        RECT 868.010 400.250 868.290 404.000 ;
        RECT 867.260 400.110 868.290 400.250 ;
        RECT 867.260 376.370 867.400 400.110 ;
        RECT 868.010 400.000 868.290 400.110 ;
        RECT 863.060 376.050 863.320 376.370 ;
        RECT 867.200 376.050 867.460 376.370 ;
        RECT 863.120 80.230 863.260 376.050 ;
        RECT 863.060 79.910 863.320 80.230 ;
        RECT 2175.440 79.910 2175.700 80.230 ;
        RECT 2175.500 1.770 2175.640 79.910 ;
        RECT 2177.590 1.770 2178.150 2.400 ;
        RECT 2175.500 1.630 2178.150 1.770 ;
        RECT 2177.590 -4.800 2178.150 1.630 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 870.390 375.940 870.710 376.000 ;
        RECT 872.230 375.940 872.550 376.000 ;
        RECT 870.390 375.800 872.550 375.940 ;
        RECT 870.390 375.740 870.710 375.800 ;
        RECT 872.230 375.740 872.550 375.800 ;
        RECT 870.390 79.800 870.710 79.860 ;
        RECT 2195.650 79.800 2195.970 79.860 ;
        RECT 870.390 79.660 2195.970 79.800 ;
        RECT 870.390 79.600 870.710 79.660 ;
        RECT 2195.650 79.600 2195.970 79.660 ;
      LAYER via ;
        RECT 870.420 375.740 870.680 376.000 ;
        RECT 872.260 375.740 872.520 376.000 ;
        RECT 870.420 79.600 870.680 79.860 ;
        RECT 2195.680 79.600 2195.940 79.860 ;
      LAYER met2 ;
        RECT 873.530 400.250 873.810 404.000 ;
        RECT 872.320 400.110 873.810 400.250 ;
        RECT 872.320 376.030 872.460 400.110 ;
        RECT 873.530 400.000 873.810 400.110 ;
        RECT 870.420 375.710 870.680 376.030 ;
        RECT 872.260 375.710 872.520 376.030 ;
        RECT 870.480 79.890 870.620 375.710 ;
        RECT 870.420 79.570 870.680 79.890 ;
        RECT 2195.680 79.570 2195.940 79.890 ;
        RECT 2195.740 2.400 2195.880 79.570 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 877.750 79.460 878.070 79.520 ;
        RECT 2213.130 79.460 2213.450 79.520 ;
        RECT 877.750 79.320 2213.450 79.460 ;
        RECT 877.750 79.260 878.070 79.320 ;
        RECT 2213.130 79.260 2213.450 79.320 ;
      LAYER via ;
        RECT 877.780 79.260 878.040 79.520 ;
        RECT 2213.160 79.260 2213.420 79.520 ;
      LAYER met2 ;
        RECT 879.050 400.250 879.330 404.000 ;
        RECT 877.840 400.110 879.330 400.250 ;
        RECT 877.840 79.550 877.980 400.110 ;
        RECT 879.050 400.000 879.330 400.110 ;
        RECT 877.780 79.230 878.040 79.550 ;
        RECT 2213.160 79.230 2213.420 79.550 ;
        RECT 2213.220 2.400 2213.360 79.230 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.690 45.460 436.010 45.520 ;
        RECT 777.010 45.460 777.330 45.520 ;
        RECT 435.690 45.320 777.330 45.460 ;
        RECT 435.690 45.260 436.010 45.320 ;
        RECT 777.010 45.260 777.330 45.320 ;
      LAYER via ;
        RECT 435.720 45.260 435.980 45.520 ;
        RECT 777.040 45.260 777.300 45.520 ;
      LAYER met2 ;
        RECT 437.910 400.250 438.190 404.000 ;
        RECT 436.700 400.110 438.190 400.250 ;
        RECT 436.700 324.370 436.840 400.110 ;
        RECT 437.910 400.000 438.190 400.110 ;
        RECT 435.780 324.230 436.840 324.370 ;
        RECT 435.780 45.550 435.920 324.230 ;
        RECT 435.720 45.230 435.980 45.550 ;
        RECT 777.040 45.230 777.300 45.550 ;
        RECT 777.100 2.400 777.240 45.230 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.570 400.250 884.850 404.000 ;
        RECT 884.280 400.110 884.850 400.250 ;
        RECT 884.280 80.085 884.420 400.110 ;
        RECT 884.570 400.000 884.850 400.110 ;
        RECT 884.210 79.715 884.490 80.085 ;
        RECT 2228.790 79.715 2229.070 80.085 ;
        RECT 2228.860 1.770 2229.000 79.715 ;
        RECT 2230.950 1.770 2231.510 2.400 ;
        RECT 2228.860 1.630 2231.510 1.770 ;
        RECT 2230.950 -4.800 2231.510 1.630 ;
      LAYER via2 ;
        RECT 884.210 79.760 884.490 80.040 ;
        RECT 2228.790 79.760 2229.070 80.040 ;
      LAYER met3 ;
        RECT 884.185 80.050 884.515 80.065 ;
        RECT 2228.765 80.050 2229.095 80.065 ;
        RECT 884.185 79.750 2229.095 80.050 ;
        RECT 884.185 79.735 884.515 79.750 ;
        RECT 2228.765 79.735 2229.095 79.750 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.630 398.720 890.950 398.780 ;
        RECT 891.550 398.720 891.870 398.780 ;
        RECT 890.630 398.580 891.870 398.720 ;
        RECT 890.630 398.520 890.950 398.580 ;
        RECT 891.550 398.520 891.870 398.580 ;
        RECT 2242.570 16.900 2242.890 16.960 ;
        RECT 2249.010 16.900 2249.330 16.960 ;
        RECT 2242.570 16.760 2249.330 16.900 ;
        RECT 2242.570 16.700 2242.890 16.760 ;
        RECT 2249.010 16.700 2249.330 16.760 ;
      LAYER via ;
        RECT 890.660 398.520 890.920 398.780 ;
        RECT 891.580 398.520 891.840 398.780 ;
        RECT 2242.600 16.700 2242.860 16.960 ;
        RECT 2249.040 16.700 2249.300 16.960 ;
      LAYER met2 ;
        RECT 890.090 400.250 890.370 404.000 ;
        RECT 890.090 400.110 890.860 400.250 ;
        RECT 890.090 400.000 890.370 400.110 ;
        RECT 890.720 398.810 890.860 400.110 ;
        RECT 890.660 398.490 890.920 398.810 ;
        RECT 891.580 398.490 891.840 398.810 ;
        RECT 891.640 351.970 891.780 398.490 ;
        RECT 891.180 351.830 891.780 351.970 ;
        RECT 891.180 79.405 891.320 351.830 ;
        RECT 891.110 79.035 891.390 79.405 ;
        RECT 2242.590 79.035 2242.870 79.405 ;
        RECT 2242.660 16.990 2242.800 79.035 ;
        RECT 2242.600 16.670 2242.860 16.990 ;
        RECT 2249.040 16.670 2249.300 16.990 ;
        RECT 2249.100 2.400 2249.240 16.670 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
      LAYER via2 ;
        RECT 891.110 79.080 891.390 79.360 ;
        RECT 2242.590 79.080 2242.870 79.360 ;
      LAYER met3 ;
        RECT 891.085 79.370 891.415 79.385 ;
        RECT 2242.565 79.370 2242.895 79.385 ;
        RECT 891.085 79.070 2242.895 79.370 ;
        RECT 891.085 79.055 891.415 79.070 ;
        RECT 2242.565 79.055 2242.895 79.070 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 891.550 122.980 891.870 123.040 ;
        RECT 2263.270 122.980 2263.590 123.040 ;
        RECT 891.550 122.840 2263.590 122.980 ;
        RECT 891.550 122.780 891.870 122.840 ;
        RECT 2263.270 122.780 2263.590 122.840 ;
      LAYER via ;
        RECT 891.580 122.780 891.840 123.040 ;
        RECT 2263.300 122.780 2263.560 123.040 ;
      LAYER met2 ;
        RECT 895.610 400.250 895.890 404.000 ;
        RECT 894.400 400.110 895.890 400.250 ;
        RECT 894.400 324.370 894.540 400.110 ;
        RECT 895.610 400.000 895.890 400.110 ;
        RECT 891.640 324.230 894.540 324.370 ;
        RECT 891.640 123.070 891.780 324.230 ;
        RECT 891.580 122.750 891.840 123.070 ;
        RECT 2263.300 122.750 2263.560 123.070 ;
        RECT 2263.360 82.870 2263.500 122.750 ;
        RECT 2263.360 82.730 2266.720 82.870 ;
        RECT 2266.580 2.400 2266.720 82.730 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 898.450 122.640 898.770 122.700 ;
        RECT 2284.430 122.640 2284.750 122.700 ;
        RECT 898.450 122.500 2284.750 122.640 ;
        RECT 898.450 122.440 898.770 122.500 ;
        RECT 2284.430 122.440 2284.750 122.500 ;
      LAYER via ;
        RECT 898.480 122.440 898.740 122.700 ;
        RECT 2284.460 122.440 2284.720 122.700 ;
      LAYER met2 ;
        RECT 900.670 400.250 900.950 404.000 ;
        RECT 899.920 400.110 900.950 400.250 ;
        RECT 899.920 324.370 900.060 400.110 ;
        RECT 900.670 400.000 900.950 400.110 ;
        RECT 898.540 324.230 900.060 324.370 ;
        RECT 898.540 122.730 898.680 324.230 ;
        RECT 898.480 122.410 898.740 122.730 ;
        RECT 2284.460 122.410 2284.720 122.730 ;
        RECT 2284.520 2.400 2284.660 122.410 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 905.350 122.300 905.670 122.360 ;
        RECT 2297.770 122.300 2298.090 122.360 ;
        RECT 905.350 122.160 2298.090 122.300 ;
        RECT 905.350 122.100 905.670 122.160 ;
        RECT 2297.770 122.100 2298.090 122.160 ;
      LAYER via ;
        RECT 905.380 122.100 905.640 122.360 ;
        RECT 2297.800 122.100 2298.060 122.360 ;
      LAYER met2 ;
        RECT 906.190 400.250 906.470 404.000 ;
        RECT 905.440 400.110 906.470 400.250 ;
        RECT 905.440 122.390 905.580 400.110 ;
        RECT 906.190 400.000 906.470 400.110 ;
        RECT 905.380 122.070 905.640 122.390 ;
        RECT 2297.800 122.070 2298.060 122.390 ;
        RECT 2297.860 82.870 2298.000 122.070 ;
        RECT 2297.860 82.730 2299.840 82.870 ;
        RECT 2299.700 1.770 2299.840 82.730 ;
        RECT 2301.790 1.770 2302.350 2.400 ;
        RECT 2299.700 1.630 2302.350 1.770 ;
        RECT 2301.790 -4.800 2302.350 1.630 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 911.790 121.960 912.110 122.020 ;
        RECT 2318.470 121.960 2318.790 122.020 ;
        RECT 911.790 121.820 2318.790 121.960 ;
        RECT 911.790 121.760 912.110 121.820 ;
        RECT 2318.470 121.760 2318.790 121.820 ;
      LAYER via ;
        RECT 911.820 121.760 912.080 122.020 ;
        RECT 2318.500 121.760 2318.760 122.020 ;
      LAYER met2 ;
        RECT 911.710 400.180 911.990 404.000 ;
        RECT 911.710 400.000 912.020 400.180 ;
        RECT 911.880 122.050 912.020 400.000 ;
        RECT 911.820 121.730 912.080 122.050 ;
        RECT 2318.500 121.730 2318.760 122.050 ;
        RECT 2318.560 82.870 2318.700 121.730 ;
        RECT 2318.560 82.730 2320.080 82.870 ;
        RECT 2319.940 2.400 2320.080 82.730 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 912.250 121.620 912.570 121.680 ;
        RECT 2332.270 121.620 2332.590 121.680 ;
        RECT 912.250 121.480 2332.590 121.620 ;
        RECT 912.250 121.420 912.570 121.480 ;
        RECT 2332.270 121.420 2332.590 121.480 ;
      LAYER via ;
        RECT 912.280 121.420 912.540 121.680 ;
        RECT 2332.300 121.420 2332.560 121.680 ;
      LAYER met2 ;
        RECT 917.230 400.250 917.510 404.000 ;
        RECT 916.020 400.110 917.510 400.250 ;
        RECT 916.020 324.370 916.160 400.110 ;
        RECT 917.230 400.000 917.510 400.110 ;
        RECT 912.340 324.230 916.160 324.370 ;
        RECT 912.340 121.710 912.480 324.230 ;
        RECT 912.280 121.390 912.540 121.710 ;
        RECT 2332.300 121.390 2332.560 121.710 ;
        RECT 2332.360 82.870 2332.500 121.390 ;
        RECT 2332.360 82.730 2337.560 82.870 ;
        RECT 2337.420 2.400 2337.560 82.730 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 918.690 84.900 919.010 84.960 ;
        RECT 2352.970 84.900 2353.290 84.960 ;
        RECT 918.690 84.760 2353.290 84.900 ;
        RECT 918.690 84.700 919.010 84.760 ;
        RECT 2352.970 84.700 2353.290 84.760 ;
      LAYER via ;
        RECT 918.720 84.700 918.980 84.960 ;
        RECT 2353.000 84.700 2353.260 84.960 ;
      LAYER met2 ;
        RECT 922.750 400.250 923.030 404.000 ;
        RECT 921.540 400.110 923.030 400.250 ;
        RECT 921.540 324.370 921.680 400.110 ;
        RECT 922.750 400.000 923.030 400.110 ;
        RECT 918.780 324.230 921.680 324.370 ;
        RECT 918.780 84.990 918.920 324.230 ;
        RECT 918.720 84.670 918.980 84.990 ;
        RECT 2353.000 84.670 2353.260 84.990 ;
        RECT 2353.060 1.770 2353.200 84.670 ;
        RECT 2355.150 1.770 2355.710 2.400 ;
        RECT 2353.060 1.630 2355.710 1.770 ;
        RECT 2355.150 -4.800 2355.710 1.630 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 926.050 85.240 926.370 85.300 ;
        RECT 2366.770 85.240 2367.090 85.300 ;
        RECT 926.050 85.100 2367.090 85.240 ;
        RECT 926.050 85.040 926.370 85.100 ;
        RECT 2366.770 85.040 2367.090 85.100 ;
        RECT 2366.770 17.580 2367.090 17.640 ;
        RECT 2370.910 17.580 2371.230 17.640 ;
        RECT 2366.770 17.440 2371.230 17.580 ;
        RECT 2366.770 17.380 2367.090 17.440 ;
        RECT 2370.910 17.380 2371.230 17.440 ;
      LAYER via ;
        RECT 926.080 85.040 926.340 85.300 ;
        RECT 2366.800 85.040 2367.060 85.300 ;
        RECT 2366.800 17.380 2367.060 17.640 ;
        RECT 2370.940 17.380 2371.200 17.640 ;
      LAYER met2 ;
        RECT 928.270 400.250 928.550 404.000 ;
        RECT 927.060 400.110 928.550 400.250 ;
        RECT 927.060 324.370 927.200 400.110 ;
        RECT 928.270 400.000 928.550 400.110 ;
        RECT 926.140 324.230 927.200 324.370 ;
        RECT 926.140 85.330 926.280 324.230 ;
        RECT 926.080 85.010 926.340 85.330 ;
        RECT 2366.800 85.010 2367.060 85.330 ;
        RECT 2366.860 17.670 2367.000 85.010 ;
        RECT 2366.800 17.350 2367.060 17.670 ;
        RECT 2370.940 17.350 2371.200 17.670 ;
        RECT 2371.000 1.770 2371.140 17.350 ;
        RECT 2372.630 1.770 2373.190 2.400 ;
        RECT 2371.000 1.630 2373.190 1.770 ;
        RECT 2372.630 -4.800 2373.190 1.630 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 932.490 85.580 932.810 85.640 ;
        RECT 2387.470 85.580 2387.790 85.640 ;
        RECT 932.490 85.440 2387.790 85.580 ;
        RECT 932.490 85.380 932.810 85.440 ;
        RECT 2387.470 85.380 2387.790 85.440 ;
      LAYER via ;
        RECT 932.520 85.380 932.780 85.640 ;
        RECT 2387.500 85.380 2387.760 85.640 ;
      LAYER met2 ;
        RECT 933.790 400.250 934.070 404.000 ;
        RECT 932.580 400.110 934.070 400.250 ;
        RECT 932.580 85.670 932.720 400.110 ;
        RECT 933.790 400.000 934.070 400.110 ;
        RECT 932.520 85.350 932.780 85.670 ;
        RECT 2387.500 85.350 2387.760 85.670 ;
        RECT 2387.560 82.870 2387.700 85.350 ;
        RECT 2387.560 82.730 2390.920 82.870 ;
        RECT 2390.780 2.400 2390.920 82.730 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 443.050 45.120 443.370 45.180 ;
        RECT 794.490 45.120 794.810 45.180 ;
        RECT 443.050 44.980 794.810 45.120 ;
        RECT 443.050 44.920 443.370 44.980 ;
        RECT 794.490 44.920 794.810 44.980 ;
      LAYER via ;
        RECT 443.080 44.920 443.340 45.180 ;
        RECT 794.520 44.920 794.780 45.180 ;
      LAYER met2 ;
        RECT 443.430 400.250 443.710 404.000 ;
        RECT 443.140 400.110 443.710 400.250 ;
        RECT 443.140 45.210 443.280 400.110 ;
        RECT 443.430 400.000 443.710 400.110 ;
        RECT 443.080 44.890 443.340 45.210 ;
        RECT 794.520 44.890 794.780 45.210 ;
        RECT 794.580 2.400 794.720 44.890 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 394.750 39.680 395.070 39.740 ;
        RECT 640.850 39.680 641.170 39.740 ;
        RECT 394.750 39.540 641.170 39.680 ;
        RECT 394.750 39.480 395.070 39.540 ;
        RECT 640.850 39.480 641.170 39.540 ;
      LAYER via ;
        RECT 394.780 39.480 395.040 39.740 ;
        RECT 640.880 39.480 641.140 39.740 ;
      LAYER met2 ;
        RECT 396.510 400.250 396.790 404.000 ;
        RECT 395.300 400.110 396.790 400.250 ;
        RECT 395.300 324.370 395.440 400.110 ;
        RECT 396.510 400.000 396.790 400.110 ;
        RECT 394.840 324.230 395.440 324.370 ;
        RECT 394.840 39.770 394.980 324.230 ;
        RECT 394.780 39.450 395.040 39.770 ;
        RECT 640.880 39.450 641.140 39.770 ;
        RECT 640.940 2.400 641.080 39.450 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 939.390 85.920 939.710 85.980 ;
        RECT 2408.170 85.920 2408.490 85.980 ;
        RECT 939.390 85.780 2408.490 85.920 ;
        RECT 939.390 85.720 939.710 85.780 ;
        RECT 2408.170 85.720 2408.490 85.780 ;
        RECT 2408.170 17.580 2408.490 17.640 ;
        RECT 2412.310 17.580 2412.630 17.640 ;
        RECT 2408.170 17.440 2412.630 17.580 ;
        RECT 2408.170 17.380 2408.490 17.440 ;
        RECT 2412.310 17.380 2412.630 17.440 ;
      LAYER via ;
        RECT 939.420 85.720 939.680 85.980 ;
        RECT 2408.200 85.720 2408.460 85.980 ;
        RECT 2408.200 17.380 2408.460 17.640 ;
        RECT 2412.340 17.380 2412.600 17.640 ;
      LAYER met2 ;
        RECT 940.690 400.250 940.970 404.000 ;
        RECT 939.480 400.110 940.970 400.250 ;
        RECT 939.480 86.010 939.620 400.110 ;
        RECT 940.690 400.000 940.970 400.110 ;
        RECT 939.420 85.690 939.680 86.010 ;
        RECT 2408.200 85.690 2408.460 86.010 ;
        RECT 2408.260 17.670 2408.400 85.690 ;
        RECT 2408.200 17.350 2408.460 17.670 ;
        RECT 2412.340 17.350 2412.600 17.670 ;
        RECT 2412.400 1.770 2412.540 17.350 ;
        RECT 2414.030 1.770 2414.590 2.400 ;
        RECT 2412.400 1.630 2414.590 1.770 ;
        RECT 2414.030 -4.800 2414.590 1.630 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 946.290 89.660 946.610 89.720 ;
        RECT 2428.870 89.660 2429.190 89.720 ;
        RECT 946.290 89.520 2429.190 89.660 ;
        RECT 946.290 89.460 946.610 89.520 ;
        RECT 2428.870 89.460 2429.190 89.520 ;
      LAYER via ;
        RECT 946.320 89.460 946.580 89.720 ;
        RECT 2428.900 89.460 2429.160 89.720 ;
      LAYER met2 ;
        RECT 946.210 400.180 946.490 404.000 ;
        RECT 946.210 400.000 946.520 400.180 ;
        RECT 946.380 89.750 946.520 400.000 ;
        RECT 946.320 89.430 946.580 89.750 ;
        RECT 2428.900 89.430 2429.160 89.750 ;
        RECT 2428.960 82.870 2429.100 89.430 ;
        RECT 2428.960 82.730 2432.320 82.870 ;
        RECT 2432.180 2.400 2432.320 82.730 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 945.830 386.140 946.150 386.200 ;
        RECT 950.430 386.140 950.750 386.200 ;
        RECT 945.830 386.000 950.750 386.140 ;
        RECT 945.830 385.940 946.150 386.000 ;
        RECT 950.430 385.940 950.750 386.000 ;
        RECT 945.830 89.320 946.150 89.380 ;
        RECT 2450.030 89.320 2450.350 89.380 ;
        RECT 945.830 89.180 2450.350 89.320 ;
        RECT 945.830 89.120 946.150 89.180 ;
        RECT 2450.030 89.120 2450.350 89.180 ;
      LAYER via ;
        RECT 945.860 385.940 946.120 386.200 ;
        RECT 950.460 385.940 950.720 386.200 ;
        RECT 945.860 89.120 946.120 89.380 ;
        RECT 2450.060 89.120 2450.320 89.380 ;
      LAYER met2 ;
        RECT 951.730 400.250 952.010 404.000 ;
        RECT 950.520 400.110 952.010 400.250 ;
        RECT 950.520 386.230 950.660 400.110 ;
        RECT 951.730 400.000 952.010 400.110 ;
        RECT 945.860 385.910 946.120 386.230 ;
        RECT 950.460 385.910 950.720 386.230 ;
        RECT 945.920 89.410 946.060 385.910 ;
        RECT 945.860 89.090 946.120 89.410 ;
        RECT 2450.060 89.090 2450.320 89.410 ;
        RECT 2450.120 16.730 2450.260 89.090 ;
        RECT 2449.660 16.590 2450.260 16.730 ;
        RECT 2449.660 2.400 2449.800 16.590 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 952.730 385.800 953.050 385.860 ;
        RECT 955.950 385.800 956.270 385.860 ;
        RECT 952.730 385.660 956.270 385.800 ;
        RECT 952.730 385.600 953.050 385.660 ;
        RECT 955.950 385.600 956.270 385.660 ;
        RECT 952.730 88.980 953.050 89.040 ;
        RECT 2463.370 88.980 2463.690 89.040 ;
        RECT 952.730 88.840 2463.690 88.980 ;
        RECT 952.730 88.780 953.050 88.840 ;
        RECT 2463.370 88.780 2463.690 88.840 ;
      LAYER via ;
        RECT 952.760 385.600 953.020 385.860 ;
        RECT 955.980 385.600 956.240 385.860 ;
        RECT 952.760 88.780 953.020 89.040 ;
        RECT 2463.400 88.780 2463.660 89.040 ;
      LAYER met2 ;
        RECT 957.250 400.250 957.530 404.000 ;
        RECT 956.040 400.110 957.530 400.250 ;
        RECT 956.040 385.890 956.180 400.110 ;
        RECT 957.250 400.000 957.530 400.110 ;
        RECT 952.760 385.570 953.020 385.890 ;
        RECT 955.980 385.570 956.240 385.890 ;
        RECT 952.820 89.070 952.960 385.570 ;
        RECT 952.760 88.750 953.020 89.070 ;
        RECT 2463.400 88.750 2463.660 89.070 ;
        RECT 2463.460 82.870 2463.600 88.750 ;
        RECT 2463.460 82.730 2465.440 82.870 ;
        RECT 2465.300 1.770 2465.440 82.730 ;
        RECT 2467.390 1.770 2467.950 2.400 ;
        RECT 2465.300 1.630 2467.950 1.770 ;
        RECT 2467.390 -4.800 2467.950 1.630 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 960.550 88.640 960.870 88.700 ;
        RECT 2484.070 88.640 2484.390 88.700 ;
        RECT 960.550 88.500 2484.390 88.640 ;
        RECT 960.550 88.440 960.870 88.500 ;
        RECT 2484.070 88.440 2484.390 88.500 ;
      LAYER via ;
        RECT 960.580 88.440 960.840 88.700 ;
        RECT 2484.100 88.440 2484.360 88.700 ;
      LAYER met2 ;
        RECT 962.770 400.250 963.050 404.000 ;
        RECT 961.560 400.110 963.050 400.250 ;
        RECT 961.560 324.370 961.700 400.110 ;
        RECT 962.770 400.000 963.050 400.110 ;
        RECT 960.640 324.230 961.700 324.370 ;
        RECT 960.640 88.730 960.780 324.230 ;
        RECT 960.580 88.410 960.840 88.730 ;
        RECT 2484.100 88.410 2484.360 88.730 ;
        RECT 2484.160 82.870 2484.300 88.410 ;
        RECT 2484.160 82.730 2485.680 82.870 ;
        RECT 2485.540 2.400 2485.680 82.730 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 966.990 88.300 967.310 88.360 ;
        RECT 2497.870 88.300 2498.190 88.360 ;
        RECT 966.990 88.160 2498.190 88.300 ;
        RECT 966.990 88.100 967.310 88.160 ;
        RECT 2497.870 88.100 2498.190 88.160 ;
      LAYER via ;
        RECT 967.020 88.100 967.280 88.360 ;
        RECT 2497.900 88.100 2498.160 88.360 ;
      LAYER met2 ;
        RECT 967.830 400.250 968.110 404.000 ;
        RECT 967.080 400.110 968.110 400.250 ;
        RECT 967.080 88.390 967.220 400.110 ;
        RECT 967.830 400.000 968.110 400.110 ;
        RECT 967.020 88.070 967.280 88.390 ;
        RECT 2497.900 88.070 2498.160 88.390 ;
        RECT 2497.960 82.870 2498.100 88.070 ;
        RECT 2497.960 82.730 2503.160 82.870 ;
        RECT 2503.020 2.400 2503.160 82.730 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.430 387.640 973.750 387.900 ;
        RECT 973.520 386.880 973.660 387.640 ;
        RECT 973.430 386.620 973.750 386.880 ;
        RECT 973.430 87.960 973.750 88.020 ;
        RECT 2518.570 87.960 2518.890 88.020 ;
        RECT 973.430 87.820 2518.890 87.960 ;
        RECT 973.430 87.760 973.750 87.820 ;
        RECT 2518.570 87.760 2518.890 87.820 ;
      LAYER via ;
        RECT 973.460 387.640 973.720 387.900 ;
        RECT 973.460 386.620 973.720 386.880 ;
        RECT 973.460 87.760 973.720 88.020 ;
        RECT 2518.600 87.760 2518.860 88.020 ;
      LAYER met2 ;
        RECT 973.350 400.180 973.630 404.000 ;
        RECT 973.350 400.000 973.660 400.180 ;
        RECT 973.520 387.930 973.660 400.000 ;
        RECT 973.460 387.610 973.720 387.930 ;
        RECT 973.460 386.590 973.720 386.910 ;
        RECT 973.520 88.050 973.660 386.590 ;
        RECT 973.460 87.730 973.720 88.050 ;
        RECT 2518.600 87.730 2518.860 88.050 ;
        RECT 2518.660 1.770 2518.800 87.730 ;
        RECT 2520.750 1.770 2521.310 2.400 ;
        RECT 2518.660 1.630 2521.310 1.770 ;
        RECT 2520.750 -4.800 2521.310 1.630 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.890 386.480 974.210 386.540 ;
        RECT 977.570 386.480 977.890 386.540 ;
        RECT 973.890 386.340 977.890 386.480 ;
        RECT 973.890 386.280 974.210 386.340 ;
        RECT 977.570 386.280 977.890 386.340 ;
        RECT 973.890 87.620 974.210 87.680 ;
        RECT 2532.830 87.620 2533.150 87.680 ;
        RECT 973.890 87.480 2533.150 87.620 ;
        RECT 973.890 87.420 974.210 87.480 ;
        RECT 2532.830 87.420 2533.150 87.480 ;
      LAYER via ;
        RECT 973.920 386.280 974.180 386.540 ;
        RECT 977.600 386.280 977.860 386.540 ;
        RECT 973.920 87.420 974.180 87.680 ;
        RECT 2532.860 87.420 2533.120 87.680 ;
      LAYER met2 ;
        RECT 978.870 400.250 979.150 404.000 ;
        RECT 977.660 400.110 979.150 400.250 ;
        RECT 977.660 386.570 977.800 400.110 ;
        RECT 978.870 400.000 979.150 400.110 ;
        RECT 973.920 386.250 974.180 386.570 ;
        RECT 977.600 386.250 977.860 386.570 ;
        RECT 973.980 87.710 974.120 386.250 ;
        RECT 973.920 87.390 974.180 87.710 ;
        RECT 2532.860 87.390 2533.120 87.710 ;
        RECT 2532.920 82.870 2533.060 87.390 ;
        RECT 2532.920 82.730 2536.280 82.870 ;
        RECT 2536.140 1.770 2536.280 82.730 ;
        RECT 2538.230 1.770 2538.790 2.400 ;
        RECT 2536.140 1.630 2538.790 1.770 ;
        RECT 2538.230 -4.800 2538.790 1.630 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 980.790 386.480 981.110 386.540 ;
        RECT 983.090 386.480 983.410 386.540 ;
        RECT 980.790 386.340 983.410 386.480 ;
        RECT 980.790 386.280 981.110 386.340 ;
        RECT 983.090 386.280 983.410 386.340 ;
        RECT 980.790 87.280 981.110 87.340 ;
        RECT 2553.070 87.280 2553.390 87.340 ;
        RECT 980.790 87.140 2553.390 87.280 ;
        RECT 980.790 87.080 981.110 87.140 ;
        RECT 2553.070 87.080 2553.390 87.140 ;
      LAYER via ;
        RECT 980.820 386.280 981.080 386.540 ;
        RECT 983.120 386.280 983.380 386.540 ;
        RECT 980.820 87.080 981.080 87.340 ;
        RECT 2553.100 87.080 2553.360 87.340 ;
      LAYER met2 ;
        RECT 984.390 400.250 984.670 404.000 ;
        RECT 983.180 400.110 984.670 400.250 ;
        RECT 983.180 386.570 983.320 400.110 ;
        RECT 984.390 400.000 984.670 400.110 ;
        RECT 980.820 386.250 981.080 386.570 ;
        RECT 983.120 386.250 983.380 386.570 ;
        RECT 980.880 87.370 981.020 386.250 ;
        RECT 980.820 87.050 981.080 87.370 ;
        RECT 2553.100 87.050 2553.360 87.370 ;
        RECT 2553.160 82.870 2553.300 87.050 ;
        RECT 2553.160 82.730 2556.520 82.870 ;
        RECT 2556.380 2.400 2556.520 82.730 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 987.230 386.480 987.550 386.540 ;
        RECT 988.610 386.480 988.930 386.540 ;
        RECT 987.230 386.340 988.930 386.480 ;
        RECT 987.230 386.280 987.550 386.340 ;
        RECT 988.610 386.280 988.930 386.340 ;
        RECT 987.230 86.940 987.550 87.000 ;
        RECT 2573.770 86.940 2574.090 87.000 ;
        RECT 987.230 86.800 2574.090 86.940 ;
        RECT 987.230 86.740 987.550 86.800 ;
        RECT 2573.770 86.740 2574.090 86.800 ;
      LAYER via ;
        RECT 987.260 386.280 987.520 386.540 ;
        RECT 988.640 386.280 988.900 386.540 ;
        RECT 987.260 86.740 987.520 87.000 ;
        RECT 2573.800 86.740 2574.060 87.000 ;
      LAYER met2 ;
        RECT 989.910 400.250 990.190 404.000 ;
        RECT 988.700 400.110 990.190 400.250 ;
        RECT 988.700 386.570 988.840 400.110 ;
        RECT 989.910 400.000 990.190 400.110 ;
        RECT 987.260 386.250 987.520 386.570 ;
        RECT 988.640 386.250 988.900 386.570 ;
        RECT 987.320 87.030 987.460 386.250 ;
        RECT 987.260 86.710 987.520 87.030 ;
        RECT 2573.800 86.710 2574.060 87.030 ;
        RECT 2573.860 2.400 2574.000 86.710 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 449.490 44.780 449.810 44.840 ;
        RECT 818.410 44.780 818.730 44.840 ;
        RECT 449.490 44.640 818.730 44.780 ;
        RECT 449.490 44.580 449.810 44.640 ;
        RECT 818.410 44.580 818.730 44.640 ;
      LAYER via ;
        RECT 449.520 44.580 449.780 44.840 ;
        RECT 818.440 44.580 818.700 44.840 ;
      LAYER met2 ;
        RECT 450.790 400.250 451.070 404.000 ;
        RECT 449.580 400.110 451.070 400.250 ;
        RECT 449.580 44.870 449.720 400.110 ;
        RECT 450.790 400.000 451.070 400.110 ;
        RECT 449.520 44.550 449.780 44.870 ;
        RECT 818.440 44.550 818.700 44.870 ;
        RECT 818.500 2.400 818.640 44.550 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 994.590 379.000 994.910 379.060 ;
        RECT 995.510 379.000 995.830 379.060 ;
        RECT 994.590 378.860 995.830 379.000 ;
        RECT 994.590 378.800 994.910 378.860 ;
        RECT 995.510 378.800 995.830 378.860 ;
        RECT 994.590 86.600 994.910 86.660 ;
        RECT 2587.570 86.600 2587.890 86.660 ;
        RECT 994.590 86.460 2587.890 86.600 ;
        RECT 994.590 86.400 994.910 86.460 ;
        RECT 2587.570 86.400 2587.890 86.460 ;
      LAYER via ;
        RECT 994.620 378.800 994.880 379.060 ;
        RECT 995.540 378.800 995.800 379.060 ;
        RECT 994.620 86.400 994.880 86.660 ;
        RECT 2587.600 86.400 2587.860 86.660 ;
      LAYER met2 ;
        RECT 995.430 400.180 995.710 404.000 ;
        RECT 995.430 400.000 995.740 400.180 ;
        RECT 995.600 379.090 995.740 400.000 ;
        RECT 994.620 378.770 994.880 379.090 ;
        RECT 995.540 378.770 995.800 379.090 ;
        RECT 994.680 86.690 994.820 378.770 ;
        RECT 994.620 86.370 994.880 86.690 ;
        RECT 2587.600 86.370 2587.860 86.690 ;
        RECT 2587.660 82.870 2587.800 86.370 ;
        RECT 2587.660 82.730 2589.640 82.870 ;
        RECT 2589.500 1.770 2589.640 82.730 ;
        RECT 2591.590 1.770 2592.150 2.400 ;
        RECT 2589.500 1.630 2592.150 1.770 ;
        RECT 2591.590 -4.800 2592.150 1.630 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1001.490 86.260 1001.810 86.320 ;
        RECT 2608.270 86.260 2608.590 86.320 ;
        RECT 1001.490 86.120 2608.590 86.260 ;
        RECT 1001.490 86.060 1001.810 86.120 ;
        RECT 2608.270 86.060 2608.590 86.120 ;
      LAYER via ;
        RECT 1001.520 86.060 1001.780 86.320 ;
        RECT 2608.300 86.060 2608.560 86.320 ;
      LAYER met2 ;
        RECT 1000.490 400.250 1000.770 404.000 ;
        RECT 1000.490 400.110 1001.720 400.250 ;
        RECT 1000.490 400.000 1000.770 400.110 ;
        RECT 1001.580 86.350 1001.720 400.110 ;
        RECT 1001.520 86.030 1001.780 86.350 ;
        RECT 2608.300 86.030 2608.560 86.350 ;
        RECT 2608.360 1.770 2608.500 86.030 ;
        RECT 2609.070 1.770 2609.630 2.400 ;
        RECT 2608.360 1.630 2609.630 1.770 ;
        RECT 2609.070 -4.800 2609.630 1.630 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.010 400.250 1006.290 404.000 ;
        RECT 1004.800 400.110 1006.290 400.250 ;
        RECT 1004.800 324.370 1004.940 400.110 ;
        RECT 1006.010 400.000 1006.290 400.110 ;
        RECT 1002.040 324.230 1004.940 324.370 ;
        RECT 1002.040 86.885 1002.180 324.230 ;
        RECT 1001.970 86.515 1002.250 86.885 ;
        RECT 2622.090 86.515 2622.370 86.885 ;
        RECT 2622.160 82.870 2622.300 86.515 ;
        RECT 2622.160 82.730 2627.360 82.870 ;
        RECT 2627.220 2.400 2627.360 82.730 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
      LAYER via2 ;
        RECT 1001.970 86.560 1002.250 86.840 ;
        RECT 2622.090 86.560 2622.370 86.840 ;
      LAYER met3 ;
        RECT 1001.945 86.850 1002.275 86.865 ;
        RECT 2622.065 86.850 2622.395 86.865 ;
        RECT 1001.945 86.550 2622.395 86.850 ;
        RECT 1001.945 86.535 1002.275 86.550 ;
        RECT 2622.065 86.535 2622.395 86.550 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.530 400.250 1011.810 404.000 ;
        RECT 1010.320 400.110 1011.810 400.250 ;
        RECT 1010.320 324.370 1010.460 400.110 ;
        RECT 1011.530 400.000 1011.810 400.110 ;
        RECT 1008.940 324.230 1010.460 324.370 ;
        RECT 1008.940 86.205 1009.080 324.230 ;
        RECT 1008.870 85.835 1009.150 86.205 ;
        RECT 2642.790 85.835 2643.070 86.205 ;
        RECT 2642.860 1.770 2643.000 85.835 ;
        RECT 2644.950 1.770 2645.510 2.400 ;
        RECT 2642.860 1.630 2645.510 1.770 ;
        RECT 2644.950 -4.800 2645.510 1.630 ;
      LAYER via2 ;
        RECT 1008.870 85.880 1009.150 86.160 ;
        RECT 2642.790 85.880 2643.070 86.160 ;
      LAYER met3 ;
        RECT 1008.845 86.170 1009.175 86.185 ;
        RECT 2642.765 86.170 2643.095 86.185 ;
        RECT 1008.845 85.870 2643.095 86.170 ;
        RECT 1008.845 85.855 1009.175 85.870 ;
        RECT 2642.765 85.855 2643.095 85.870 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1015.750 121.280 1016.070 121.340 ;
        RECT 2656.570 121.280 2656.890 121.340 ;
        RECT 1015.750 121.140 2656.890 121.280 ;
        RECT 1015.750 121.080 1016.070 121.140 ;
        RECT 2656.570 121.080 2656.890 121.140 ;
        RECT 2656.570 17.580 2656.890 17.640 ;
        RECT 2660.710 17.580 2661.030 17.640 ;
        RECT 2656.570 17.440 2661.030 17.580 ;
        RECT 2656.570 17.380 2656.890 17.440 ;
        RECT 2660.710 17.380 2661.030 17.440 ;
      LAYER via ;
        RECT 1015.780 121.080 1016.040 121.340 ;
        RECT 2656.600 121.080 2656.860 121.340 ;
        RECT 2656.600 17.380 2656.860 17.640 ;
        RECT 2660.740 17.380 2661.000 17.640 ;
      LAYER met2 ;
        RECT 1017.050 400.250 1017.330 404.000 ;
        RECT 1015.840 400.110 1017.330 400.250 ;
        RECT 1015.840 121.370 1015.980 400.110 ;
        RECT 1017.050 400.000 1017.330 400.110 ;
        RECT 1015.780 121.050 1016.040 121.370 ;
        RECT 2656.600 121.050 2656.860 121.370 ;
        RECT 2656.660 17.670 2656.800 121.050 ;
        RECT 2656.600 17.350 2656.860 17.670 ;
        RECT 2660.740 17.350 2661.000 17.670 ;
        RECT 2660.800 1.770 2660.940 17.350 ;
        RECT 2662.430 1.770 2662.990 2.400 ;
        RECT 2660.800 1.630 2662.990 1.770 ;
        RECT 2662.430 -4.800 2662.990 1.630 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.190 120.940 1022.510 121.000 ;
        RECT 2677.270 120.940 2677.590 121.000 ;
        RECT 1022.190 120.800 2677.590 120.940 ;
        RECT 1022.190 120.740 1022.510 120.800 ;
        RECT 2677.270 120.740 2677.590 120.800 ;
      LAYER via ;
        RECT 1022.220 120.740 1022.480 121.000 ;
        RECT 2677.300 120.740 2677.560 121.000 ;
      LAYER met2 ;
        RECT 1022.570 400.250 1022.850 404.000 ;
        RECT 1022.280 400.110 1022.850 400.250 ;
        RECT 1022.280 121.030 1022.420 400.110 ;
        RECT 1022.570 400.000 1022.850 400.110 ;
        RECT 1022.220 120.710 1022.480 121.030 ;
        RECT 2677.300 120.710 2677.560 121.030 ;
        RECT 2677.360 82.870 2677.500 120.710 ;
        RECT 2677.360 82.730 2680.720 82.870 ;
        RECT 2680.580 2.400 2680.720 82.730 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1027.710 386.480 1028.030 386.540 ;
        RECT 1029.550 386.480 1029.870 386.540 ;
        RECT 1027.710 386.340 1029.870 386.480 ;
        RECT 1027.710 386.280 1028.030 386.340 ;
        RECT 1029.550 386.280 1029.870 386.340 ;
        RECT 1029.550 120.600 1029.870 120.660 ;
        RECT 2697.970 120.600 2698.290 120.660 ;
        RECT 1029.550 120.460 2698.290 120.600 ;
        RECT 1029.550 120.400 1029.870 120.460 ;
        RECT 2697.970 120.400 2698.290 120.460 ;
      LAYER via ;
        RECT 1027.740 386.280 1028.000 386.540 ;
        RECT 1029.580 386.280 1029.840 386.540 ;
        RECT 1029.580 120.400 1029.840 120.660 ;
        RECT 2698.000 120.400 2698.260 120.660 ;
      LAYER met2 ;
        RECT 1028.090 400.180 1028.370 404.000 ;
        RECT 1028.090 400.000 1028.400 400.180 ;
        RECT 1028.260 389.370 1028.400 400.000 ;
        RECT 1028.030 389.230 1028.400 389.370 ;
        RECT 1028.030 388.690 1028.170 389.230 ;
        RECT 1027.800 388.550 1028.170 388.690 ;
        RECT 1027.800 386.570 1027.940 388.550 ;
        RECT 1027.740 386.250 1028.000 386.570 ;
        RECT 1029.580 386.250 1029.840 386.570 ;
        RECT 1029.640 120.690 1029.780 386.250 ;
        RECT 1029.580 120.370 1029.840 120.690 ;
        RECT 2698.000 120.370 2698.260 120.690 ;
        RECT 2698.060 2.400 2698.200 120.370 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1029.090 376.280 1029.410 376.340 ;
        RECT 1032.310 376.280 1032.630 376.340 ;
        RECT 1029.090 376.140 1032.630 376.280 ;
        RECT 1029.090 376.080 1029.410 376.140 ;
        RECT 1032.310 376.080 1032.630 376.140 ;
      LAYER via ;
        RECT 1029.120 376.080 1029.380 376.340 ;
        RECT 1032.340 376.080 1032.600 376.340 ;
      LAYER met2 ;
        RECT 1033.610 400.250 1033.890 404.000 ;
        RECT 1032.400 400.110 1033.890 400.250 ;
        RECT 1032.400 376.370 1032.540 400.110 ;
        RECT 1033.610 400.000 1033.890 400.110 ;
        RECT 1029.120 376.050 1029.380 376.370 ;
        RECT 1032.340 376.050 1032.600 376.370 ;
        RECT 1029.180 120.885 1029.320 376.050 ;
        RECT 1029.110 120.515 1029.390 120.885 ;
        RECT 2711.790 120.515 2712.070 120.885 ;
        RECT 2711.860 82.870 2712.000 120.515 ;
        RECT 2711.860 82.730 2713.840 82.870 ;
        RECT 2713.700 1.770 2713.840 82.730 ;
        RECT 2715.790 1.770 2716.350 2.400 ;
        RECT 2713.700 1.630 2716.350 1.770 ;
        RECT 2715.790 -4.800 2716.350 1.630 ;
      LAYER via2 ;
        RECT 1029.110 120.560 1029.390 120.840 ;
        RECT 2711.790 120.560 2712.070 120.840 ;
      LAYER met3 ;
        RECT 1029.085 120.850 1029.415 120.865 ;
        RECT 2711.765 120.850 2712.095 120.865 ;
        RECT 1029.085 120.550 2712.095 120.850 ;
        RECT 1029.085 120.535 1029.415 120.550 ;
        RECT 2711.765 120.535 2712.095 120.550 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1036.450 95.100 1036.770 95.160 ;
        RECT 2732.470 95.100 2732.790 95.160 ;
        RECT 1036.450 94.960 2732.790 95.100 ;
        RECT 1036.450 94.900 1036.770 94.960 ;
        RECT 2732.470 94.900 2732.790 94.960 ;
      LAYER via ;
        RECT 1036.480 94.900 1036.740 95.160 ;
        RECT 2732.500 94.900 2732.760 95.160 ;
      LAYER met2 ;
        RECT 1038.670 400.250 1038.950 404.000 ;
        RECT 1037.460 400.110 1038.950 400.250 ;
        RECT 1037.460 303.670 1037.600 400.110 ;
        RECT 1038.670 400.000 1038.950 400.110 ;
        RECT 1036.540 303.530 1037.600 303.670 ;
        RECT 1036.540 95.190 1036.680 303.530 ;
        RECT 1036.480 94.870 1036.740 95.190 ;
        RECT 2732.500 94.870 2732.760 95.190 ;
        RECT 2732.560 1.770 2732.700 94.870 ;
        RECT 2733.270 1.770 2733.830 2.400 ;
        RECT 2732.560 1.630 2733.830 1.770 ;
        RECT 2733.270 -4.800 2733.830 1.630 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1043.350 94.760 1043.670 94.820 ;
        RECT 2746.270 94.760 2746.590 94.820 ;
        RECT 1043.350 94.620 2746.590 94.760 ;
        RECT 1043.350 94.560 1043.670 94.620 ;
        RECT 2746.270 94.560 2746.590 94.620 ;
      LAYER via ;
        RECT 1043.380 94.560 1043.640 94.820 ;
        RECT 2746.300 94.560 2746.560 94.820 ;
      LAYER met2 ;
        RECT 1044.190 400.250 1044.470 404.000 ;
        RECT 1043.440 400.110 1044.470 400.250 ;
        RECT 1043.440 94.850 1043.580 400.110 ;
        RECT 1044.190 400.000 1044.470 400.110 ;
        RECT 1043.380 94.530 1043.640 94.850 ;
        RECT 2746.300 94.530 2746.560 94.850 ;
        RECT 2746.360 82.870 2746.500 94.530 ;
        RECT 2746.360 82.730 2751.560 82.870 ;
        RECT 2751.420 2.400 2751.560 82.730 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 455.930 40.020 456.250 40.080 ;
        RECT 669.370 40.020 669.690 40.080 ;
        RECT 455.930 39.880 669.690 40.020 ;
        RECT 455.930 39.820 456.250 39.880 ;
        RECT 669.370 39.820 669.690 39.880 ;
        RECT 669.370 16.900 669.690 16.960 ;
        RECT 835.890 16.900 836.210 16.960 ;
        RECT 669.370 16.760 836.210 16.900 ;
        RECT 669.370 16.700 669.690 16.760 ;
        RECT 835.890 16.700 836.210 16.760 ;
      LAYER via ;
        RECT 455.960 39.820 456.220 40.080 ;
        RECT 669.400 39.820 669.660 40.080 ;
        RECT 669.400 16.700 669.660 16.960 ;
        RECT 835.920 16.700 836.180 16.960 ;
      LAYER met2 ;
        RECT 456.310 400.250 456.590 404.000 ;
        RECT 456.020 400.110 456.590 400.250 ;
        RECT 456.020 40.110 456.160 400.110 ;
        RECT 456.310 400.000 456.590 400.110 ;
        RECT 455.960 39.790 456.220 40.110 ;
        RECT 669.400 39.790 669.660 40.110 ;
        RECT 669.460 16.990 669.600 39.790 ;
        RECT 669.400 16.670 669.660 16.990 ;
        RECT 835.920 16.670 836.180 16.990 ;
        RECT 835.980 2.400 836.120 16.670 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.790 94.420 1050.110 94.480 ;
        RECT 2766.970 94.420 2767.290 94.480 ;
        RECT 1049.790 94.280 2767.290 94.420 ;
        RECT 1049.790 94.220 1050.110 94.280 ;
        RECT 2766.970 94.220 2767.290 94.280 ;
      LAYER via ;
        RECT 1049.820 94.220 1050.080 94.480 ;
        RECT 2767.000 94.220 2767.260 94.480 ;
      LAYER met2 ;
        RECT 1049.710 400.180 1049.990 404.000 ;
        RECT 1049.710 400.000 1050.020 400.180 ;
        RECT 1049.880 94.510 1050.020 400.000 ;
        RECT 1049.820 94.190 1050.080 94.510 ;
        RECT 2767.000 94.190 2767.260 94.510 ;
        RECT 2767.060 82.870 2767.200 94.190 ;
        RECT 2767.060 82.730 2769.040 82.870 ;
        RECT 2768.900 2.400 2769.040 82.730 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.330 375.940 1049.650 376.000 ;
        RECT 1053.930 375.940 1054.250 376.000 ;
        RECT 1049.330 375.800 1054.250 375.940 ;
        RECT 1049.330 375.740 1049.650 375.800 ;
        RECT 1053.930 375.740 1054.250 375.800 ;
        RECT 1049.330 94.080 1049.650 94.140 ;
        RECT 2780.770 94.080 2781.090 94.140 ;
        RECT 1049.330 93.940 2781.090 94.080 ;
        RECT 1049.330 93.880 1049.650 93.940 ;
        RECT 2780.770 93.880 2781.090 93.940 ;
        RECT 2780.770 17.580 2781.090 17.640 ;
        RECT 2784.910 17.580 2785.230 17.640 ;
        RECT 2780.770 17.440 2785.230 17.580 ;
        RECT 2780.770 17.380 2781.090 17.440 ;
        RECT 2784.910 17.380 2785.230 17.440 ;
      LAYER via ;
        RECT 1049.360 375.740 1049.620 376.000 ;
        RECT 1053.960 375.740 1054.220 376.000 ;
        RECT 1049.360 93.880 1049.620 94.140 ;
        RECT 2780.800 93.880 2781.060 94.140 ;
        RECT 2780.800 17.380 2781.060 17.640 ;
        RECT 2784.940 17.380 2785.200 17.640 ;
      LAYER met2 ;
        RECT 1055.230 400.250 1055.510 404.000 ;
        RECT 1054.020 400.110 1055.510 400.250 ;
        RECT 1054.020 376.030 1054.160 400.110 ;
        RECT 1055.230 400.000 1055.510 400.110 ;
        RECT 1049.360 375.710 1049.620 376.030 ;
        RECT 1053.960 375.710 1054.220 376.030 ;
        RECT 1049.420 94.170 1049.560 375.710 ;
        RECT 1049.360 93.850 1049.620 94.170 ;
        RECT 2780.800 93.850 2781.060 94.170 ;
        RECT 2780.860 17.670 2781.000 93.850 ;
        RECT 2780.800 17.350 2781.060 17.670 ;
        RECT 2784.940 17.350 2785.200 17.670 ;
        RECT 2785.000 1.770 2785.140 17.350 ;
        RECT 2786.630 1.770 2787.190 2.400 ;
        RECT 2785.000 1.630 2787.190 1.770 ;
        RECT 2786.630 -4.800 2787.190 1.630 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1056.230 376.280 1056.550 376.340 ;
        RECT 1059.450 376.280 1059.770 376.340 ;
        RECT 1056.230 376.140 1059.770 376.280 ;
        RECT 1056.230 376.080 1056.550 376.140 ;
        RECT 1059.450 376.080 1059.770 376.140 ;
        RECT 1056.230 93.740 1056.550 93.800 ;
        RECT 2801.470 93.740 2801.790 93.800 ;
        RECT 1056.230 93.600 2801.790 93.740 ;
        RECT 1056.230 93.540 1056.550 93.600 ;
        RECT 2801.470 93.540 2801.790 93.600 ;
      LAYER via ;
        RECT 1056.260 376.080 1056.520 376.340 ;
        RECT 1059.480 376.080 1059.740 376.340 ;
        RECT 1056.260 93.540 1056.520 93.800 ;
        RECT 2801.500 93.540 2801.760 93.800 ;
      LAYER met2 ;
        RECT 1060.750 400.250 1061.030 404.000 ;
        RECT 1059.540 400.110 1061.030 400.250 ;
        RECT 1059.540 376.370 1059.680 400.110 ;
        RECT 1060.750 400.000 1061.030 400.110 ;
        RECT 1056.260 376.050 1056.520 376.370 ;
        RECT 1059.480 376.050 1059.740 376.370 ;
        RECT 1056.320 93.830 1056.460 376.050 ;
        RECT 1056.260 93.510 1056.520 93.830 ;
        RECT 2801.500 93.510 2801.760 93.830 ;
        RECT 2801.560 82.870 2801.700 93.510 ;
        RECT 2801.560 82.730 2802.160 82.870 ;
        RECT 2802.020 1.770 2802.160 82.730 ;
        RECT 2804.110 1.770 2804.670 2.400 ;
        RECT 2802.020 1.630 2804.670 1.770 ;
        RECT 2804.110 -4.800 2804.670 1.630 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1063.130 303.520 1063.450 303.580 ;
        RECT 1064.050 303.520 1064.370 303.580 ;
        RECT 1063.130 303.380 1064.370 303.520 ;
        RECT 1063.130 303.320 1063.450 303.380 ;
        RECT 1064.050 303.320 1064.370 303.380 ;
        RECT 1063.130 93.400 1063.450 93.460 ;
        RECT 2822.630 93.400 2822.950 93.460 ;
        RECT 1063.130 93.260 2822.950 93.400 ;
        RECT 1063.130 93.200 1063.450 93.260 ;
        RECT 2822.630 93.200 2822.950 93.260 ;
      LAYER via ;
        RECT 1063.160 303.320 1063.420 303.580 ;
        RECT 1064.080 303.320 1064.340 303.580 ;
        RECT 1063.160 93.200 1063.420 93.460 ;
        RECT 2822.660 93.200 2822.920 93.460 ;
      LAYER met2 ;
        RECT 1066.270 400.250 1066.550 404.000 ;
        RECT 1065.060 400.110 1066.550 400.250 ;
        RECT 1065.060 351.970 1065.200 400.110 ;
        RECT 1066.270 400.000 1066.550 400.110 ;
        RECT 1064.140 351.830 1065.200 351.970 ;
        RECT 1064.140 303.610 1064.280 351.830 ;
        RECT 1063.160 303.290 1063.420 303.610 ;
        RECT 1064.080 303.290 1064.340 303.610 ;
        RECT 1063.220 93.490 1063.360 303.290 ;
        RECT 1063.160 93.170 1063.420 93.490 ;
        RECT 2822.660 93.170 2822.920 93.490 ;
        RECT 2822.720 34.570 2822.860 93.170 ;
        RECT 2822.260 34.430 2822.860 34.570 ;
        RECT 2822.260 2.400 2822.400 34.430 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1070.490 93.060 1070.810 93.120 ;
        RECT 2835.970 93.060 2836.290 93.120 ;
        RECT 1070.490 92.920 2836.290 93.060 ;
        RECT 1070.490 92.860 1070.810 92.920 ;
        RECT 2835.970 92.860 2836.290 92.920 ;
      LAYER via ;
        RECT 1070.520 92.860 1070.780 93.120 ;
        RECT 2836.000 92.860 2836.260 93.120 ;
      LAYER met2 ;
        RECT 1071.330 400.250 1071.610 404.000 ;
        RECT 1070.580 400.110 1071.610 400.250 ;
        RECT 1070.580 93.150 1070.720 400.110 ;
        RECT 1071.330 400.000 1071.610 400.110 ;
        RECT 1070.520 92.830 1070.780 93.150 ;
        RECT 2836.000 92.830 2836.260 93.150 ;
        RECT 2836.060 82.870 2836.200 92.830 ;
        RECT 2836.060 82.730 2838.040 82.870 ;
        RECT 2837.900 1.770 2838.040 82.730 ;
        RECT 2839.990 1.770 2840.550 2.400 ;
        RECT 2837.900 1.630 2840.550 1.770 ;
        RECT 2839.990 -4.800 2840.550 1.630 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.850 400.250 1077.130 404.000 ;
        RECT 1076.850 400.110 1077.620 400.250 ;
        RECT 1076.850 400.000 1077.130 400.110 ;
        RECT 1077.480 93.685 1077.620 400.110 ;
        RECT 1077.410 93.315 1077.690 93.685 ;
        RECT 2856.690 93.315 2856.970 93.685 ;
        RECT 2856.760 1.770 2856.900 93.315 ;
        RECT 2857.470 1.770 2858.030 2.400 ;
        RECT 2856.760 1.630 2858.030 1.770 ;
        RECT 2857.470 -4.800 2858.030 1.630 ;
      LAYER via2 ;
        RECT 1077.410 93.360 1077.690 93.640 ;
        RECT 2856.690 93.360 2856.970 93.640 ;
      LAYER met3 ;
        RECT 1077.385 93.650 1077.715 93.665 ;
        RECT 2856.665 93.650 2856.995 93.665 ;
        RECT 1077.385 93.350 2856.995 93.650 ;
        RECT 1077.385 93.335 1077.715 93.350 ;
        RECT 2856.665 93.335 2856.995 93.350 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.370 400.250 1082.650 404.000 ;
        RECT 1081.160 400.110 1082.650 400.250 ;
        RECT 1081.160 324.370 1081.300 400.110 ;
        RECT 1082.370 400.000 1082.650 400.110 ;
        RECT 1078.400 324.230 1081.300 324.370 ;
        RECT 1078.400 93.005 1078.540 324.230 ;
        RECT 1078.330 92.635 1078.610 93.005 ;
        RECT 2870.490 92.635 2870.770 93.005 ;
        RECT 2870.560 82.870 2870.700 92.635 ;
        RECT 2870.560 82.730 2875.760 82.870 ;
        RECT 2875.620 2.400 2875.760 82.730 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
      LAYER via2 ;
        RECT 1078.330 92.680 1078.610 92.960 ;
        RECT 2870.490 92.680 2870.770 92.960 ;
      LAYER met3 ;
        RECT 1078.305 92.970 1078.635 92.985 ;
        RECT 2870.465 92.970 2870.795 92.985 ;
        RECT 1078.305 92.670 2870.795 92.970 ;
        RECT 1078.305 92.655 1078.635 92.670 ;
        RECT 2870.465 92.655 2870.795 92.670 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.750 58.720 1085.070 58.780 ;
        RECT 2893.010 58.720 2893.330 58.780 ;
        RECT 1084.750 58.580 2893.330 58.720 ;
        RECT 1084.750 58.520 1085.070 58.580 ;
        RECT 2893.010 58.520 2893.330 58.580 ;
      LAYER via ;
        RECT 1084.780 58.520 1085.040 58.780 ;
        RECT 2893.040 58.520 2893.300 58.780 ;
      LAYER met2 ;
        RECT 1087.890 400.250 1088.170 404.000 ;
        RECT 1086.680 400.110 1088.170 400.250 ;
        RECT 1086.680 324.370 1086.820 400.110 ;
        RECT 1087.890 400.000 1088.170 400.110 ;
        RECT 1084.840 324.230 1086.820 324.370 ;
        RECT 1084.840 58.810 1084.980 324.230 ;
        RECT 1084.780 58.490 1085.040 58.810 ;
        RECT 2893.040 58.490 2893.300 58.810 ;
        RECT 2893.100 2.400 2893.240 58.490 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 456.390 376.280 456.710 376.340 ;
        RECT 460.530 376.280 460.850 376.340 ;
        RECT 456.390 376.140 460.850 376.280 ;
        RECT 456.390 376.080 456.710 376.140 ;
        RECT 460.530 376.080 460.850 376.140 ;
        RECT 456.390 53.620 456.710 53.680 ;
        RECT 851.530 53.620 851.850 53.680 ;
        RECT 456.390 53.480 851.850 53.620 ;
        RECT 456.390 53.420 456.710 53.480 ;
        RECT 851.530 53.420 851.850 53.480 ;
      LAYER via ;
        RECT 456.420 376.080 456.680 376.340 ;
        RECT 460.560 376.080 460.820 376.340 ;
        RECT 456.420 53.420 456.680 53.680 ;
        RECT 851.560 53.420 851.820 53.680 ;
      LAYER met2 ;
        RECT 461.830 400.250 462.110 404.000 ;
        RECT 460.620 400.110 462.110 400.250 ;
        RECT 460.620 376.370 460.760 400.110 ;
        RECT 461.830 400.000 462.110 400.110 ;
        RECT 456.420 376.050 456.680 376.370 ;
        RECT 460.560 376.050 460.820 376.370 ;
        RECT 456.480 53.710 456.620 376.050 ;
        RECT 456.420 53.390 456.680 53.710 ;
        RECT 851.560 53.390 851.820 53.710 ;
        RECT 851.620 1.770 851.760 53.390 ;
        RECT 853.710 1.770 854.270 2.400 ;
        RECT 851.620 1.630 854.270 1.770 ;
        RECT 853.710 -4.800 854.270 1.630 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 463.290 53.280 463.610 53.340 ;
        RECT 870.390 53.280 870.710 53.340 ;
        RECT 463.290 53.140 870.710 53.280 ;
        RECT 463.290 53.080 463.610 53.140 ;
        RECT 870.390 53.080 870.710 53.140 ;
      LAYER via ;
        RECT 463.320 53.080 463.580 53.340 ;
        RECT 870.420 53.080 870.680 53.340 ;
      LAYER met2 ;
        RECT 466.890 400.250 467.170 404.000 ;
        RECT 466.140 400.110 467.170 400.250 ;
        RECT 466.140 351.970 466.280 400.110 ;
        RECT 466.890 400.000 467.170 400.110 ;
        RECT 463.380 351.830 466.280 351.970 ;
        RECT 463.380 53.370 463.520 351.830 ;
        RECT 463.320 53.050 463.580 53.370 ;
        RECT 870.420 53.050 870.680 53.370 ;
        RECT 870.480 1.770 870.620 53.050 ;
        RECT 871.190 1.770 871.750 2.400 ;
        RECT 870.480 1.630 871.750 1.770 ;
        RECT 871.190 -4.800 871.750 1.630 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 469.730 52.940 470.050 53.000 ;
        RECT 884.190 52.940 884.510 53.000 ;
        RECT 469.730 52.800 884.510 52.940 ;
        RECT 469.730 52.740 470.050 52.800 ;
        RECT 884.190 52.740 884.510 52.800 ;
        RECT 884.190 18.600 884.510 18.660 ;
        RECT 889.250 18.600 889.570 18.660 ;
        RECT 884.190 18.460 889.570 18.600 ;
        RECT 884.190 18.400 884.510 18.460 ;
        RECT 889.250 18.400 889.570 18.460 ;
      LAYER via ;
        RECT 469.760 52.740 470.020 53.000 ;
        RECT 884.220 52.740 884.480 53.000 ;
        RECT 884.220 18.400 884.480 18.660 ;
        RECT 889.280 18.400 889.540 18.660 ;
      LAYER met2 ;
        RECT 472.410 400.250 472.690 404.000 ;
        RECT 471.200 400.110 472.690 400.250 ;
        RECT 471.200 324.370 471.340 400.110 ;
        RECT 472.410 400.000 472.690 400.110 ;
        RECT 469.820 324.230 471.340 324.370 ;
        RECT 469.820 53.030 469.960 324.230 ;
        RECT 469.760 52.710 470.020 53.030 ;
        RECT 884.220 52.710 884.480 53.030 ;
        RECT 884.280 18.690 884.420 52.710 ;
        RECT 884.220 18.370 884.480 18.690 ;
        RECT 889.280 18.370 889.540 18.690 ;
        RECT 889.340 2.400 889.480 18.370 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 476.630 52.260 476.950 52.320 ;
        RECT 904.890 52.260 905.210 52.320 ;
        RECT 476.630 52.120 905.210 52.260 ;
        RECT 476.630 52.060 476.950 52.120 ;
        RECT 904.890 52.060 905.210 52.120 ;
      LAYER via ;
        RECT 476.660 52.060 476.920 52.320 ;
        RECT 904.920 52.060 905.180 52.320 ;
      LAYER met2 ;
        RECT 477.930 400.250 478.210 404.000 ;
        RECT 476.720 400.110 478.210 400.250 ;
        RECT 476.720 52.350 476.860 400.110 ;
        RECT 477.930 400.000 478.210 400.110 ;
        RECT 476.660 52.030 476.920 52.350 ;
        RECT 904.920 52.030 905.180 52.350 ;
        RECT 904.980 1.770 905.120 52.030 ;
        RECT 907.070 1.770 907.630 2.400 ;
        RECT 904.980 1.630 907.630 1.770 ;
        RECT 907.070 -4.800 907.630 1.630 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.990 51.920 484.310 51.980 ;
        RECT 925.590 51.920 925.910 51.980 ;
        RECT 483.990 51.780 925.910 51.920 ;
        RECT 483.990 51.720 484.310 51.780 ;
        RECT 925.590 51.720 925.910 51.780 ;
      LAYER via ;
        RECT 484.020 51.720 484.280 51.980 ;
        RECT 925.620 51.720 925.880 51.980 ;
      LAYER met2 ;
        RECT 483.450 400.250 483.730 404.000 ;
        RECT 483.450 400.110 485.140 400.250 ;
        RECT 483.450 400.000 483.730 400.110 ;
        RECT 485.000 324.370 485.140 400.110 ;
        RECT 484.080 324.230 485.140 324.370 ;
        RECT 484.080 52.010 484.220 324.230 ;
        RECT 484.020 51.690 484.280 52.010 ;
        RECT 925.620 51.690 925.880 52.010 ;
        RECT 925.680 17.410 925.820 51.690 ;
        RECT 924.760 17.270 925.820 17.410 ;
        RECT 924.760 2.400 924.900 17.270 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 483.530 376.280 483.850 376.340 ;
        RECT 487.670 376.280 487.990 376.340 ;
        RECT 483.530 376.140 487.990 376.280 ;
        RECT 483.530 376.080 483.850 376.140 ;
        RECT 487.670 376.080 487.990 376.140 ;
        RECT 483.530 43.080 483.850 43.140 ;
        RECT 942.610 43.080 942.930 43.140 ;
        RECT 483.530 42.940 942.930 43.080 ;
        RECT 483.530 42.880 483.850 42.940 ;
        RECT 942.610 42.880 942.930 42.940 ;
      LAYER via ;
        RECT 483.560 376.080 483.820 376.340 ;
        RECT 487.700 376.080 487.960 376.340 ;
        RECT 483.560 42.880 483.820 43.140 ;
        RECT 942.640 42.880 942.900 43.140 ;
      LAYER met2 ;
        RECT 488.970 400.250 489.250 404.000 ;
        RECT 487.760 400.110 489.250 400.250 ;
        RECT 487.760 376.370 487.900 400.110 ;
        RECT 488.970 400.000 489.250 400.110 ;
        RECT 483.560 376.050 483.820 376.370 ;
        RECT 487.700 376.050 487.960 376.370 ;
        RECT 483.620 43.170 483.760 376.050 ;
        RECT 483.560 42.850 483.820 43.170 ;
        RECT 942.640 42.850 942.900 43.170 ;
        RECT 942.700 2.400 942.840 42.850 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 490.890 49.540 491.210 49.600 ;
        RECT 960.090 49.540 960.410 49.600 ;
        RECT 490.890 49.400 960.410 49.540 ;
        RECT 490.890 49.340 491.210 49.400 ;
        RECT 960.090 49.340 960.410 49.400 ;
      LAYER via ;
        RECT 490.920 49.340 491.180 49.600 ;
        RECT 960.120 49.340 960.380 49.600 ;
      LAYER met2 ;
        RECT 494.490 400.250 494.770 404.000 ;
        RECT 493.280 400.110 494.770 400.250 ;
        RECT 493.280 399.570 493.420 400.110 ;
        RECT 494.490 400.000 494.770 400.110 ;
        RECT 492.820 399.430 493.420 399.570 ;
        RECT 492.820 351.970 492.960 399.430 ;
        RECT 490.980 351.830 492.960 351.970 ;
        RECT 490.980 49.630 491.120 351.830 ;
        RECT 490.920 49.310 491.180 49.630 ;
        RECT 960.120 49.310 960.380 49.630 ;
        RECT 960.180 2.400 960.320 49.310 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 497.790 60.760 498.110 60.820 ;
        RECT 975.730 60.760 976.050 60.820 ;
        RECT 497.790 60.620 976.050 60.760 ;
        RECT 497.790 60.560 498.110 60.620 ;
        RECT 975.730 60.560 976.050 60.620 ;
      LAYER via ;
        RECT 497.820 60.560 498.080 60.820 ;
        RECT 975.760 60.560 976.020 60.820 ;
      LAYER met2 ;
        RECT 500.010 400.250 500.290 404.000 ;
        RECT 498.800 400.110 500.290 400.250 ;
        RECT 498.800 324.370 498.940 400.110 ;
        RECT 500.010 400.000 500.290 400.110 ;
        RECT 497.880 324.230 498.940 324.370 ;
        RECT 497.880 60.850 498.020 324.230 ;
        RECT 497.820 60.530 498.080 60.850 ;
        RECT 975.760 60.530 976.020 60.850 ;
        RECT 975.820 1.770 975.960 60.530 ;
        RECT 977.910 1.770 978.470 2.400 ;
        RECT 975.820 1.630 978.470 1.770 ;
        RECT 977.910 -4.800 978.470 1.630 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 401.650 391.240 401.970 391.300 ;
        RECT 616.930 391.240 617.250 391.300 ;
        RECT 401.650 391.100 617.250 391.240 ;
        RECT 401.650 391.040 401.970 391.100 ;
        RECT 616.930 391.040 617.250 391.100 ;
        RECT 616.930 16.900 617.250 16.960 ;
        RECT 658.790 16.900 659.110 16.960 ;
        RECT 616.930 16.760 659.110 16.900 ;
        RECT 616.930 16.700 617.250 16.760 ;
        RECT 658.790 16.700 659.110 16.760 ;
      LAYER via ;
        RECT 401.680 391.040 401.940 391.300 ;
        RECT 616.960 391.040 617.220 391.300 ;
        RECT 616.960 16.700 617.220 16.960 ;
        RECT 658.820 16.700 659.080 16.960 ;
      LAYER met2 ;
        RECT 401.570 400.180 401.850 404.000 ;
        RECT 401.570 400.000 401.880 400.180 ;
        RECT 401.740 391.330 401.880 400.000 ;
        RECT 401.680 391.010 401.940 391.330 ;
        RECT 616.960 391.010 617.220 391.330 ;
        RECT 617.020 351.970 617.160 391.010 ;
        RECT 617.020 351.830 617.620 351.970 ;
        RECT 617.480 34.570 617.620 351.830 ;
        RECT 617.020 34.430 617.620 34.570 ;
        RECT 617.020 16.990 617.160 34.430 ;
        RECT 616.960 16.670 617.220 16.990 ;
        RECT 658.820 16.670 659.080 16.990 ;
        RECT 658.880 2.400 659.020 16.670 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 504.690 60.420 505.010 60.480 ;
        RECT 994.590 60.420 994.910 60.480 ;
        RECT 504.690 60.280 994.910 60.420 ;
        RECT 504.690 60.220 505.010 60.280 ;
        RECT 994.590 60.220 994.910 60.280 ;
      LAYER via ;
        RECT 504.720 60.220 504.980 60.480 ;
        RECT 994.620 60.220 994.880 60.480 ;
      LAYER met2 ;
        RECT 505.070 400.250 505.350 404.000 ;
        RECT 504.780 400.110 505.350 400.250 ;
        RECT 504.780 60.510 504.920 400.110 ;
        RECT 505.070 400.000 505.350 400.110 ;
        RECT 504.720 60.190 504.980 60.510 ;
        RECT 994.620 60.190 994.880 60.510 ;
        RECT 994.680 1.770 994.820 60.190 ;
        RECT 995.390 1.770 995.950 2.400 ;
        RECT 994.680 1.630 995.950 1.770 ;
        RECT 995.390 -4.800 995.950 1.630 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.130 60.080 511.450 60.140 ;
        RECT 1008.850 60.080 1009.170 60.140 ;
        RECT 511.130 59.940 1009.170 60.080 ;
        RECT 511.130 59.880 511.450 59.940 ;
        RECT 1008.850 59.880 1009.170 59.940 ;
      LAYER via ;
        RECT 511.160 59.880 511.420 60.140 ;
        RECT 1008.880 59.880 1009.140 60.140 ;
      LAYER met2 ;
        RECT 510.590 400.250 510.870 404.000 ;
        RECT 510.590 400.110 511.360 400.250 ;
        RECT 510.590 400.000 510.870 400.110 ;
        RECT 511.220 60.170 511.360 400.110 ;
        RECT 511.160 59.850 511.420 60.170 ;
        RECT 1008.880 59.850 1009.140 60.170 ;
        RECT 1008.940 17.410 1009.080 59.850 ;
        RECT 1008.940 17.270 1013.680 17.410 ;
        RECT 1013.540 2.400 1013.680 17.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.590 59.400 511.910 59.460 ;
        RECT 1030.930 59.400 1031.250 59.460 ;
        RECT 511.590 59.260 1031.250 59.400 ;
        RECT 511.590 59.200 511.910 59.260 ;
        RECT 1030.930 59.200 1031.250 59.260 ;
      LAYER via ;
        RECT 511.620 59.200 511.880 59.460 ;
        RECT 1030.960 59.200 1031.220 59.460 ;
      LAYER met2 ;
        RECT 516.110 400.250 516.390 404.000 ;
        RECT 514.900 400.110 516.390 400.250 ;
        RECT 514.900 388.690 515.040 400.110 ;
        RECT 516.110 400.000 516.390 400.110 ;
        RECT 512.600 388.550 515.040 388.690 ;
        RECT 512.600 324.370 512.740 388.550 ;
        RECT 511.680 324.230 512.740 324.370 ;
        RECT 511.680 59.490 511.820 324.230 ;
        RECT 511.620 59.170 511.880 59.490 ;
        RECT 1030.960 59.170 1031.220 59.490 ;
        RECT 1031.020 2.400 1031.160 59.170 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 518.030 386.480 518.350 386.540 ;
        RECT 520.330 386.480 520.650 386.540 ;
        RECT 518.030 386.340 520.650 386.480 ;
        RECT 518.030 386.280 518.350 386.340 ;
        RECT 520.330 386.280 520.650 386.340 ;
        RECT 518.030 59.060 518.350 59.120 ;
        RECT 1048.870 59.060 1049.190 59.120 ;
        RECT 518.030 58.920 1049.190 59.060 ;
        RECT 518.030 58.860 518.350 58.920 ;
        RECT 1048.870 58.860 1049.190 58.920 ;
      LAYER via ;
        RECT 518.060 386.280 518.320 386.540 ;
        RECT 520.360 386.280 520.620 386.540 ;
        RECT 518.060 58.860 518.320 59.120 ;
        RECT 1048.900 58.860 1049.160 59.120 ;
      LAYER met2 ;
        RECT 521.630 400.250 521.910 404.000 ;
        RECT 520.420 400.110 521.910 400.250 ;
        RECT 520.420 386.570 520.560 400.110 ;
        RECT 521.630 400.000 521.910 400.110 ;
        RECT 518.060 386.250 518.320 386.570 ;
        RECT 520.360 386.250 520.620 386.570 ;
        RECT 518.120 59.150 518.260 386.250 ;
        RECT 518.060 58.830 518.320 59.150 ;
        RECT 1048.900 58.830 1049.160 59.150 ;
        RECT 1048.960 2.400 1049.100 58.830 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 524.470 56.340 524.790 56.400 ;
        RECT 1066.810 56.340 1067.130 56.400 ;
        RECT 524.470 56.200 1067.130 56.340 ;
        RECT 524.470 56.140 524.790 56.200 ;
        RECT 1066.810 56.140 1067.130 56.200 ;
      LAYER via ;
        RECT 524.500 56.140 524.760 56.400 ;
        RECT 1066.840 56.140 1067.100 56.400 ;
      LAYER met2 ;
        RECT 527.150 400.250 527.430 404.000 ;
        RECT 525.940 400.110 527.430 400.250 ;
        RECT 525.940 386.470 526.080 400.110 ;
        RECT 527.150 400.000 527.430 400.110 ;
        RECT 524.560 386.330 526.080 386.470 ;
        RECT 524.560 56.430 524.700 386.330 ;
        RECT 524.500 56.110 524.760 56.430 ;
        RECT 1066.840 56.110 1067.100 56.430 ;
        RECT 1066.900 2.400 1067.040 56.110 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 531.830 58.720 532.150 58.780 ;
        RECT 1083.370 58.720 1083.690 58.780 ;
        RECT 531.830 58.580 1083.690 58.720 ;
        RECT 531.830 58.520 532.150 58.580 ;
        RECT 1083.370 58.520 1083.690 58.580 ;
      LAYER via ;
        RECT 531.860 58.520 532.120 58.780 ;
        RECT 1083.400 58.520 1083.660 58.780 ;
      LAYER met2 ;
        RECT 532.670 400.250 532.950 404.000 ;
        RECT 531.920 400.110 532.950 400.250 ;
        RECT 531.920 58.810 532.060 400.110 ;
        RECT 532.670 400.000 532.950 400.110 ;
        RECT 531.860 58.490 532.120 58.810 ;
        RECT 1083.400 58.490 1083.660 58.810 ;
        RECT 1083.460 17.410 1083.600 58.490 ;
        RECT 1083.460 17.270 1084.520 17.410 ;
        RECT 1084.380 2.400 1084.520 17.270 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 532.290 386.480 532.610 386.540 ;
        RECT 536.430 386.480 536.750 386.540 ;
        RECT 532.290 386.340 536.750 386.480 ;
        RECT 532.290 386.280 532.610 386.340 ;
        RECT 536.430 386.280 536.750 386.340 ;
        RECT 532.290 77.760 532.610 77.820 ;
        RECT 1099.930 77.760 1100.250 77.820 ;
        RECT 532.290 77.620 1100.250 77.760 ;
        RECT 532.290 77.560 532.610 77.620 ;
        RECT 1099.930 77.560 1100.250 77.620 ;
      LAYER via ;
        RECT 532.320 386.280 532.580 386.540 ;
        RECT 536.460 386.280 536.720 386.540 ;
        RECT 532.320 77.560 532.580 77.820 ;
        RECT 1099.960 77.560 1100.220 77.820 ;
      LAYER met2 ;
        RECT 537.730 400.250 538.010 404.000 ;
        RECT 536.520 400.110 538.010 400.250 ;
        RECT 536.520 386.570 536.660 400.110 ;
        RECT 537.730 400.000 538.010 400.110 ;
        RECT 532.320 386.250 532.580 386.570 ;
        RECT 536.460 386.250 536.720 386.570 ;
        RECT 532.380 77.850 532.520 386.250 ;
        RECT 532.320 77.530 532.580 77.850 ;
        RECT 1099.960 77.530 1100.220 77.850 ;
        RECT 1100.020 1.770 1100.160 77.530 ;
        RECT 1102.110 1.770 1102.670 2.400 ;
        RECT 1100.020 1.630 1102.670 1.770 ;
        RECT 1102.110 -4.800 1102.670 1.630 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.270 386.480 538.590 386.540 ;
        RECT 541.950 386.480 542.270 386.540 ;
        RECT 538.270 386.340 542.270 386.480 ;
        RECT 538.270 386.280 538.590 386.340 ;
        RECT 541.950 386.280 542.270 386.340 ;
        RECT 538.270 84.560 538.590 84.620 ;
        RECT 1117.870 84.560 1118.190 84.620 ;
        RECT 538.270 84.420 1118.190 84.560 ;
        RECT 538.270 84.360 538.590 84.420 ;
        RECT 1117.870 84.360 1118.190 84.420 ;
      LAYER via ;
        RECT 538.300 386.280 538.560 386.540 ;
        RECT 541.980 386.280 542.240 386.540 ;
        RECT 538.300 84.360 538.560 84.620 ;
        RECT 1117.900 84.360 1118.160 84.620 ;
      LAYER met2 ;
        RECT 543.250 400.250 543.530 404.000 ;
        RECT 542.040 400.110 543.530 400.250 ;
        RECT 542.040 386.570 542.180 400.110 ;
        RECT 543.250 400.000 543.530 400.110 ;
        RECT 538.300 386.250 538.560 386.570 ;
        RECT 541.980 386.250 542.240 386.570 ;
        RECT 538.360 84.650 538.500 386.250 ;
        RECT 538.300 84.330 538.560 84.650 ;
        RECT 1117.900 84.330 1118.160 84.650 ;
        RECT 1117.960 1.770 1118.100 84.330 ;
        RECT 1119.590 1.770 1120.150 2.400 ;
        RECT 1117.960 1.630 1120.150 1.770 ;
        RECT 1119.590 -4.800 1120.150 1.630 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 546.090 376.280 546.410 376.340 ;
        RECT 547.470 376.280 547.790 376.340 ;
        RECT 546.090 376.140 547.790 376.280 ;
        RECT 546.090 376.080 546.410 376.140 ;
        RECT 547.470 376.080 547.790 376.140 ;
        RECT 546.090 91.360 546.410 91.420 ;
        RECT 1132.130 91.360 1132.450 91.420 ;
        RECT 546.090 91.220 1132.450 91.360 ;
        RECT 546.090 91.160 546.410 91.220 ;
        RECT 1132.130 91.160 1132.450 91.220 ;
      LAYER via ;
        RECT 546.120 376.080 546.380 376.340 ;
        RECT 547.500 376.080 547.760 376.340 ;
        RECT 546.120 91.160 546.380 91.420 ;
        RECT 1132.160 91.160 1132.420 91.420 ;
      LAYER met2 ;
        RECT 548.770 400.250 549.050 404.000 ;
        RECT 547.560 400.110 549.050 400.250 ;
        RECT 547.560 376.370 547.700 400.110 ;
        RECT 548.770 400.000 549.050 400.110 ;
        RECT 546.120 376.050 546.380 376.370 ;
        RECT 547.500 376.050 547.760 376.370 ;
        RECT 546.180 91.450 546.320 376.050 ;
        RECT 546.120 91.130 546.380 91.450 ;
        RECT 1132.160 91.130 1132.420 91.450 ;
        RECT 1132.220 82.870 1132.360 91.130 ;
        RECT 1132.220 82.730 1137.880 82.870 ;
        RECT 1137.740 2.400 1137.880 82.730 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 552.530 376.280 552.850 376.340 ;
        RECT 553.450 376.280 553.770 376.340 ;
        RECT 552.530 376.140 553.770 376.280 ;
        RECT 552.530 376.080 552.850 376.140 ;
        RECT 553.450 376.080 553.770 376.140 ;
        RECT 552.530 91.700 552.850 91.760 ;
        RECT 1152.370 91.700 1152.690 91.760 ;
        RECT 552.530 91.560 1152.690 91.700 ;
        RECT 552.530 91.500 552.850 91.560 ;
        RECT 1152.370 91.500 1152.690 91.560 ;
      LAYER via ;
        RECT 552.560 376.080 552.820 376.340 ;
        RECT 553.480 376.080 553.740 376.340 ;
        RECT 552.560 91.500 552.820 91.760 ;
        RECT 1152.400 91.500 1152.660 91.760 ;
      LAYER met2 ;
        RECT 554.290 400.250 554.570 404.000 ;
        RECT 553.540 400.110 554.570 400.250 ;
        RECT 553.540 376.370 553.680 400.110 ;
        RECT 554.290 400.000 554.570 400.110 ;
        RECT 552.560 376.050 552.820 376.370 ;
        RECT 553.480 376.050 553.740 376.370 ;
        RECT 552.620 91.790 552.760 376.050 ;
        RECT 552.560 91.470 552.820 91.790 ;
        RECT 1152.400 91.470 1152.660 91.790 ;
        RECT 1152.460 82.870 1152.600 91.470 ;
        RECT 1152.460 82.730 1155.360 82.870 ;
        RECT 1155.220 2.400 1155.360 82.730 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.090 38.660 408.410 38.720 ;
        RECT 676.270 38.660 676.590 38.720 ;
        RECT 408.090 38.520 676.590 38.660 ;
        RECT 408.090 38.460 408.410 38.520 ;
        RECT 676.270 38.460 676.590 38.520 ;
      LAYER via ;
        RECT 408.120 38.460 408.380 38.720 ;
        RECT 676.300 38.460 676.560 38.720 ;
      LAYER met2 ;
        RECT 407.090 400.250 407.370 404.000 ;
        RECT 407.090 400.110 408.320 400.250 ;
        RECT 407.090 400.000 407.370 400.110 ;
        RECT 408.180 38.750 408.320 400.110 ;
        RECT 408.120 38.430 408.380 38.750 ;
        RECT 676.300 38.430 676.560 38.750 ;
        RECT 676.360 2.400 676.500 38.430 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 559.890 92.040 560.210 92.100 ;
        RECT 1173.070 92.040 1173.390 92.100 ;
        RECT 559.890 91.900 1173.390 92.040 ;
        RECT 559.890 91.840 560.210 91.900 ;
        RECT 1173.070 91.840 1173.390 91.900 ;
      LAYER via ;
        RECT 559.920 91.840 560.180 92.100 ;
        RECT 1173.100 91.840 1173.360 92.100 ;
      LAYER met2 ;
        RECT 559.810 400.250 560.090 404.000 ;
        RECT 559.520 400.110 560.090 400.250 ;
        RECT 559.520 386.470 559.660 400.110 ;
        RECT 559.810 400.000 560.090 400.110 ;
        RECT 559.520 386.330 560.120 386.470 ;
        RECT 559.980 92.130 560.120 386.330 ;
        RECT 559.920 91.810 560.180 92.130 ;
        RECT 1173.100 91.810 1173.360 92.130 ;
        RECT 1173.160 2.400 1173.300 91.810 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.350 92.380 560.670 92.440 ;
        RECT 1186.870 92.380 1187.190 92.440 ;
        RECT 560.350 92.240 1187.190 92.380 ;
        RECT 560.350 92.180 560.670 92.240 ;
        RECT 1186.870 92.180 1187.190 92.240 ;
      LAYER via ;
        RECT 560.380 92.180 560.640 92.440 ;
        RECT 1186.900 92.180 1187.160 92.440 ;
      LAYER met2 ;
        RECT 565.330 400.250 565.610 404.000 ;
        RECT 564.120 400.110 565.610 400.250 ;
        RECT 564.120 324.370 564.260 400.110 ;
        RECT 565.330 400.000 565.610 400.110 ;
        RECT 560.440 324.230 564.260 324.370 ;
        RECT 560.440 92.470 560.580 324.230 ;
        RECT 560.380 92.150 560.640 92.470 ;
        RECT 1186.900 92.150 1187.160 92.470 ;
        RECT 1186.960 82.870 1187.100 92.150 ;
        RECT 1186.960 82.730 1188.480 82.870 ;
        RECT 1188.340 1.770 1188.480 82.730 ;
        RECT 1190.430 1.770 1190.990 2.400 ;
        RECT 1188.340 1.630 1190.990 1.770 ;
        RECT 1190.430 -4.800 1190.990 1.630 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 567.250 92.720 567.570 92.780 ;
        RECT 1207.570 92.720 1207.890 92.780 ;
        RECT 567.250 92.580 1207.890 92.720 ;
        RECT 567.250 92.520 567.570 92.580 ;
        RECT 1207.570 92.520 1207.890 92.580 ;
      LAYER via ;
        RECT 567.280 92.520 567.540 92.780 ;
        RECT 1207.600 92.520 1207.860 92.780 ;
      LAYER met2 ;
        RECT 570.390 400.250 570.670 404.000 ;
        RECT 569.180 400.110 570.670 400.250 ;
        RECT 569.180 324.370 569.320 400.110 ;
        RECT 570.390 400.000 570.670 400.110 ;
        RECT 567.340 324.230 569.320 324.370 ;
        RECT 567.340 92.810 567.480 324.230 ;
        RECT 567.280 92.490 567.540 92.810 ;
        RECT 1207.600 92.490 1207.860 92.810 ;
        RECT 1207.660 82.870 1207.800 92.490 ;
        RECT 1207.660 82.730 1208.720 82.870 ;
        RECT 1208.580 2.400 1208.720 82.730 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 573.690 96.460 574.010 96.520 ;
        RECT 1221.370 96.460 1221.690 96.520 ;
        RECT 573.690 96.320 1221.690 96.460 ;
        RECT 573.690 96.260 574.010 96.320 ;
        RECT 1221.370 96.260 1221.690 96.320 ;
      LAYER via ;
        RECT 573.720 96.260 573.980 96.520 ;
        RECT 1221.400 96.260 1221.660 96.520 ;
      LAYER met2 ;
        RECT 575.910 400.250 576.190 404.000 ;
        RECT 574.700 400.110 576.190 400.250 ;
        RECT 574.700 324.370 574.840 400.110 ;
        RECT 575.910 400.000 576.190 400.110 ;
        RECT 573.780 324.230 574.840 324.370 ;
        RECT 573.780 96.550 573.920 324.230 ;
        RECT 573.720 96.230 573.980 96.550 ;
        RECT 1221.400 96.230 1221.660 96.550 ;
        RECT 1221.460 82.870 1221.600 96.230 ;
        RECT 1221.460 82.730 1226.200 82.870 ;
        RECT 1226.060 2.400 1226.200 82.730 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 581.050 96.120 581.370 96.180 ;
        RECT 1242.070 96.120 1242.390 96.180 ;
        RECT 581.050 95.980 1242.390 96.120 ;
        RECT 581.050 95.920 581.370 95.980 ;
        RECT 1242.070 95.920 1242.390 95.980 ;
      LAYER via ;
        RECT 581.080 95.920 581.340 96.180 ;
        RECT 1242.100 95.920 1242.360 96.180 ;
      LAYER met2 ;
        RECT 581.430 400.250 581.710 404.000 ;
        RECT 581.140 400.110 581.710 400.250 ;
        RECT 581.140 96.210 581.280 400.110 ;
        RECT 581.430 400.000 581.710 400.110 ;
        RECT 581.080 95.890 581.340 96.210 ;
        RECT 1242.100 95.890 1242.360 96.210 ;
        RECT 1242.160 1.770 1242.300 95.890 ;
        RECT 1243.790 1.770 1244.350 2.400 ;
        RECT 1242.160 1.630 1244.350 1.770 ;
        RECT 1243.790 -4.800 1244.350 1.630 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.950 95.780 588.270 95.840 ;
        RECT 1255.870 95.780 1256.190 95.840 ;
        RECT 587.950 95.640 1256.190 95.780 ;
        RECT 587.950 95.580 588.270 95.640 ;
        RECT 1255.870 95.580 1256.190 95.640 ;
        RECT 1255.870 20.980 1256.190 21.040 ;
        RECT 1261.850 20.980 1262.170 21.040 ;
        RECT 1255.870 20.840 1262.170 20.980 ;
        RECT 1255.870 20.780 1256.190 20.840 ;
        RECT 1261.850 20.780 1262.170 20.840 ;
      LAYER via ;
        RECT 587.980 95.580 588.240 95.840 ;
        RECT 1255.900 95.580 1256.160 95.840 ;
        RECT 1255.900 20.780 1256.160 21.040 ;
        RECT 1261.880 20.780 1262.140 21.040 ;
      LAYER met2 ;
        RECT 586.950 400.250 587.230 404.000 ;
        RECT 586.950 400.110 588.640 400.250 ;
        RECT 586.950 400.000 587.230 400.110 ;
        RECT 588.500 351.970 588.640 400.110 ;
        RECT 588.500 351.830 589.100 351.970 ;
        RECT 588.960 324.370 589.100 351.830 ;
        RECT 588.040 324.230 589.100 324.370 ;
        RECT 588.040 95.870 588.180 324.230 ;
        RECT 587.980 95.550 588.240 95.870 ;
        RECT 1255.900 95.550 1256.160 95.870 ;
        RECT 1255.960 21.070 1256.100 95.550 ;
        RECT 1255.900 20.750 1256.160 21.070 ;
        RECT 1261.880 20.750 1262.140 21.070 ;
        RECT 1261.940 2.400 1262.080 20.750 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 587.490 376.280 587.810 376.340 ;
        RECT 591.170 376.280 591.490 376.340 ;
        RECT 587.490 376.140 591.490 376.280 ;
        RECT 587.490 376.080 587.810 376.140 ;
        RECT 591.170 376.080 591.490 376.140 ;
        RECT 587.490 95.440 587.810 95.500 ;
        RECT 1276.570 95.440 1276.890 95.500 ;
        RECT 587.490 95.300 1276.890 95.440 ;
        RECT 587.490 95.240 587.810 95.300 ;
        RECT 1276.570 95.240 1276.890 95.300 ;
      LAYER via ;
        RECT 587.520 376.080 587.780 376.340 ;
        RECT 591.200 376.080 591.460 376.340 ;
        RECT 587.520 95.240 587.780 95.500 ;
        RECT 1276.600 95.240 1276.860 95.500 ;
      LAYER met2 ;
        RECT 592.470 400.250 592.750 404.000 ;
        RECT 591.260 400.110 592.750 400.250 ;
        RECT 591.260 376.370 591.400 400.110 ;
        RECT 592.470 400.000 592.750 400.110 ;
        RECT 587.520 376.050 587.780 376.370 ;
        RECT 591.200 376.050 591.460 376.370 ;
        RECT 587.580 95.530 587.720 376.050 ;
        RECT 587.520 95.210 587.780 95.530 ;
        RECT 1276.600 95.210 1276.860 95.530 ;
        RECT 1276.660 82.870 1276.800 95.210 ;
        RECT 1276.660 82.730 1279.560 82.870 ;
        RECT 1279.420 2.400 1279.560 82.730 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 594.850 98.160 595.170 98.220 ;
        RECT 1297.270 98.160 1297.590 98.220 ;
        RECT 594.850 98.020 1297.590 98.160 ;
        RECT 594.850 97.960 595.170 98.020 ;
        RECT 1297.270 97.960 1297.590 98.020 ;
      LAYER via ;
        RECT 594.880 97.960 595.140 98.220 ;
        RECT 1297.300 97.960 1297.560 98.220 ;
      LAYER met2 ;
        RECT 597.990 400.250 598.270 404.000 ;
        RECT 596.780 400.110 598.270 400.250 ;
        RECT 596.780 399.570 596.920 400.110 ;
        RECT 597.990 400.000 598.270 400.110 ;
        RECT 595.860 399.430 596.920 399.570 ;
        RECT 595.860 324.370 596.000 399.430 ;
        RECT 594.940 324.230 596.000 324.370 ;
        RECT 594.940 98.250 595.080 324.230 ;
        RECT 594.880 97.930 595.140 98.250 ;
        RECT 1297.300 97.930 1297.560 98.250 ;
        RECT 1297.360 2.400 1297.500 97.930 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 601.750 98.500 602.070 98.560 ;
        RECT 1311.070 98.500 1311.390 98.560 ;
        RECT 601.750 98.360 1311.390 98.500 ;
        RECT 601.750 98.300 602.070 98.360 ;
        RECT 1311.070 98.300 1311.390 98.360 ;
      LAYER via ;
        RECT 601.780 98.300 602.040 98.560 ;
        RECT 1311.100 98.300 1311.360 98.560 ;
      LAYER met2 ;
        RECT 603.050 400.250 603.330 404.000 ;
        RECT 601.840 400.110 603.330 400.250 ;
        RECT 601.840 98.590 601.980 400.110 ;
        RECT 603.050 400.000 603.330 400.110 ;
        RECT 601.780 98.270 602.040 98.590 ;
        RECT 1311.100 98.270 1311.360 98.590 ;
        RECT 1311.160 82.870 1311.300 98.270 ;
        RECT 1311.160 82.730 1312.680 82.870 ;
        RECT 1312.540 1.770 1312.680 82.730 ;
        RECT 1314.630 1.770 1315.190 2.400 ;
        RECT 1312.540 1.630 1315.190 1.770 ;
        RECT 1314.630 -4.800 1315.190 1.630 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 607.730 98.840 608.050 98.900 ;
        RECT 1331.770 98.840 1332.090 98.900 ;
        RECT 607.730 98.700 1332.090 98.840 ;
        RECT 607.730 98.640 608.050 98.700 ;
        RECT 1331.770 98.640 1332.090 98.700 ;
      LAYER via ;
        RECT 607.760 98.640 608.020 98.900 ;
        RECT 1331.800 98.640 1332.060 98.900 ;
      LAYER met2 ;
        RECT 608.570 400.250 608.850 404.000 ;
        RECT 607.820 400.110 608.850 400.250 ;
        RECT 607.820 98.930 607.960 400.110 ;
        RECT 608.570 400.000 608.850 400.110 ;
        RECT 607.760 98.610 608.020 98.930 ;
        RECT 1331.800 98.610 1332.060 98.930 ;
        RECT 1331.860 82.870 1332.000 98.610 ;
        RECT 1331.860 82.730 1332.920 82.870 ;
        RECT 1332.780 2.400 1332.920 82.730 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 407.630 386.140 407.950 386.200 ;
        RECT 411.310 386.140 411.630 386.200 ;
        RECT 407.630 386.000 411.630 386.140 ;
        RECT 407.630 385.940 407.950 386.000 ;
        RECT 411.310 385.940 411.630 386.000 ;
        RECT 407.630 32.540 407.950 32.600 ;
        RECT 553.450 32.540 553.770 32.600 ;
        RECT 407.630 32.400 553.770 32.540 ;
        RECT 407.630 32.340 407.950 32.400 ;
        RECT 553.450 32.340 553.770 32.400 ;
        RECT 553.450 16.220 553.770 16.280 ;
        RECT 694.210 16.220 694.530 16.280 ;
        RECT 553.450 16.080 694.530 16.220 ;
        RECT 553.450 16.020 553.770 16.080 ;
        RECT 694.210 16.020 694.530 16.080 ;
      LAYER via ;
        RECT 407.660 385.940 407.920 386.200 ;
        RECT 411.340 385.940 411.600 386.200 ;
        RECT 407.660 32.340 407.920 32.600 ;
        RECT 553.480 32.340 553.740 32.600 ;
        RECT 553.480 16.020 553.740 16.280 ;
        RECT 694.240 16.020 694.500 16.280 ;
      LAYER met2 ;
        RECT 412.610 400.250 412.890 404.000 ;
        RECT 411.400 400.110 412.890 400.250 ;
        RECT 411.400 386.230 411.540 400.110 ;
        RECT 412.610 400.000 412.890 400.110 ;
        RECT 407.660 385.910 407.920 386.230 ;
        RECT 411.340 385.910 411.600 386.230 ;
        RECT 407.720 32.630 407.860 385.910 ;
        RECT 407.660 32.310 407.920 32.630 ;
        RECT 553.480 32.310 553.740 32.630 ;
        RECT 553.540 16.310 553.680 32.310 ;
        RECT 553.480 15.990 553.740 16.310 ;
        RECT 694.240 15.990 694.500 16.310 ;
        RECT 694.300 2.400 694.440 15.990 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 615.090 99.180 615.410 99.240 ;
        RECT 1345.570 99.180 1345.890 99.240 ;
        RECT 615.090 99.040 1345.890 99.180 ;
        RECT 615.090 98.980 615.410 99.040 ;
        RECT 1345.570 98.980 1345.890 99.040 ;
      LAYER via ;
        RECT 615.120 98.980 615.380 99.240 ;
        RECT 1345.600 98.980 1345.860 99.240 ;
      LAYER met2 ;
        RECT 614.090 400.250 614.370 404.000 ;
        RECT 614.090 400.110 615.320 400.250 ;
        RECT 614.090 400.000 614.370 400.110 ;
        RECT 615.180 99.270 615.320 400.110 ;
        RECT 615.120 98.950 615.380 99.270 ;
        RECT 1345.600 98.950 1345.860 99.270 ;
        RECT 1345.660 82.870 1345.800 98.950 ;
        RECT 1345.660 82.730 1350.400 82.870 ;
        RECT 1350.260 2.400 1350.400 82.730 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 614.630 376.280 614.950 376.340 ;
        RECT 618.310 376.280 618.630 376.340 ;
        RECT 614.630 376.140 618.630 376.280 ;
        RECT 614.630 376.080 614.950 376.140 ;
        RECT 618.310 376.080 618.630 376.140 ;
        RECT 614.630 99.520 614.950 99.580 ;
        RECT 1366.270 99.520 1366.590 99.580 ;
        RECT 614.630 99.380 1366.590 99.520 ;
        RECT 614.630 99.320 614.950 99.380 ;
        RECT 1366.270 99.320 1366.590 99.380 ;
      LAYER via ;
        RECT 614.660 376.080 614.920 376.340 ;
        RECT 618.340 376.080 618.600 376.340 ;
        RECT 614.660 99.320 614.920 99.580 ;
        RECT 1366.300 99.320 1366.560 99.580 ;
      LAYER met2 ;
        RECT 619.610 400.250 619.890 404.000 ;
        RECT 618.400 400.110 619.890 400.250 ;
        RECT 618.400 376.370 618.540 400.110 ;
        RECT 619.610 400.000 619.890 400.110 ;
        RECT 614.660 376.050 614.920 376.370 ;
        RECT 618.340 376.050 618.600 376.370 ;
        RECT 614.720 99.610 614.860 376.050 ;
        RECT 614.660 99.290 614.920 99.610 ;
        RECT 1366.300 99.290 1366.560 99.610 ;
        RECT 1366.360 1.770 1366.500 99.290 ;
        RECT 1367.990 1.770 1368.550 2.400 ;
        RECT 1366.360 1.630 1368.550 1.770 ;
        RECT 1367.990 -4.800 1368.550 1.630 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.530 375.940 621.850 376.000 ;
        RECT 623.830 375.940 624.150 376.000 ;
        RECT 621.530 375.800 624.150 375.940 ;
        RECT 621.530 375.740 621.850 375.800 ;
        RECT 623.830 375.740 624.150 375.800 ;
        RECT 621.530 103.260 621.850 103.320 ;
        RECT 1380.070 103.260 1380.390 103.320 ;
        RECT 621.530 103.120 1380.390 103.260 ;
        RECT 621.530 103.060 621.850 103.120 ;
        RECT 1380.070 103.060 1380.390 103.120 ;
        RECT 1380.070 20.980 1380.390 21.040 ;
        RECT 1383.750 20.980 1384.070 21.040 ;
        RECT 1380.070 20.840 1384.070 20.980 ;
        RECT 1380.070 20.780 1380.390 20.840 ;
        RECT 1383.750 20.780 1384.070 20.840 ;
      LAYER via ;
        RECT 621.560 375.740 621.820 376.000 ;
        RECT 623.860 375.740 624.120 376.000 ;
        RECT 621.560 103.060 621.820 103.320 ;
        RECT 1380.100 103.060 1380.360 103.320 ;
        RECT 1380.100 20.780 1380.360 21.040 ;
        RECT 1383.780 20.780 1384.040 21.040 ;
      LAYER met2 ;
        RECT 625.130 400.250 625.410 404.000 ;
        RECT 623.920 400.110 625.410 400.250 ;
        RECT 623.920 376.030 624.060 400.110 ;
        RECT 625.130 400.000 625.410 400.110 ;
        RECT 621.560 375.710 621.820 376.030 ;
        RECT 623.860 375.710 624.120 376.030 ;
        RECT 621.620 103.350 621.760 375.710 ;
        RECT 621.560 103.030 621.820 103.350 ;
        RECT 1380.100 103.030 1380.360 103.350 ;
        RECT 1380.160 21.070 1380.300 103.030 ;
        RECT 1380.100 20.750 1380.360 21.070 ;
        RECT 1383.780 20.750 1384.040 21.070 ;
        RECT 1383.840 1.770 1383.980 20.750 ;
        RECT 1385.470 1.770 1386.030 2.400 ;
        RECT 1383.840 1.630 1386.030 1.770 ;
        RECT 1385.470 -4.800 1386.030 1.630 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 628.890 102.920 629.210 102.980 ;
        RECT 1400.770 102.920 1401.090 102.980 ;
        RECT 628.890 102.780 1401.090 102.920 ;
        RECT 628.890 102.720 629.210 102.780 ;
        RECT 1400.770 102.720 1401.090 102.780 ;
      LAYER via ;
        RECT 628.920 102.720 629.180 102.980 ;
        RECT 1400.800 102.720 1401.060 102.980 ;
      LAYER met2 ;
        RECT 630.650 400.250 630.930 404.000 ;
        RECT 629.440 400.110 630.930 400.250 ;
        RECT 629.440 351.970 629.580 400.110 ;
        RECT 630.650 400.000 630.930 400.110 ;
        RECT 628.980 351.830 629.580 351.970 ;
        RECT 628.980 103.010 629.120 351.830 ;
        RECT 628.920 102.690 629.180 103.010 ;
        RECT 1400.800 102.690 1401.060 103.010 ;
        RECT 1400.860 82.870 1401.000 102.690 ;
        RECT 1400.860 82.730 1403.760 82.870 ;
        RECT 1403.620 2.400 1403.760 82.730 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 636.250 102.580 636.570 102.640 ;
        RECT 1421.470 102.580 1421.790 102.640 ;
        RECT 636.250 102.440 1421.790 102.580 ;
        RECT 636.250 102.380 636.570 102.440 ;
        RECT 1421.470 102.380 1421.790 102.440 ;
      LAYER via ;
        RECT 636.280 102.380 636.540 102.640 ;
        RECT 1421.500 102.380 1421.760 102.640 ;
      LAYER met2 ;
        RECT 635.710 400.180 635.990 404.000 ;
        RECT 635.710 400.000 636.020 400.180 ;
        RECT 635.880 376.450 636.020 400.000 ;
        RECT 635.880 376.310 636.480 376.450 ;
        RECT 636.340 102.670 636.480 376.310 ;
        RECT 636.280 102.350 636.540 102.670 ;
        RECT 1421.500 102.350 1421.760 102.670 ;
        RECT 1421.560 2.400 1421.700 102.350 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 635.790 375.940 636.110 376.000 ;
        RECT 639.930 375.940 640.250 376.000 ;
        RECT 635.790 375.800 640.250 375.940 ;
        RECT 635.790 375.740 636.110 375.800 ;
        RECT 639.930 375.740 640.250 375.800 ;
        RECT 635.790 102.240 636.110 102.300 ;
        RECT 1435.270 102.240 1435.590 102.300 ;
        RECT 635.790 102.100 1435.590 102.240 ;
        RECT 635.790 102.040 636.110 102.100 ;
        RECT 1435.270 102.040 1435.590 102.100 ;
      LAYER via ;
        RECT 635.820 375.740 636.080 376.000 ;
        RECT 639.960 375.740 640.220 376.000 ;
        RECT 635.820 102.040 636.080 102.300 ;
        RECT 1435.300 102.040 1435.560 102.300 ;
      LAYER met2 ;
        RECT 641.230 400.250 641.510 404.000 ;
        RECT 640.020 400.110 641.510 400.250 ;
        RECT 640.020 376.030 640.160 400.110 ;
        RECT 641.230 400.000 641.510 400.110 ;
        RECT 635.820 375.710 636.080 376.030 ;
        RECT 639.960 375.710 640.220 376.030 ;
        RECT 635.880 102.330 636.020 375.710 ;
        RECT 635.820 102.010 636.080 102.330 ;
        RECT 1435.300 102.010 1435.560 102.330 ;
        RECT 1435.360 82.870 1435.500 102.010 ;
        RECT 1435.360 82.730 1436.880 82.870 ;
        RECT 1436.740 1.770 1436.880 82.730 ;
        RECT 1438.830 1.770 1439.390 2.400 ;
        RECT 1436.740 1.630 1439.390 1.770 ;
        RECT 1438.830 -4.800 1439.390 1.630 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 642.690 101.900 643.010 101.960 ;
        RECT 1455.970 101.900 1456.290 101.960 ;
        RECT 642.690 101.760 1456.290 101.900 ;
        RECT 642.690 101.700 643.010 101.760 ;
        RECT 1455.970 101.700 1456.290 101.760 ;
      LAYER via ;
        RECT 642.720 101.700 642.980 101.960 ;
        RECT 1456.000 101.700 1456.260 101.960 ;
      LAYER met2 ;
        RECT 646.750 400.250 647.030 404.000 ;
        RECT 645.540 400.110 647.030 400.250 ;
        RECT 645.540 324.370 645.680 400.110 ;
        RECT 646.750 400.000 647.030 400.110 ;
        RECT 642.780 324.230 645.680 324.370 ;
        RECT 642.780 101.990 642.920 324.230 ;
        RECT 642.720 101.670 642.980 101.990 ;
        RECT 1456.000 101.670 1456.260 101.990 ;
        RECT 1456.060 82.870 1456.200 101.670 ;
        RECT 1456.060 82.730 1457.120 82.870 ;
        RECT 1456.980 2.400 1457.120 82.730 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 650.050 101.560 650.370 101.620 ;
        RECT 1469.770 101.560 1470.090 101.620 ;
        RECT 650.050 101.420 1470.090 101.560 ;
        RECT 650.050 101.360 650.370 101.420 ;
        RECT 1469.770 101.360 1470.090 101.420 ;
      LAYER via ;
        RECT 650.080 101.360 650.340 101.620 ;
        RECT 1469.800 101.360 1470.060 101.620 ;
      LAYER met2 ;
        RECT 652.270 400.250 652.550 404.000 ;
        RECT 651.060 400.110 652.550 400.250 ;
        RECT 651.060 324.370 651.200 400.110 ;
        RECT 652.270 400.000 652.550 400.110 ;
        RECT 650.140 324.230 651.200 324.370 ;
        RECT 650.140 101.650 650.280 324.230 ;
        RECT 650.080 101.330 650.340 101.650 ;
        RECT 1469.800 101.330 1470.060 101.650 ;
        RECT 1469.860 82.870 1470.000 101.330 ;
        RECT 1469.860 82.730 1474.600 82.870 ;
        RECT 1474.460 2.400 1474.600 82.730 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 656.030 101.220 656.350 101.280 ;
        RECT 1490.470 101.220 1490.790 101.280 ;
        RECT 656.030 101.080 1490.790 101.220 ;
        RECT 656.030 101.020 656.350 101.080 ;
        RECT 1490.470 101.020 1490.790 101.080 ;
      LAYER via ;
        RECT 656.060 101.020 656.320 101.280 ;
        RECT 1490.500 101.020 1490.760 101.280 ;
      LAYER met2 ;
        RECT 657.790 400.250 658.070 404.000 ;
        RECT 656.580 400.110 658.070 400.250 ;
        RECT 656.580 386.650 656.720 400.110 ;
        RECT 657.790 400.000 658.070 400.110 ;
        RECT 656.120 386.510 656.720 386.650 ;
        RECT 656.120 101.310 656.260 386.510 ;
        RECT 656.060 100.990 656.320 101.310 ;
        RECT 1490.500 100.990 1490.760 101.310 ;
        RECT 1490.560 1.770 1490.700 100.990 ;
        RECT 1492.190 1.770 1492.750 2.400 ;
        RECT 1490.560 1.630 1492.750 1.770 ;
        RECT 1492.190 -4.800 1492.750 1.630 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 663.390 387.640 663.710 387.900 ;
        RECT 663.480 386.880 663.620 387.640 ;
        RECT 663.390 386.620 663.710 386.880 ;
        RECT 663.390 100.880 663.710 100.940 ;
        RECT 1504.270 100.880 1504.590 100.940 ;
        RECT 663.390 100.740 1504.590 100.880 ;
        RECT 663.390 100.680 663.710 100.740 ;
        RECT 1504.270 100.680 1504.590 100.740 ;
      LAYER via ;
        RECT 663.420 387.640 663.680 387.900 ;
        RECT 663.420 386.620 663.680 386.880 ;
        RECT 663.420 100.680 663.680 100.940 ;
        RECT 1504.300 100.680 1504.560 100.940 ;
      LAYER met2 ;
        RECT 663.310 400.180 663.590 404.000 ;
        RECT 663.310 400.000 663.620 400.180 ;
        RECT 663.480 387.930 663.620 400.000 ;
        RECT 663.420 387.610 663.680 387.930 ;
        RECT 663.420 386.590 663.680 386.910 ;
        RECT 663.480 100.970 663.620 386.590 ;
        RECT 663.420 100.650 663.680 100.970 ;
        RECT 1504.300 100.650 1504.560 100.970 ;
        RECT 1504.360 82.870 1504.500 100.650 ;
        RECT 1504.360 82.730 1507.720 82.870 ;
        RECT 1507.580 1.770 1507.720 82.730 ;
        RECT 1509.670 1.770 1510.230 2.400 ;
        RECT 1507.580 1.630 1510.230 1.770 ;
        RECT 1509.670 -4.800 1510.230 1.630 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 414.990 386.480 415.310 386.540 ;
        RECT 416.830 386.480 417.150 386.540 ;
        RECT 414.990 386.340 417.150 386.480 ;
        RECT 414.990 386.280 415.310 386.340 ;
        RECT 416.830 386.280 417.150 386.340 ;
        RECT 414.990 32.880 415.310 32.940 ;
        RECT 552.990 32.880 553.310 32.940 ;
        RECT 414.990 32.740 553.310 32.880 ;
        RECT 414.990 32.680 415.310 32.740 ;
        RECT 552.990 32.680 553.310 32.740 ;
        RECT 552.990 16.560 553.310 16.620 ;
        RECT 712.150 16.560 712.470 16.620 ;
        RECT 552.990 16.420 712.470 16.560 ;
        RECT 552.990 16.360 553.310 16.420 ;
        RECT 712.150 16.360 712.470 16.420 ;
      LAYER via ;
        RECT 415.020 386.280 415.280 386.540 ;
        RECT 416.860 386.280 417.120 386.540 ;
        RECT 415.020 32.680 415.280 32.940 ;
        RECT 553.020 32.680 553.280 32.940 ;
        RECT 553.020 16.360 553.280 16.620 ;
        RECT 712.180 16.360 712.440 16.620 ;
      LAYER met2 ;
        RECT 418.130 400.250 418.410 404.000 ;
        RECT 416.920 400.110 418.410 400.250 ;
        RECT 416.920 386.570 417.060 400.110 ;
        RECT 418.130 400.000 418.410 400.110 ;
        RECT 415.020 386.250 415.280 386.570 ;
        RECT 416.860 386.250 417.120 386.570 ;
        RECT 415.080 32.970 415.220 386.250 ;
        RECT 415.020 32.650 415.280 32.970 ;
        RECT 553.020 32.650 553.280 32.970 ;
        RECT 553.080 16.650 553.220 32.650 ;
        RECT 553.020 16.330 553.280 16.650 ;
        RECT 712.180 16.330 712.440 16.650 ;
        RECT 712.240 2.400 712.380 16.330 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 662.930 386.480 663.250 386.540 ;
        RECT 667.530 386.480 667.850 386.540 ;
        RECT 662.930 386.340 667.850 386.480 ;
        RECT 662.930 386.280 663.250 386.340 ;
        RECT 667.530 386.280 667.850 386.340 ;
        RECT 662.930 100.540 663.250 100.600 ;
        RECT 1524.970 100.540 1525.290 100.600 ;
        RECT 662.930 100.400 1525.290 100.540 ;
        RECT 662.930 100.340 663.250 100.400 ;
        RECT 1524.970 100.340 1525.290 100.400 ;
      LAYER via ;
        RECT 662.960 386.280 663.220 386.540 ;
        RECT 667.560 386.280 667.820 386.540 ;
        RECT 662.960 100.340 663.220 100.600 ;
        RECT 1525.000 100.340 1525.260 100.600 ;
      LAYER met2 ;
        RECT 668.370 400.250 668.650 404.000 ;
        RECT 667.620 400.110 668.650 400.250 ;
        RECT 667.620 386.570 667.760 400.110 ;
        RECT 668.370 400.000 668.650 400.110 ;
        RECT 662.960 386.250 663.220 386.570 ;
        RECT 667.560 386.250 667.820 386.570 ;
        RECT 663.020 100.630 663.160 386.250 ;
        RECT 662.960 100.310 663.220 100.630 ;
        RECT 1525.000 100.310 1525.260 100.630 ;
        RECT 1525.060 82.870 1525.200 100.310 ;
        RECT 1525.060 82.730 1527.960 82.870 ;
        RECT 1527.820 2.400 1527.960 82.730 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 670.290 386.480 670.610 386.540 ;
        RECT 672.590 386.480 672.910 386.540 ;
        RECT 670.290 386.340 672.910 386.480 ;
        RECT 670.290 386.280 670.610 386.340 ;
        RECT 672.590 386.280 672.910 386.340 ;
        RECT 670.290 100.200 670.610 100.260 ;
        RECT 1539.230 100.200 1539.550 100.260 ;
        RECT 670.290 100.060 1539.550 100.200 ;
        RECT 670.290 100.000 670.610 100.060 ;
        RECT 1539.230 100.000 1539.550 100.060 ;
        RECT 1539.230 20.980 1539.550 21.040 ;
        RECT 1545.210 20.980 1545.530 21.040 ;
        RECT 1539.230 20.840 1545.530 20.980 ;
        RECT 1539.230 20.780 1539.550 20.840 ;
        RECT 1545.210 20.780 1545.530 20.840 ;
      LAYER via ;
        RECT 670.320 386.280 670.580 386.540 ;
        RECT 672.620 386.280 672.880 386.540 ;
        RECT 670.320 100.000 670.580 100.260 ;
        RECT 1539.260 100.000 1539.520 100.260 ;
        RECT 1539.260 20.780 1539.520 21.040 ;
        RECT 1545.240 20.780 1545.500 21.040 ;
      LAYER met2 ;
        RECT 673.890 400.250 674.170 404.000 ;
        RECT 672.680 400.110 674.170 400.250 ;
        RECT 672.680 386.570 672.820 400.110 ;
        RECT 673.890 400.000 674.170 400.110 ;
        RECT 670.320 386.250 670.580 386.570 ;
        RECT 672.620 386.250 672.880 386.570 ;
        RECT 670.380 100.290 670.520 386.250 ;
        RECT 670.320 99.970 670.580 100.290 ;
        RECT 1539.260 99.970 1539.520 100.290 ;
        RECT 1539.320 21.070 1539.460 99.970 ;
        RECT 1539.260 20.750 1539.520 21.070 ;
        RECT 1545.240 20.750 1545.500 21.070 ;
        RECT 1545.300 2.400 1545.440 20.750 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.730 374.580 677.050 374.640 ;
        RECT 678.110 374.580 678.430 374.640 ;
        RECT 676.730 374.440 678.430 374.580 ;
        RECT 676.730 374.380 677.050 374.440 ;
        RECT 678.110 374.380 678.430 374.440 ;
        RECT 676.730 99.860 677.050 99.920 ;
        RECT 1559.470 99.860 1559.790 99.920 ;
        RECT 676.730 99.720 1559.790 99.860 ;
        RECT 676.730 99.660 677.050 99.720 ;
        RECT 1559.470 99.660 1559.790 99.720 ;
      LAYER via ;
        RECT 676.760 374.380 677.020 374.640 ;
        RECT 678.140 374.380 678.400 374.640 ;
        RECT 676.760 99.660 677.020 99.920 ;
        RECT 1559.500 99.660 1559.760 99.920 ;
      LAYER met2 ;
        RECT 679.410 400.250 679.690 404.000 ;
        RECT 678.200 400.110 679.690 400.250 ;
        RECT 678.200 374.670 678.340 400.110 ;
        RECT 679.410 400.000 679.690 400.110 ;
        RECT 676.760 374.350 677.020 374.670 ;
        RECT 678.140 374.350 678.400 374.670 ;
        RECT 676.820 99.950 676.960 374.350 ;
        RECT 676.760 99.630 677.020 99.950 ;
        RECT 1559.500 99.630 1559.760 99.950 ;
        RECT 1559.560 82.870 1559.700 99.630 ;
        RECT 1559.560 82.730 1561.080 82.870 ;
        RECT 1560.940 1.770 1561.080 82.730 ;
        RECT 1563.030 1.770 1563.590 2.400 ;
        RECT 1560.940 1.630 1563.590 1.770 ;
        RECT 1563.030 -4.800 1563.590 1.630 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.930 400.250 685.210 404.000 ;
        RECT 684.640 400.110 685.210 400.250 ;
        RECT 684.640 99.805 684.780 400.110 ;
        RECT 684.930 400.000 685.210 400.110 ;
        RECT 684.570 99.435 684.850 99.805 ;
        RECT 1580.190 99.435 1580.470 99.805 ;
        RECT 1580.260 82.870 1580.400 99.435 ;
        RECT 1580.260 82.730 1581.320 82.870 ;
        RECT 1581.180 2.400 1581.320 82.730 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
      LAYER via2 ;
        RECT 684.570 99.480 684.850 99.760 ;
        RECT 1580.190 99.480 1580.470 99.760 ;
      LAYER met3 ;
        RECT 684.545 99.770 684.875 99.785 ;
        RECT 1580.165 99.770 1580.495 99.785 ;
        RECT 684.545 99.470 1580.495 99.770 ;
        RECT 684.545 99.455 684.875 99.470 ;
        RECT 1580.165 99.455 1580.495 99.470 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 691.450 126.040 691.770 126.100 ;
        RECT 1593.970 126.040 1594.290 126.100 ;
        RECT 691.450 125.900 1594.290 126.040 ;
        RECT 691.450 125.840 691.770 125.900 ;
        RECT 1593.970 125.840 1594.290 125.900 ;
      LAYER via ;
        RECT 691.480 125.840 691.740 126.100 ;
        RECT 1594.000 125.840 1594.260 126.100 ;
      LAYER met2 ;
        RECT 690.450 400.250 690.730 404.000 ;
        RECT 690.450 400.110 691.680 400.250 ;
        RECT 690.450 400.000 690.730 400.110 ;
        RECT 691.540 126.130 691.680 400.110 ;
        RECT 691.480 125.810 691.740 126.130 ;
        RECT 1594.000 125.810 1594.260 126.130 ;
        RECT 1594.060 82.870 1594.200 125.810 ;
        RECT 1594.060 82.730 1598.800 82.870 ;
        RECT 1598.660 2.400 1598.800 82.730 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 690.990 386.140 691.310 386.200 ;
        RECT 694.670 386.140 694.990 386.200 ;
        RECT 690.990 386.000 694.990 386.140 ;
        RECT 690.990 385.940 691.310 386.000 ;
        RECT 694.670 385.940 694.990 386.000 ;
        RECT 690.990 126.380 691.310 126.440 ;
        RECT 1614.670 126.380 1614.990 126.440 ;
        RECT 690.990 126.240 1614.990 126.380 ;
        RECT 690.990 126.180 691.310 126.240 ;
        RECT 1614.670 126.180 1614.990 126.240 ;
      LAYER via ;
        RECT 691.020 385.940 691.280 386.200 ;
        RECT 694.700 385.940 694.960 386.200 ;
        RECT 691.020 126.180 691.280 126.440 ;
        RECT 1614.700 126.180 1614.960 126.440 ;
      LAYER met2 ;
        RECT 695.970 400.250 696.250 404.000 ;
        RECT 694.760 400.110 696.250 400.250 ;
        RECT 694.760 386.230 694.900 400.110 ;
        RECT 695.970 400.000 696.250 400.110 ;
        RECT 691.020 385.910 691.280 386.230 ;
        RECT 694.700 385.910 694.960 386.230 ;
        RECT 691.080 126.470 691.220 385.910 ;
        RECT 691.020 126.150 691.280 126.470 ;
        RECT 1614.700 126.150 1614.960 126.470 ;
        RECT 1614.760 1.770 1614.900 126.150 ;
        RECT 1616.390 1.770 1616.950 2.400 ;
        RECT 1614.760 1.630 1616.950 1.770 ;
        RECT 1616.390 -4.800 1616.950 1.630 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 698.350 126.720 698.670 126.780 ;
        RECT 1628.470 126.720 1628.790 126.780 ;
        RECT 698.350 126.580 1628.790 126.720 ;
        RECT 698.350 126.520 698.670 126.580 ;
        RECT 1628.470 126.520 1628.790 126.580 ;
      LAYER via ;
        RECT 698.380 126.520 698.640 126.780 ;
        RECT 1628.500 126.520 1628.760 126.780 ;
      LAYER met2 ;
        RECT 701.030 400.250 701.310 404.000 ;
        RECT 700.280 400.110 701.310 400.250 ;
        RECT 700.280 324.370 700.420 400.110 ;
        RECT 701.030 400.000 701.310 400.110 ;
        RECT 698.440 324.230 700.420 324.370 ;
        RECT 698.440 126.810 698.580 324.230 ;
        RECT 698.380 126.490 698.640 126.810 ;
        RECT 1628.500 126.490 1628.760 126.810 ;
        RECT 1628.560 82.870 1628.700 126.490 ;
        RECT 1628.560 82.730 1631.920 82.870 ;
        RECT 1631.780 1.770 1631.920 82.730 ;
        RECT 1633.870 1.770 1634.430 2.400 ;
        RECT 1631.780 1.630 1634.430 1.770 ;
        RECT 1633.870 -4.800 1634.430 1.630 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 705.250 127.060 705.570 127.120 ;
        RECT 1649.170 127.060 1649.490 127.120 ;
        RECT 705.250 126.920 1649.490 127.060 ;
        RECT 705.250 126.860 705.570 126.920 ;
        RECT 1649.170 126.860 1649.490 126.920 ;
      LAYER via ;
        RECT 705.280 126.860 705.540 127.120 ;
        RECT 1649.200 126.860 1649.460 127.120 ;
      LAYER met2 ;
        RECT 706.550 400.250 706.830 404.000 ;
        RECT 705.340 400.110 706.830 400.250 ;
        RECT 705.340 127.150 705.480 400.110 ;
        RECT 706.550 400.000 706.830 400.110 ;
        RECT 705.280 126.830 705.540 127.150 ;
        RECT 1649.200 126.830 1649.460 127.150 ;
        RECT 1649.260 82.870 1649.400 126.830 ;
        RECT 1649.260 82.730 1652.160 82.870 ;
        RECT 1652.020 2.400 1652.160 82.730 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 711.690 127.400 712.010 127.460 ;
        RECT 1662.970 127.400 1663.290 127.460 ;
        RECT 711.690 127.260 1663.290 127.400 ;
        RECT 711.690 127.200 712.010 127.260 ;
        RECT 1662.970 127.200 1663.290 127.260 ;
        RECT 1662.970 15.200 1663.290 15.260 ;
        RECT 1669.410 15.200 1669.730 15.260 ;
        RECT 1662.970 15.060 1669.730 15.200 ;
        RECT 1662.970 15.000 1663.290 15.060 ;
        RECT 1669.410 15.000 1669.730 15.060 ;
      LAYER via ;
        RECT 711.720 127.200 711.980 127.460 ;
        RECT 1663.000 127.200 1663.260 127.460 ;
        RECT 1663.000 15.000 1663.260 15.260 ;
        RECT 1669.440 15.000 1669.700 15.260 ;
      LAYER met2 ;
        RECT 712.070 400.250 712.350 404.000 ;
        RECT 711.780 400.110 712.350 400.250 ;
        RECT 711.780 127.490 711.920 400.110 ;
        RECT 712.070 400.000 712.350 400.110 ;
        RECT 711.720 127.170 711.980 127.490 ;
        RECT 1663.000 127.170 1663.260 127.490 ;
        RECT 1663.060 15.290 1663.200 127.170 ;
        RECT 1663.000 14.970 1663.260 15.290 ;
        RECT 1669.440 14.970 1669.700 15.290 ;
        RECT 1669.500 2.400 1669.640 14.970 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 719.050 131.140 719.370 131.200 ;
        RECT 1683.670 131.140 1683.990 131.200 ;
        RECT 719.050 131.000 1683.990 131.140 ;
        RECT 719.050 130.940 719.370 131.000 ;
        RECT 1683.670 130.940 1683.990 131.000 ;
      LAYER via ;
        RECT 719.080 130.940 719.340 131.200 ;
        RECT 1683.700 130.940 1683.960 131.200 ;
      LAYER met2 ;
        RECT 717.590 400.930 717.870 404.000 ;
        RECT 717.590 400.790 719.280 400.930 ;
        RECT 717.590 400.000 717.870 400.790 ;
        RECT 719.140 131.230 719.280 400.790 ;
        RECT 719.080 130.910 719.340 131.230 ;
        RECT 1683.700 130.910 1683.960 131.230 ;
        RECT 1683.760 82.870 1683.900 130.910 ;
        RECT 1683.760 82.730 1685.280 82.870 ;
        RECT 1685.140 1.770 1685.280 82.730 ;
        RECT 1687.230 1.770 1687.790 2.400 ;
        RECT 1685.140 1.630 1687.790 1.770 ;
        RECT 1687.230 -4.800 1687.790 1.630 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 421.430 386.480 421.750 386.540 ;
        RECT 422.350 386.480 422.670 386.540 ;
        RECT 421.430 386.340 422.670 386.480 ;
        RECT 421.430 386.280 421.750 386.340 ;
        RECT 422.350 386.280 422.670 386.340 ;
        RECT 421.430 33.220 421.750 33.280 ;
        RECT 558.510 33.220 558.830 33.280 ;
        RECT 421.430 33.080 558.830 33.220 ;
        RECT 421.430 33.020 421.750 33.080 ;
        RECT 558.510 33.020 558.830 33.080 ;
        RECT 558.510 20.640 558.830 20.700 ;
        RECT 729.630 20.640 729.950 20.700 ;
        RECT 558.510 20.500 729.950 20.640 ;
        RECT 558.510 20.440 558.830 20.500 ;
        RECT 729.630 20.440 729.950 20.500 ;
      LAYER via ;
        RECT 421.460 386.280 421.720 386.540 ;
        RECT 422.380 386.280 422.640 386.540 ;
        RECT 421.460 33.020 421.720 33.280 ;
        RECT 558.540 33.020 558.800 33.280 ;
        RECT 558.540 20.440 558.800 20.700 ;
        RECT 729.660 20.440 729.920 20.700 ;
      LAYER met2 ;
        RECT 423.650 400.250 423.930 404.000 ;
        RECT 422.440 400.110 423.930 400.250 ;
        RECT 422.440 386.570 422.580 400.110 ;
        RECT 423.650 400.000 423.930 400.110 ;
        RECT 421.460 386.250 421.720 386.570 ;
        RECT 422.380 386.250 422.640 386.570 ;
        RECT 421.520 33.310 421.660 386.250 ;
        RECT 421.460 32.990 421.720 33.310 ;
        RECT 558.540 32.990 558.800 33.310 ;
        RECT 558.600 20.730 558.740 32.990 ;
        RECT 558.540 20.410 558.800 20.730 ;
        RECT 729.660 20.410 729.920 20.730 ;
        RECT 729.720 2.400 729.860 20.410 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 718.590 386.480 718.910 386.540 ;
        RECT 721.810 386.480 722.130 386.540 ;
        RECT 718.590 386.340 722.130 386.480 ;
        RECT 718.590 386.280 718.910 386.340 ;
        RECT 721.810 386.280 722.130 386.340 ;
        RECT 718.590 130.800 718.910 130.860 ;
        RECT 1704.370 130.800 1704.690 130.860 ;
        RECT 718.590 130.660 1704.690 130.800 ;
        RECT 718.590 130.600 718.910 130.660 ;
        RECT 1704.370 130.600 1704.690 130.660 ;
      LAYER via ;
        RECT 718.620 386.280 718.880 386.540 ;
        RECT 721.840 386.280 722.100 386.540 ;
        RECT 718.620 130.600 718.880 130.860 ;
        RECT 1704.400 130.600 1704.660 130.860 ;
      LAYER met2 ;
        RECT 723.110 400.250 723.390 404.000 ;
        RECT 721.900 400.110 723.390 400.250 ;
        RECT 721.900 386.570 722.040 400.110 ;
        RECT 723.110 400.000 723.390 400.110 ;
        RECT 718.620 386.250 718.880 386.570 ;
        RECT 721.840 386.250 722.100 386.570 ;
        RECT 718.680 130.890 718.820 386.250 ;
        RECT 718.620 130.570 718.880 130.890 ;
        RECT 1704.400 130.570 1704.660 130.890 ;
        RECT 1704.460 82.870 1704.600 130.570 ;
        RECT 1704.460 82.730 1705.060 82.870 ;
        RECT 1704.920 2.400 1705.060 82.730 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 725.950 130.460 726.270 130.520 ;
        RECT 1718.170 130.460 1718.490 130.520 ;
        RECT 725.950 130.320 1718.490 130.460 ;
        RECT 725.950 130.260 726.270 130.320 ;
        RECT 1718.170 130.260 1718.490 130.320 ;
      LAYER via ;
        RECT 725.980 130.260 726.240 130.520 ;
        RECT 1718.200 130.260 1718.460 130.520 ;
      LAYER met2 ;
        RECT 728.630 400.250 728.910 404.000 ;
        RECT 727.420 400.110 728.910 400.250 ;
        RECT 727.420 324.370 727.560 400.110 ;
        RECT 728.630 400.000 728.910 400.110 ;
        RECT 726.040 324.230 727.560 324.370 ;
        RECT 726.040 130.550 726.180 324.230 ;
        RECT 725.980 130.230 726.240 130.550 ;
        RECT 1718.200 130.230 1718.460 130.550 ;
        RECT 1718.260 82.870 1718.400 130.230 ;
        RECT 1718.260 82.730 1723.000 82.870 ;
        RECT 1722.860 2.400 1723.000 82.730 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 732.850 130.120 733.170 130.180 ;
        RECT 1738.870 130.120 1739.190 130.180 ;
        RECT 732.850 129.980 1739.190 130.120 ;
        RECT 732.850 129.920 733.170 129.980 ;
        RECT 1738.870 129.920 1739.190 129.980 ;
      LAYER via ;
        RECT 732.880 129.920 733.140 130.180 ;
        RECT 1738.900 129.920 1739.160 130.180 ;
      LAYER met2 ;
        RECT 733.690 400.250 733.970 404.000 ;
        RECT 732.940 400.110 733.970 400.250 ;
        RECT 732.940 130.210 733.080 400.110 ;
        RECT 733.690 400.000 733.970 400.110 ;
        RECT 732.880 129.890 733.140 130.210 ;
        RECT 1738.900 129.890 1739.160 130.210 ;
        RECT 1738.960 82.870 1739.100 129.890 ;
        RECT 1738.960 82.730 1740.480 82.870 ;
        RECT 1740.340 2.400 1740.480 82.730 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 739.290 129.780 739.610 129.840 ;
        RECT 1752.670 129.780 1752.990 129.840 ;
        RECT 739.290 129.640 1752.990 129.780 ;
        RECT 739.290 129.580 739.610 129.640 ;
        RECT 1752.670 129.580 1752.990 129.640 ;
      LAYER via ;
        RECT 739.320 129.580 739.580 129.840 ;
        RECT 1752.700 129.580 1752.960 129.840 ;
      LAYER met2 ;
        RECT 739.210 400.180 739.490 404.000 ;
        RECT 739.210 400.000 739.520 400.180 ;
        RECT 739.380 129.870 739.520 400.000 ;
        RECT 739.320 129.550 739.580 129.870 ;
        RECT 1752.700 129.550 1752.960 129.870 ;
        RECT 1752.760 82.870 1752.900 129.550 ;
        RECT 1752.760 82.730 1756.120 82.870 ;
        RECT 1755.980 1.770 1756.120 82.730 ;
        RECT 1758.070 1.770 1758.630 2.400 ;
        RECT 1755.980 1.630 1758.630 1.770 ;
        RECT 1758.070 -4.800 1758.630 1.630 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 739.750 129.440 740.070 129.500 ;
        RECT 1773.370 129.440 1773.690 129.500 ;
        RECT 739.750 129.300 1773.690 129.440 ;
        RECT 739.750 129.240 740.070 129.300 ;
        RECT 1773.370 129.240 1773.690 129.300 ;
      LAYER via ;
        RECT 739.780 129.240 740.040 129.500 ;
        RECT 1773.400 129.240 1773.660 129.500 ;
      LAYER met2 ;
        RECT 744.730 400.250 745.010 404.000 ;
        RECT 743.520 400.110 745.010 400.250 ;
        RECT 743.520 324.370 743.660 400.110 ;
        RECT 744.730 400.000 745.010 400.110 ;
        RECT 739.840 324.230 743.660 324.370 ;
        RECT 739.840 129.530 739.980 324.230 ;
        RECT 739.780 129.210 740.040 129.530 ;
        RECT 1773.400 129.210 1773.660 129.530 ;
        RECT 1773.460 82.870 1773.600 129.210 ;
        RECT 1773.460 82.730 1776.360 82.870 ;
        RECT 1776.220 2.400 1776.360 82.730 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 746.190 129.100 746.510 129.160 ;
        RECT 1787.170 129.100 1787.490 129.160 ;
        RECT 746.190 128.960 1787.490 129.100 ;
        RECT 746.190 128.900 746.510 128.960 ;
        RECT 1787.170 128.900 1787.490 128.960 ;
        RECT 1787.170 15.200 1787.490 15.260 ;
        RECT 1793.610 15.200 1793.930 15.260 ;
        RECT 1787.170 15.060 1793.930 15.200 ;
        RECT 1787.170 15.000 1787.490 15.060 ;
        RECT 1793.610 15.000 1793.930 15.060 ;
      LAYER via ;
        RECT 746.220 128.900 746.480 129.160 ;
        RECT 1787.200 128.900 1787.460 129.160 ;
        RECT 1787.200 15.000 1787.460 15.260 ;
        RECT 1793.640 15.000 1793.900 15.260 ;
      LAYER met2 ;
        RECT 750.250 400.250 750.530 404.000 ;
        RECT 749.040 400.110 750.530 400.250 ;
        RECT 749.040 386.480 749.180 400.110 ;
        RECT 750.250 400.000 750.530 400.110 ;
        RECT 746.280 386.340 749.180 386.480 ;
        RECT 746.280 129.190 746.420 386.340 ;
        RECT 746.220 128.870 746.480 129.190 ;
        RECT 1787.200 128.870 1787.460 129.190 ;
        RECT 1787.260 15.290 1787.400 128.870 ;
        RECT 1787.200 14.970 1787.460 15.290 ;
        RECT 1793.640 14.970 1793.900 15.290 ;
        RECT 1793.700 2.400 1793.840 14.970 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 755.850 393.280 756.170 393.340 ;
        RECT 1807.870 393.280 1808.190 393.340 ;
        RECT 755.850 393.140 1808.190 393.280 ;
        RECT 755.850 393.080 756.170 393.140 ;
        RECT 1807.870 393.080 1808.190 393.140 ;
      LAYER via ;
        RECT 755.880 393.080 756.140 393.340 ;
        RECT 1807.900 393.080 1808.160 393.340 ;
      LAYER met2 ;
        RECT 755.770 400.180 756.050 404.000 ;
        RECT 755.770 400.000 756.080 400.180 ;
        RECT 755.940 393.370 756.080 400.000 ;
        RECT 755.880 393.050 756.140 393.370 ;
        RECT 1807.900 393.050 1808.160 393.370 ;
        RECT 1807.960 82.870 1808.100 393.050 ;
        RECT 1807.960 82.730 1809.480 82.870 ;
        RECT 1809.340 1.770 1809.480 82.730 ;
        RECT 1811.430 1.770 1811.990 2.400 ;
        RECT 1809.340 1.630 1811.990 1.770 ;
        RECT 1811.430 -4.800 1811.990 1.630 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 760.450 128.760 760.770 128.820 ;
        RECT 1828.570 128.760 1828.890 128.820 ;
        RECT 760.450 128.620 1828.890 128.760 ;
        RECT 760.450 128.560 760.770 128.620 ;
        RECT 1828.570 128.560 1828.890 128.620 ;
      LAYER via ;
        RECT 760.480 128.560 760.740 128.820 ;
        RECT 1828.600 128.560 1828.860 128.820 ;
      LAYER met2 ;
        RECT 761.290 400.250 761.570 404.000 ;
        RECT 760.540 400.110 761.570 400.250 ;
        RECT 760.540 128.850 760.680 400.110 ;
        RECT 761.290 400.000 761.570 400.110 ;
        RECT 760.480 128.530 760.740 128.850 ;
        RECT 1828.600 128.530 1828.860 128.850 ;
        RECT 1828.660 82.870 1828.800 128.530 ;
        RECT 1828.660 82.730 1829.260 82.870 ;
        RECT 1829.120 2.400 1829.260 82.730 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.890 392.940 767.210 393.000 ;
        RECT 1842.370 392.940 1842.690 393.000 ;
        RECT 766.890 392.800 1842.690 392.940 ;
        RECT 766.890 392.740 767.210 392.800 ;
        RECT 1842.370 392.740 1842.690 392.800 ;
      LAYER via ;
        RECT 766.920 392.740 767.180 393.000 ;
        RECT 1842.400 392.740 1842.660 393.000 ;
      LAYER met2 ;
        RECT 766.810 400.180 767.090 404.000 ;
        RECT 766.810 400.000 767.120 400.180 ;
        RECT 766.980 393.030 767.120 400.000 ;
        RECT 766.920 392.710 767.180 393.030 ;
        RECT 1842.400 392.710 1842.660 393.030 ;
        RECT 1842.460 82.870 1842.600 392.710 ;
        RECT 1842.460 82.730 1847.200 82.870 ;
        RECT 1847.060 2.400 1847.200 82.730 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 766.890 385.460 767.210 385.520 ;
        RECT 770.570 385.460 770.890 385.520 ;
        RECT 766.890 385.320 770.890 385.460 ;
        RECT 766.890 385.260 767.210 385.320 ;
        RECT 770.570 385.260 770.890 385.320 ;
        RECT 766.890 128.420 767.210 128.480 ;
        RECT 1863.070 128.420 1863.390 128.480 ;
        RECT 766.890 128.280 1863.390 128.420 ;
        RECT 766.890 128.220 767.210 128.280 ;
        RECT 1863.070 128.220 1863.390 128.280 ;
      LAYER via ;
        RECT 766.920 385.260 767.180 385.520 ;
        RECT 770.600 385.260 770.860 385.520 ;
        RECT 766.920 128.220 767.180 128.480 ;
        RECT 1863.100 128.220 1863.360 128.480 ;
      LAYER met2 ;
        RECT 771.870 400.250 772.150 404.000 ;
        RECT 770.660 400.110 772.150 400.250 ;
        RECT 770.660 385.550 770.800 400.110 ;
        RECT 771.870 400.000 772.150 400.110 ;
        RECT 766.920 385.230 767.180 385.550 ;
        RECT 770.600 385.230 770.860 385.550 ;
        RECT 766.980 128.510 767.120 385.230 ;
        RECT 766.920 128.190 767.180 128.510 ;
        RECT 1863.100 128.190 1863.360 128.510 ;
        RECT 1863.160 82.870 1863.300 128.190 ;
        RECT 1863.160 82.730 1864.680 82.870 ;
        RECT 1864.540 2.400 1864.680 82.730 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 428.330 22.000 428.650 22.060 ;
        RECT 503.770 22.000 504.090 22.060 ;
        RECT 428.330 21.860 504.090 22.000 ;
        RECT 428.330 21.800 428.650 21.860 ;
        RECT 503.770 21.800 504.090 21.860 ;
        RECT 503.770 18.260 504.090 18.320 ;
        RECT 747.570 18.260 747.890 18.320 ;
        RECT 503.770 18.120 747.890 18.260 ;
        RECT 503.770 18.060 504.090 18.120 ;
        RECT 747.570 18.060 747.890 18.120 ;
      LAYER via ;
        RECT 428.360 21.800 428.620 22.060 ;
        RECT 503.800 21.800 504.060 22.060 ;
        RECT 503.800 18.060 504.060 18.320 ;
        RECT 747.600 18.060 747.860 18.320 ;
      LAYER met2 ;
        RECT 429.170 400.250 429.450 404.000 ;
        RECT 428.420 400.110 429.450 400.250 ;
        RECT 428.420 22.090 428.560 400.110 ;
        RECT 429.170 400.000 429.450 400.110 ;
        RECT 428.360 21.770 428.620 22.090 ;
        RECT 503.800 21.770 504.060 22.090 ;
        RECT 503.860 18.350 504.000 21.770 ;
        RECT 503.800 18.030 504.060 18.350 ;
        RECT 747.600 18.030 747.860 18.350 ;
        RECT 747.660 2.400 747.800 18.030 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1876.870 392.600 1877.190 392.660 ;
        RECT 786.530 392.460 1877.190 392.600 ;
        RECT 777.470 391.920 777.790 391.980 ;
        RECT 786.530 391.920 786.670 392.460 ;
        RECT 1876.870 392.400 1877.190 392.460 ;
        RECT 777.470 391.780 786.670 391.920 ;
        RECT 777.470 391.720 777.790 391.780 ;
      LAYER via ;
        RECT 777.500 391.720 777.760 391.980 ;
        RECT 1876.900 392.400 1877.160 392.660 ;
      LAYER met2 ;
        RECT 777.390 400.180 777.670 404.000 ;
        RECT 777.390 400.000 777.700 400.180 ;
        RECT 777.560 392.010 777.700 400.000 ;
        RECT 1876.900 392.370 1877.160 392.690 ;
        RECT 777.500 391.690 777.760 392.010 ;
        RECT 1876.960 82.870 1877.100 392.370 ;
        RECT 1876.960 82.730 1880.320 82.870 ;
        RECT 1880.180 1.770 1880.320 82.730 ;
        RECT 1882.270 1.770 1882.830 2.400 ;
        RECT 1880.180 1.630 1882.830 1.770 ;
        RECT 1882.270 -4.800 1882.830 1.630 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 780.690 128.080 781.010 128.140 ;
        RECT 1897.570 128.080 1897.890 128.140 ;
        RECT 780.690 127.940 1897.890 128.080 ;
        RECT 780.690 127.880 781.010 127.940 ;
        RECT 1897.570 127.880 1897.890 127.940 ;
      LAYER via ;
        RECT 780.720 127.880 780.980 128.140 ;
        RECT 1897.600 127.880 1897.860 128.140 ;
      LAYER met2 ;
        RECT 782.910 400.250 783.190 404.000 ;
        RECT 781.700 400.110 783.190 400.250 ;
        RECT 781.700 324.370 781.840 400.110 ;
        RECT 782.910 400.000 783.190 400.110 ;
        RECT 780.780 324.230 781.840 324.370 ;
        RECT 780.780 128.170 780.920 324.230 ;
        RECT 780.720 127.850 780.980 128.170 ;
        RECT 1897.600 127.850 1897.860 128.170 ;
        RECT 1897.660 1.770 1897.800 127.850 ;
        RECT 1899.750 1.770 1900.310 2.400 ;
        RECT 1897.660 1.630 1900.310 1.770 ;
        RECT 1899.750 -4.800 1900.310 1.630 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 788.510 392.260 788.830 392.320 ;
        RECT 1911.370 392.260 1911.690 392.320 ;
        RECT 788.510 392.120 1911.690 392.260 ;
        RECT 788.510 392.060 788.830 392.120 ;
        RECT 1911.370 392.060 1911.690 392.120 ;
        RECT 1911.370 15.200 1911.690 15.260 ;
        RECT 1917.810 15.200 1918.130 15.260 ;
        RECT 1911.370 15.060 1918.130 15.200 ;
        RECT 1911.370 15.000 1911.690 15.060 ;
        RECT 1917.810 15.000 1918.130 15.060 ;
      LAYER via ;
        RECT 788.540 392.060 788.800 392.320 ;
        RECT 1911.400 392.060 1911.660 392.320 ;
        RECT 1911.400 15.000 1911.660 15.260 ;
        RECT 1917.840 15.000 1918.100 15.260 ;
      LAYER met2 ;
        RECT 788.430 400.180 788.710 404.000 ;
        RECT 788.430 400.000 788.740 400.180 ;
        RECT 788.600 392.350 788.740 400.000 ;
        RECT 788.540 392.030 788.800 392.350 ;
        RECT 1911.400 392.030 1911.660 392.350 ;
        RECT 1911.460 15.290 1911.600 392.030 ;
        RECT 1911.400 14.970 1911.660 15.290 ;
        RECT 1917.840 14.970 1918.100 15.290 ;
        RECT 1917.900 2.400 1918.040 14.970 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 794.490 127.740 794.810 127.800 ;
        RECT 1932.070 127.740 1932.390 127.800 ;
        RECT 794.490 127.600 1932.390 127.740 ;
        RECT 794.490 127.540 794.810 127.600 ;
        RECT 1932.070 127.540 1932.390 127.600 ;
      LAYER via ;
        RECT 794.520 127.540 794.780 127.800 ;
        RECT 1932.100 127.540 1932.360 127.800 ;
      LAYER met2 ;
        RECT 793.950 400.250 794.230 404.000 ;
        RECT 793.660 400.110 794.230 400.250 ;
        RECT 793.660 398.890 793.800 400.110 ;
        RECT 793.950 400.000 794.230 400.110 ;
        RECT 793.660 398.750 794.260 398.890 ;
        RECT 794.120 377.130 794.260 398.750 ;
        RECT 794.120 376.990 794.720 377.130 ;
        RECT 794.580 127.830 794.720 376.990 ;
        RECT 794.520 127.510 794.780 127.830 ;
        RECT 1932.100 127.510 1932.360 127.830 ;
        RECT 1932.160 82.870 1932.300 127.510 ;
        RECT 1932.160 82.730 1933.680 82.870 ;
        RECT 1933.540 1.770 1933.680 82.730 ;
        RECT 1935.630 1.770 1936.190 2.400 ;
        RECT 1933.540 1.630 1936.190 1.770 ;
        RECT 1935.630 -4.800 1936.190 1.630 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 799.550 391.580 799.870 391.640 ;
        RECT 1952.770 391.580 1953.090 391.640 ;
        RECT 799.550 391.440 1953.090 391.580 ;
        RECT 799.550 391.380 799.870 391.440 ;
        RECT 1952.770 391.380 1953.090 391.440 ;
      LAYER via ;
        RECT 799.580 391.380 799.840 391.640 ;
        RECT 1952.800 391.380 1953.060 391.640 ;
      LAYER met2 ;
        RECT 799.470 400.180 799.750 404.000 ;
        RECT 799.470 400.000 799.780 400.180 ;
        RECT 799.640 391.670 799.780 400.000 ;
        RECT 799.580 391.350 799.840 391.670 ;
        RECT 1952.800 391.350 1953.060 391.670 ;
        RECT 1952.860 82.870 1953.000 391.350 ;
        RECT 1952.860 82.730 1953.460 82.870 ;
        RECT 1953.320 2.400 1953.460 82.730 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.530 400.250 804.810 404.000 ;
        RECT 803.320 400.110 804.810 400.250 ;
        RECT 803.320 324.370 803.460 400.110 ;
        RECT 804.530 400.000 804.810 400.110 ;
        RECT 801.940 324.230 803.460 324.370 ;
        RECT 801.940 127.685 802.080 324.230 ;
        RECT 801.870 127.315 802.150 127.685 ;
        RECT 1966.590 127.315 1966.870 127.685 ;
        RECT 1966.660 82.870 1966.800 127.315 ;
        RECT 1966.660 82.730 1971.400 82.870 ;
        RECT 1971.260 2.400 1971.400 82.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
      LAYER via2 ;
        RECT 801.870 127.360 802.150 127.640 ;
        RECT 1966.590 127.360 1966.870 127.640 ;
      LAYER met3 ;
        RECT 801.845 127.650 802.175 127.665 ;
        RECT 1966.565 127.650 1966.895 127.665 ;
        RECT 801.845 127.350 1966.895 127.650 ;
        RECT 801.845 127.335 802.175 127.350 ;
        RECT 1966.565 127.335 1966.895 127.350 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 810.130 391.240 810.450 391.300 ;
        RECT 1987.270 391.240 1987.590 391.300 ;
        RECT 810.130 391.100 1987.590 391.240 ;
        RECT 810.130 391.040 810.450 391.100 ;
        RECT 1987.270 391.040 1987.590 391.100 ;
      LAYER via ;
        RECT 810.160 391.040 810.420 391.300 ;
        RECT 1987.300 391.040 1987.560 391.300 ;
      LAYER met2 ;
        RECT 810.050 400.180 810.330 404.000 ;
        RECT 810.050 400.000 810.360 400.180 ;
        RECT 810.220 391.330 810.360 400.000 ;
        RECT 810.160 391.010 810.420 391.330 ;
        RECT 1987.300 391.010 1987.560 391.330 ;
        RECT 1987.360 82.870 1987.500 391.010 ;
        RECT 1987.360 82.730 1988.880 82.870 ;
        RECT 1988.740 2.400 1988.880 82.730 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 815.190 135.560 815.510 135.620 ;
        RECT 2001.070 135.560 2001.390 135.620 ;
        RECT 815.190 135.420 2001.390 135.560 ;
        RECT 815.190 135.360 815.510 135.420 ;
        RECT 2001.070 135.360 2001.390 135.420 ;
      LAYER via ;
        RECT 815.220 135.360 815.480 135.620 ;
        RECT 2001.100 135.360 2001.360 135.620 ;
      LAYER met2 ;
        RECT 815.570 400.180 815.850 404.000 ;
        RECT 815.570 400.000 815.880 400.180 ;
        RECT 815.740 324.370 815.880 400.000 ;
        RECT 815.280 324.230 815.880 324.370 ;
        RECT 815.280 135.650 815.420 324.230 ;
        RECT 815.220 135.330 815.480 135.650 ;
        RECT 2001.100 135.330 2001.360 135.650 ;
        RECT 2001.160 82.870 2001.300 135.330 ;
        RECT 2001.160 82.730 2004.520 82.870 ;
        RECT 2004.380 1.770 2004.520 82.730 ;
        RECT 2006.470 1.770 2007.030 2.400 ;
        RECT 2004.380 1.630 2007.030 1.770 ;
        RECT 2006.470 -4.800 2007.030 1.630 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 822.090 390.900 822.410 390.960 ;
        RECT 2021.770 390.900 2022.090 390.960 ;
        RECT 822.090 390.760 2022.090 390.900 ;
        RECT 822.090 390.700 822.410 390.760 ;
        RECT 2021.770 390.700 2022.090 390.760 ;
      LAYER via ;
        RECT 822.120 390.700 822.380 390.960 ;
        RECT 2021.800 390.700 2022.060 390.960 ;
      LAYER met2 ;
        RECT 821.090 400.250 821.370 404.000 ;
        RECT 821.090 400.110 822.320 400.250 ;
        RECT 821.090 400.000 821.370 400.110 ;
        RECT 822.180 390.990 822.320 400.110 ;
        RECT 822.120 390.670 822.380 390.990 ;
        RECT 2021.800 390.670 2022.060 390.990 ;
        RECT 2021.860 1.770 2022.000 390.670 ;
        RECT 2023.950 1.770 2024.510 2.400 ;
        RECT 2021.860 1.630 2024.510 1.770 ;
        RECT 2023.950 -4.800 2024.510 1.630 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 822.090 135.220 822.410 135.280 ;
        RECT 2035.570 135.220 2035.890 135.280 ;
        RECT 822.090 135.080 2035.890 135.220 ;
        RECT 822.090 135.020 822.410 135.080 ;
        RECT 2035.570 135.020 2035.890 135.080 ;
        RECT 2035.570 15.200 2035.890 15.260 ;
        RECT 2042.010 15.200 2042.330 15.260 ;
        RECT 2035.570 15.060 2042.330 15.200 ;
        RECT 2035.570 15.000 2035.890 15.060 ;
        RECT 2042.010 15.000 2042.330 15.060 ;
      LAYER via ;
        RECT 822.120 135.020 822.380 135.280 ;
        RECT 2035.600 135.020 2035.860 135.280 ;
        RECT 2035.600 15.000 2035.860 15.260 ;
        RECT 2042.040 15.000 2042.300 15.260 ;
      LAYER met2 ;
        RECT 826.610 400.250 826.890 404.000 ;
        RECT 825.400 400.110 826.890 400.250 ;
        RECT 825.400 324.370 825.540 400.110 ;
        RECT 826.610 400.000 826.890 400.110 ;
        RECT 822.180 324.230 825.540 324.370 ;
        RECT 822.180 135.310 822.320 324.230 ;
        RECT 822.120 134.990 822.380 135.310 ;
        RECT 2035.600 134.990 2035.860 135.310 ;
        RECT 2035.660 15.290 2035.800 134.990 ;
        RECT 2035.600 14.970 2035.860 15.290 ;
        RECT 2042.040 14.970 2042.300 15.290 ;
        RECT 2042.100 2.400 2042.240 14.970 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.310 386.820 434.630 386.880 ;
        RECT 444.890 386.820 445.210 386.880 ;
        RECT 434.310 386.680 445.210 386.820 ;
        RECT 434.310 386.620 434.630 386.680 ;
        RECT 444.890 386.620 445.210 386.680 ;
      LAYER via ;
        RECT 434.340 386.620 434.600 386.880 ;
        RECT 444.920 386.620 445.180 386.880 ;
      LAYER met2 ;
        RECT 434.230 400.180 434.510 404.000 ;
        RECT 434.230 400.000 434.540 400.180 ;
        RECT 434.400 386.910 434.540 400.000 ;
        RECT 434.340 386.590 434.600 386.910 ;
        RECT 444.920 386.590 445.180 386.910 ;
        RECT 444.980 17.525 445.120 386.590 ;
        RECT 444.910 17.155 445.190 17.525 ;
        RECT 765.070 17.155 765.350 17.525 ;
        RECT 765.140 2.400 765.280 17.155 ;
        RECT 764.930 -4.800 765.490 2.400 ;
      LAYER via2 ;
        RECT 444.910 17.200 445.190 17.480 ;
        RECT 765.070 17.200 765.350 17.480 ;
      LAYER met3 ;
        RECT 444.885 17.490 445.215 17.505 ;
        RECT 765.045 17.490 765.375 17.505 ;
        RECT 444.885 17.190 765.375 17.490 ;
        RECT 444.885 17.175 445.215 17.190 ;
        RECT 765.045 17.175 765.375 17.190 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 832.210 390.560 832.530 390.620 ;
        RECT 2056.270 390.560 2056.590 390.620 ;
        RECT 832.210 390.420 2056.590 390.560 ;
        RECT 832.210 390.360 832.530 390.420 ;
        RECT 2056.270 390.360 2056.590 390.420 ;
      LAYER via ;
        RECT 832.240 390.360 832.500 390.620 ;
        RECT 2056.300 390.360 2056.560 390.620 ;
      LAYER met2 ;
        RECT 832.130 400.180 832.410 404.000 ;
        RECT 832.130 400.000 832.440 400.180 ;
        RECT 832.300 390.650 832.440 400.000 ;
        RECT 832.240 390.330 832.500 390.650 ;
        RECT 2056.300 390.330 2056.560 390.650 ;
        RECT 2056.360 82.870 2056.500 390.330 ;
        RECT 2056.360 82.730 2059.720 82.870 ;
        RECT 2059.580 2.400 2059.720 82.730 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 836.350 134.880 836.670 134.940 ;
        RECT 2076.970 134.880 2077.290 134.940 ;
        RECT 836.350 134.740 2077.290 134.880 ;
        RECT 836.350 134.680 836.670 134.740 ;
        RECT 2076.970 134.680 2077.290 134.740 ;
      LAYER via ;
        RECT 836.380 134.680 836.640 134.940 ;
        RECT 2077.000 134.680 2077.260 134.940 ;
      LAYER met2 ;
        RECT 837.190 400.250 837.470 404.000 ;
        RECT 836.440 400.110 837.470 400.250 ;
        RECT 836.440 134.970 836.580 400.110 ;
        RECT 837.190 400.000 837.470 400.110 ;
        RECT 836.380 134.650 836.640 134.970 ;
        RECT 2077.000 134.650 2077.260 134.970 ;
        RECT 2077.060 82.870 2077.200 134.650 ;
        RECT 2077.060 82.730 2077.660 82.870 ;
        RECT 2077.520 2.400 2077.660 82.730 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.790 390.220 843.110 390.280 ;
        RECT 2090.770 390.220 2091.090 390.280 ;
        RECT 842.790 390.080 2091.090 390.220 ;
        RECT 842.790 390.020 843.110 390.080 ;
        RECT 2090.770 390.020 2091.090 390.080 ;
      LAYER via ;
        RECT 842.820 390.020 843.080 390.280 ;
        RECT 2090.800 390.020 2091.060 390.280 ;
      LAYER met2 ;
        RECT 842.710 400.180 842.990 404.000 ;
        RECT 842.710 400.000 843.020 400.180 ;
        RECT 842.880 390.310 843.020 400.000 ;
        RECT 842.820 389.990 843.080 390.310 ;
        RECT 2090.800 389.990 2091.060 390.310 ;
        RECT 2090.860 82.870 2091.000 389.990 ;
        RECT 2090.860 82.730 2092.840 82.870 ;
        RECT 2092.700 1.770 2092.840 82.730 ;
        RECT 2094.790 1.770 2095.350 2.400 ;
        RECT 2092.700 1.630 2095.350 1.770 ;
        RECT 2094.790 -4.800 2095.350 1.630 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.790 134.540 843.110 134.600 ;
        RECT 2111.470 134.540 2111.790 134.600 ;
        RECT 842.790 134.400 2111.790 134.540 ;
        RECT 842.790 134.340 843.110 134.400 ;
        RECT 2111.470 134.340 2111.790 134.400 ;
      LAYER via ;
        RECT 842.820 134.340 843.080 134.600 ;
        RECT 2111.500 134.340 2111.760 134.600 ;
      LAYER met2 ;
        RECT 848.230 400.250 848.510 404.000 ;
        RECT 847.020 400.110 848.510 400.250 ;
        RECT 847.020 324.370 847.160 400.110 ;
        RECT 848.230 400.000 848.510 400.110 ;
        RECT 842.880 324.230 847.160 324.370 ;
        RECT 842.880 134.630 843.020 324.230 ;
        RECT 842.820 134.310 843.080 134.630 ;
        RECT 2111.500 134.310 2111.760 134.630 ;
        RECT 2111.560 82.870 2111.700 134.310 ;
        RECT 2111.560 82.730 2113.080 82.870 ;
        RECT 2112.940 2.400 2113.080 82.730 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 853.830 389.880 854.150 389.940 ;
        RECT 2125.270 389.880 2125.590 389.940 ;
        RECT 853.830 389.740 2125.590 389.880 ;
        RECT 853.830 389.680 854.150 389.740 ;
        RECT 2125.270 389.680 2125.590 389.740 ;
      LAYER via ;
        RECT 853.860 389.680 854.120 389.940 ;
        RECT 2125.300 389.680 2125.560 389.940 ;
      LAYER met2 ;
        RECT 853.750 400.180 854.030 404.000 ;
        RECT 853.750 400.000 854.060 400.180 ;
        RECT 853.920 389.970 854.060 400.000 ;
        RECT 853.860 389.650 854.120 389.970 ;
        RECT 2125.300 389.650 2125.560 389.970 ;
        RECT 2125.360 82.870 2125.500 389.650 ;
        RECT 2125.360 82.730 2128.720 82.870 ;
        RECT 2128.580 1.770 2128.720 82.730 ;
        RECT 2130.670 1.770 2131.230 2.400 ;
        RECT 2128.580 1.630 2131.230 1.770 ;
        RECT 2130.670 -4.800 2131.230 1.630 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 855.670 375.600 855.990 375.660 ;
        RECT 857.970 375.600 858.290 375.660 ;
        RECT 855.670 375.460 858.290 375.600 ;
        RECT 855.670 375.400 855.990 375.460 ;
        RECT 857.970 375.400 858.290 375.460 ;
        RECT 855.670 15.540 855.990 15.600 ;
        RECT 855.670 15.400 2063.170 15.540 ;
        RECT 855.670 15.340 855.990 15.400 ;
        RECT 2063.030 15.200 2063.170 15.400 ;
        RECT 2148.270 15.200 2148.590 15.260 ;
        RECT 2063.030 15.060 2148.590 15.200 ;
        RECT 2148.270 15.000 2148.590 15.060 ;
      LAYER via ;
        RECT 855.700 375.400 855.960 375.660 ;
        RECT 858.000 375.400 858.260 375.660 ;
        RECT 855.700 15.340 855.960 15.600 ;
        RECT 2148.300 15.000 2148.560 15.260 ;
      LAYER met2 ;
        RECT 859.270 400.250 859.550 404.000 ;
        RECT 858.060 400.110 859.550 400.250 ;
        RECT 858.060 375.690 858.200 400.110 ;
        RECT 859.270 400.000 859.550 400.110 ;
        RECT 855.700 375.370 855.960 375.690 ;
        RECT 858.000 375.370 858.260 375.690 ;
        RECT 855.760 15.630 855.900 375.370 ;
        RECT 855.700 15.310 855.960 15.630 ;
        RECT 2148.300 14.970 2148.560 15.290 ;
        RECT 2148.360 2.400 2148.500 14.970 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 862.570 377.640 862.890 377.700 ;
        RECT 863.490 377.640 863.810 377.700 ;
        RECT 862.570 377.500 863.810 377.640 ;
        RECT 862.570 377.440 862.890 377.500 ;
        RECT 863.490 377.440 863.810 377.500 ;
        RECT 862.570 15.880 862.890 15.940 ;
        RECT 2166.210 15.880 2166.530 15.940 ;
        RECT 862.570 15.740 2166.530 15.880 ;
        RECT 862.570 15.680 862.890 15.740 ;
        RECT 2166.210 15.680 2166.530 15.740 ;
      LAYER via ;
        RECT 862.600 377.440 862.860 377.700 ;
        RECT 863.520 377.440 863.780 377.700 ;
        RECT 862.600 15.680 862.860 15.940 ;
        RECT 2166.240 15.680 2166.500 15.940 ;
      LAYER met2 ;
        RECT 864.790 400.250 865.070 404.000 ;
        RECT 863.580 400.110 865.070 400.250 ;
        RECT 863.580 377.730 863.720 400.110 ;
        RECT 864.790 400.000 865.070 400.110 ;
        RECT 862.600 377.410 862.860 377.730 ;
        RECT 863.520 377.410 863.780 377.730 ;
        RECT 862.660 15.970 862.800 377.410 ;
        RECT 862.600 15.650 862.860 15.970 ;
        RECT 2166.240 15.650 2166.500 15.970 ;
        RECT 2166.300 2.400 2166.440 15.650 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.470 16.220 869.790 16.280 ;
        RECT 2183.690 16.220 2184.010 16.280 ;
        RECT 869.470 16.080 2184.010 16.220 ;
        RECT 869.470 16.020 869.790 16.080 ;
        RECT 2183.690 16.020 2184.010 16.080 ;
      LAYER via ;
        RECT 869.500 16.020 869.760 16.280 ;
        RECT 2183.720 16.020 2183.980 16.280 ;
      LAYER met2 ;
        RECT 869.850 400.250 870.130 404.000 ;
        RECT 869.560 400.110 870.130 400.250 ;
        RECT 869.560 16.310 869.700 400.110 ;
        RECT 869.850 400.000 870.130 400.110 ;
        RECT 869.500 15.990 869.760 16.310 ;
        RECT 2183.720 15.990 2183.980 16.310 ;
        RECT 2183.780 2.400 2183.920 15.990 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 869.930 376.280 870.250 376.340 ;
        RECT 874.070 376.280 874.390 376.340 ;
        RECT 869.930 376.140 874.390 376.280 ;
        RECT 869.930 376.080 870.250 376.140 ;
        RECT 874.070 376.080 874.390 376.140 ;
        RECT 869.930 16.560 870.250 16.620 ;
        RECT 2201.170 16.560 2201.490 16.620 ;
        RECT 869.930 16.420 2201.490 16.560 ;
        RECT 869.930 16.360 870.250 16.420 ;
        RECT 2201.170 16.360 2201.490 16.420 ;
      LAYER via ;
        RECT 869.960 376.080 870.220 376.340 ;
        RECT 874.100 376.080 874.360 376.340 ;
        RECT 869.960 16.360 870.220 16.620 ;
        RECT 2201.200 16.360 2201.460 16.620 ;
      LAYER met2 ;
        RECT 875.370 400.250 875.650 404.000 ;
        RECT 874.160 400.110 875.650 400.250 ;
        RECT 874.160 376.370 874.300 400.110 ;
        RECT 875.370 400.000 875.650 400.110 ;
        RECT 869.960 376.050 870.220 376.370 ;
        RECT 874.100 376.050 874.360 376.370 ;
        RECT 870.020 16.650 870.160 376.050 ;
        RECT 869.960 16.330 870.220 16.650 ;
        RECT 2201.200 16.330 2201.460 16.650 ;
        RECT 2201.260 8.570 2201.400 16.330 ;
        RECT 2201.260 8.430 2201.860 8.570 ;
        RECT 2201.720 2.400 2201.860 8.430 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 876.370 376.280 876.690 376.340 ;
        RECT 879.590 376.280 879.910 376.340 ;
        RECT 876.370 376.140 879.910 376.280 ;
        RECT 876.370 376.080 876.690 376.140 ;
        RECT 879.590 376.080 879.910 376.140 ;
        RECT 876.370 16.900 876.690 16.960 ;
        RECT 2219.110 16.900 2219.430 16.960 ;
        RECT 876.370 16.760 2219.430 16.900 ;
        RECT 876.370 16.700 876.690 16.760 ;
        RECT 2219.110 16.700 2219.430 16.760 ;
      LAYER via ;
        RECT 876.400 376.080 876.660 376.340 ;
        RECT 879.620 376.080 879.880 376.340 ;
        RECT 876.400 16.700 876.660 16.960 ;
        RECT 2219.140 16.700 2219.400 16.960 ;
      LAYER met2 ;
        RECT 880.890 400.250 881.170 404.000 ;
        RECT 879.680 400.110 881.170 400.250 ;
        RECT 879.680 376.370 879.820 400.110 ;
        RECT 880.890 400.000 881.170 400.110 ;
        RECT 876.400 376.050 876.660 376.370 ;
        RECT 879.620 376.050 879.880 376.370 ;
        RECT 876.460 16.990 876.600 376.050 ;
        RECT 876.400 16.670 876.660 16.990 ;
        RECT 2219.140 16.670 2219.400 16.990 ;
        RECT 2219.200 2.400 2219.340 16.670 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 434.770 386.480 435.090 386.540 ;
        RECT 438.450 386.480 438.770 386.540 ;
        RECT 434.770 386.340 438.770 386.480 ;
        RECT 434.770 386.280 435.090 386.340 ;
        RECT 438.450 386.280 438.770 386.340 ;
      LAYER via ;
        RECT 434.800 386.280 435.060 386.540 ;
        RECT 438.480 386.280 438.740 386.540 ;
      LAYER met2 ;
        RECT 439.750 400.250 440.030 404.000 ;
        RECT 438.540 400.110 440.030 400.250 ;
        RECT 438.540 386.570 438.680 400.110 ;
        RECT 439.750 400.000 440.030 400.110 ;
        RECT 434.800 386.250 435.060 386.570 ;
        RECT 438.480 386.250 438.740 386.570 ;
        RECT 434.860 16.845 435.000 386.250 ;
        RECT 434.790 16.475 435.070 16.845 ;
        RECT 783.010 16.475 783.290 16.845 ;
        RECT 783.080 2.400 783.220 16.475 ;
        RECT 782.870 -4.800 783.430 2.400 ;
      LAYER via2 ;
        RECT 434.790 16.520 435.070 16.800 ;
        RECT 783.010 16.520 783.290 16.800 ;
      LAYER met3 ;
        RECT 434.765 16.810 435.095 16.825 ;
        RECT 782.985 16.810 783.315 16.825 ;
        RECT 434.765 16.510 783.315 16.810 ;
        RECT 434.765 16.495 435.095 16.510 ;
        RECT 782.985 16.495 783.315 16.510 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 883.270 376.280 883.590 376.340 ;
        RECT 885.110 376.280 885.430 376.340 ;
        RECT 883.270 376.140 885.430 376.280 ;
        RECT 883.270 376.080 883.590 376.140 ;
        RECT 885.110 376.080 885.430 376.140 ;
        RECT 883.270 20.640 883.590 20.700 ;
        RECT 2237.050 20.640 2237.370 20.700 ;
        RECT 883.270 20.500 2237.370 20.640 ;
        RECT 883.270 20.440 883.590 20.500 ;
        RECT 2237.050 20.440 2237.370 20.500 ;
      LAYER via ;
        RECT 883.300 376.080 883.560 376.340 ;
        RECT 885.140 376.080 885.400 376.340 ;
        RECT 883.300 20.440 883.560 20.700 ;
        RECT 2237.080 20.440 2237.340 20.700 ;
      LAYER met2 ;
        RECT 886.410 400.250 886.690 404.000 ;
        RECT 885.200 400.110 886.690 400.250 ;
        RECT 885.200 376.370 885.340 400.110 ;
        RECT 886.410 400.000 886.690 400.110 ;
        RECT 883.300 376.050 883.560 376.370 ;
        RECT 885.140 376.050 885.400 376.370 ;
        RECT 883.360 20.730 883.500 376.050 ;
        RECT 883.300 20.410 883.560 20.730 ;
        RECT 2237.080 20.410 2237.340 20.730 ;
        RECT 2237.140 2.400 2237.280 20.410 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 890.170 398.380 890.490 398.440 ;
        RECT 891.090 398.380 891.410 398.440 ;
        RECT 890.170 398.240 891.410 398.380 ;
        RECT 890.170 398.180 890.490 398.240 ;
        RECT 891.090 398.180 891.410 398.240 ;
        RECT 890.170 20.300 890.490 20.360 ;
        RECT 2254.530 20.300 2254.850 20.360 ;
        RECT 890.170 20.160 2254.850 20.300 ;
        RECT 890.170 20.100 890.490 20.160 ;
        RECT 2254.530 20.100 2254.850 20.160 ;
      LAYER via ;
        RECT 890.200 398.180 890.460 398.440 ;
        RECT 891.120 398.180 891.380 398.440 ;
        RECT 890.200 20.100 890.460 20.360 ;
        RECT 2254.560 20.100 2254.820 20.360 ;
      LAYER met2 ;
        RECT 891.930 400.250 892.210 404.000 ;
        RECT 891.180 400.110 892.210 400.250 ;
        RECT 891.180 398.470 891.320 400.110 ;
        RECT 891.930 400.000 892.210 400.110 ;
        RECT 890.200 398.150 890.460 398.470 ;
        RECT 891.120 398.150 891.380 398.470 ;
        RECT 890.260 20.390 890.400 398.150 ;
        RECT 890.200 20.070 890.460 20.390 ;
        RECT 2254.560 20.070 2254.820 20.390 ;
        RECT 2254.620 2.400 2254.760 20.070 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.530 19.960 897.850 20.020 ;
        RECT 2272.470 19.960 2272.790 20.020 ;
        RECT 897.530 19.820 2272.790 19.960 ;
        RECT 897.530 19.760 897.850 19.820 ;
        RECT 2272.470 19.760 2272.790 19.820 ;
      LAYER via ;
        RECT 897.560 19.760 897.820 20.020 ;
        RECT 2272.500 19.760 2272.760 20.020 ;
      LAYER met2 ;
        RECT 897.450 400.180 897.730 404.000 ;
        RECT 897.450 400.000 897.760 400.180 ;
        RECT 897.620 20.050 897.760 400.000 ;
        RECT 897.560 19.730 897.820 20.050 ;
        RECT 2272.500 19.730 2272.760 20.050 ;
        RECT 2272.560 2.400 2272.700 19.730 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.070 376.280 897.390 376.340 ;
        RECT 901.210 376.280 901.530 376.340 ;
        RECT 897.070 376.140 901.530 376.280 ;
        RECT 897.070 376.080 897.390 376.140 ;
        RECT 901.210 376.080 901.530 376.140 ;
        RECT 897.070 19.620 897.390 19.680 ;
        RECT 2290.410 19.620 2290.730 19.680 ;
        RECT 897.070 19.480 2290.730 19.620 ;
        RECT 897.070 19.420 897.390 19.480 ;
        RECT 2290.410 19.420 2290.730 19.480 ;
      LAYER via ;
        RECT 897.100 376.080 897.360 376.340 ;
        RECT 901.240 376.080 901.500 376.340 ;
        RECT 897.100 19.420 897.360 19.680 ;
        RECT 2290.440 19.420 2290.700 19.680 ;
      LAYER met2 ;
        RECT 902.510 400.250 902.790 404.000 ;
        RECT 901.300 400.110 902.790 400.250 ;
        RECT 901.300 376.370 901.440 400.110 ;
        RECT 902.510 400.000 902.790 400.110 ;
        RECT 897.100 376.050 897.360 376.370 ;
        RECT 901.240 376.050 901.500 376.370 ;
        RECT 897.160 19.710 897.300 376.050 ;
        RECT 897.100 19.390 897.360 19.710 ;
        RECT 2290.440 19.390 2290.700 19.710 ;
        RECT 2290.500 2.400 2290.640 19.390 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 903.970 376.280 904.290 376.340 ;
        RECT 906.730 376.280 907.050 376.340 ;
        RECT 903.970 376.140 907.050 376.280 ;
        RECT 903.970 376.080 904.290 376.140 ;
        RECT 906.730 376.080 907.050 376.140 ;
        RECT 903.970 19.280 904.290 19.340 ;
        RECT 2307.890 19.280 2308.210 19.340 ;
        RECT 903.970 19.140 2308.210 19.280 ;
        RECT 903.970 19.080 904.290 19.140 ;
        RECT 2307.890 19.080 2308.210 19.140 ;
      LAYER via ;
        RECT 904.000 376.080 904.260 376.340 ;
        RECT 906.760 376.080 907.020 376.340 ;
        RECT 904.000 19.080 904.260 19.340 ;
        RECT 2307.920 19.080 2308.180 19.340 ;
      LAYER met2 ;
        RECT 908.030 400.250 908.310 404.000 ;
        RECT 906.820 400.110 908.310 400.250 ;
        RECT 906.820 376.370 906.960 400.110 ;
        RECT 908.030 400.000 908.310 400.110 ;
        RECT 904.000 376.050 904.260 376.370 ;
        RECT 906.760 376.050 907.020 376.370 ;
        RECT 904.060 19.370 904.200 376.050 ;
        RECT 904.000 19.050 904.260 19.370 ;
        RECT 2307.920 19.050 2308.180 19.370 ;
        RECT 2307.980 2.400 2308.120 19.050 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 910.870 376.280 911.190 376.340 ;
        RECT 912.250 376.280 912.570 376.340 ;
        RECT 910.870 376.140 912.570 376.280 ;
        RECT 910.870 376.080 911.190 376.140 ;
        RECT 912.250 376.080 912.570 376.140 ;
        RECT 910.870 18.940 911.190 19.000 ;
        RECT 2325.830 18.940 2326.150 19.000 ;
        RECT 910.870 18.800 2326.150 18.940 ;
        RECT 910.870 18.740 911.190 18.800 ;
        RECT 2325.830 18.740 2326.150 18.800 ;
      LAYER via ;
        RECT 910.900 376.080 911.160 376.340 ;
        RECT 912.280 376.080 912.540 376.340 ;
        RECT 910.900 18.740 911.160 19.000 ;
        RECT 2325.860 18.740 2326.120 19.000 ;
      LAYER met2 ;
        RECT 913.550 400.250 913.830 404.000 ;
        RECT 912.340 400.110 913.830 400.250 ;
        RECT 912.340 376.370 912.480 400.110 ;
        RECT 913.550 400.000 913.830 400.110 ;
        RECT 910.900 376.050 911.160 376.370 ;
        RECT 912.280 376.050 912.540 376.370 ;
        RECT 910.960 19.030 911.100 376.050 ;
        RECT 910.900 18.710 911.160 19.030 ;
        RECT 2325.860 18.710 2326.120 19.030 ;
        RECT 2325.920 2.400 2326.060 18.710 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 917.770 18.600 918.090 18.660 ;
        RECT 2343.310 18.600 2343.630 18.660 ;
        RECT 917.770 18.460 2343.630 18.600 ;
        RECT 917.770 18.400 918.090 18.460 ;
        RECT 2343.310 18.400 2343.630 18.460 ;
      LAYER via ;
        RECT 917.800 18.400 918.060 18.660 ;
        RECT 2343.340 18.400 2343.600 18.660 ;
      LAYER met2 ;
        RECT 919.070 400.250 919.350 404.000 ;
        RECT 917.860 400.110 919.350 400.250 ;
        RECT 917.860 18.690 918.000 400.110 ;
        RECT 919.070 400.000 919.350 400.110 ;
        RECT 917.800 18.370 918.060 18.690 ;
        RECT 2343.340 18.370 2343.600 18.690 ;
        RECT 2343.400 2.400 2343.540 18.370 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 925.130 18.260 925.450 18.320 ;
        RECT 2361.250 18.260 2361.570 18.320 ;
        RECT 925.130 18.120 2361.570 18.260 ;
        RECT 925.130 18.060 925.450 18.120 ;
        RECT 2361.250 18.060 2361.570 18.120 ;
      LAYER via ;
        RECT 925.160 18.060 925.420 18.320 ;
        RECT 2361.280 18.060 2361.540 18.320 ;
      LAYER met2 ;
        RECT 924.590 400.250 924.870 404.000 ;
        RECT 924.590 400.110 925.360 400.250 ;
        RECT 924.590 400.000 924.870 400.110 ;
        RECT 925.220 18.350 925.360 400.110 ;
        RECT 925.160 18.030 925.420 18.350 ;
        RECT 2361.280 18.030 2361.540 18.350 ;
        RECT 2361.340 2.400 2361.480 18.030 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 924.670 376.280 924.990 376.340 ;
        RECT 928.810 376.280 929.130 376.340 ;
        RECT 924.670 376.140 929.130 376.280 ;
        RECT 924.670 376.080 924.990 376.140 ;
        RECT 928.810 376.080 929.130 376.140 ;
        RECT 924.670 17.920 924.990 17.980 ;
        RECT 2378.730 17.920 2379.050 17.980 ;
        RECT 924.670 17.780 2379.050 17.920 ;
        RECT 924.670 17.720 924.990 17.780 ;
        RECT 2378.730 17.720 2379.050 17.780 ;
      LAYER via ;
        RECT 924.700 376.080 924.960 376.340 ;
        RECT 928.840 376.080 929.100 376.340 ;
        RECT 924.700 17.720 924.960 17.980 ;
        RECT 2378.760 17.720 2379.020 17.980 ;
      LAYER met2 ;
        RECT 930.110 400.250 930.390 404.000 ;
        RECT 928.900 400.110 930.390 400.250 ;
        RECT 928.900 376.370 929.040 400.110 ;
        RECT 930.110 400.000 930.390 400.110 ;
        RECT 924.700 376.050 924.960 376.370 ;
        RECT 928.840 376.050 929.100 376.370 ;
        RECT 924.760 18.010 924.900 376.050 ;
        RECT 924.700 17.690 924.960 18.010 ;
        RECT 2378.760 17.690 2379.020 18.010 ;
        RECT 2378.820 2.400 2378.960 17.690 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 931.570 386.480 931.890 386.540 ;
        RECT 934.330 386.480 934.650 386.540 ;
        RECT 931.570 386.340 934.650 386.480 ;
        RECT 931.570 386.280 931.890 386.340 ;
        RECT 934.330 386.280 934.650 386.340 ;
        RECT 931.570 17.580 931.890 17.640 ;
        RECT 2366.310 17.580 2366.630 17.640 ;
        RECT 931.570 17.440 2366.630 17.580 ;
        RECT 931.570 17.380 931.890 17.440 ;
        RECT 2366.310 17.380 2366.630 17.440 ;
        RECT 2366.310 16.560 2366.630 16.620 ;
        RECT 2396.670 16.560 2396.990 16.620 ;
        RECT 2366.310 16.420 2396.990 16.560 ;
        RECT 2366.310 16.360 2366.630 16.420 ;
        RECT 2396.670 16.360 2396.990 16.420 ;
      LAYER via ;
        RECT 931.600 386.280 931.860 386.540 ;
        RECT 934.360 386.280 934.620 386.540 ;
        RECT 931.600 17.380 931.860 17.640 ;
        RECT 2366.340 17.380 2366.600 17.640 ;
        RECT 2366.340 16.360 2366.600 16.620 ;
        RECT 2396.700 16.360 2396.960 16.620 ;
      LAYER met2 ;
        RECT 935.170 400.250 935.450 404.000 ;
        RECT 934.420 400.110 935.450 400.250 ;
        RECT 934.420 386.570 934.560 400.110 ;
        RECT 935.170 400.000 935.450 400.110 ;
        RECT 931.600 386.250 931.860 386.570 ;
        RECT 934.360 386.250 934.620 386.570 ;
        RECT 931.660 17.670 931.800 386.250 ;
        RECT 931.600 17.350 931.860 17.670 ;
        RECT 2366.340 17.350 2366.600 17.670 ;
        RECT 2366.400 16.650 2366.540 17.350 ;
        RECT 2366.340 16.330 2366.600 16.650 ;
        RECT 2396.700 16.330 2396.960 16.650 ;
        RECT 2396.760 2.400 2396.900 16.330 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.670 386.140 441.990 386.200 ;
        RECT 443.970 386.140 444.290 386.200 ;
        RECT 441.670 386.000 444.290 386.140 ;
        RECT 441.670 385.940 441.990 386.000 ;
        RECT 443.970 385.940 444.290 386.000 ;
        RECT 441.670 33.560 441.990 33.620 ;
        RECT 559.430 33.560 559.750 33.620 ;
        RECT 441.670 33.420 559.750 33.560 ;
        RECT 441.670 33.360 441.990 33.420 ;
        RECT 559.430 33.360 559.750 33.420 ;
        RECT 559.430 18.600 559.750 18.660 ;
        RECT 800.470 18.600 800.790 18.660 ;
        RECT 559.430 18.460 800.790 18.600 ;
        RECT 559.430 18.400 559.750 18.460 ;
        RECT 800.470 18.400 800.790 18.460 ;
      LAYER via ;
        RECT 441.700 385.940 441.960 386.200 ;
        RECT 444.000 385.940 444.260 386.200 ;
        RECT 441.700 33.360 441.960 33.620 ;
        RECT 559.460 33.360 559.720 33.620 ;
        RECT 559.460 18.400 559.720 18.660 ;
        RECT 800.500 18.400 800.760 18.660 ;
      LAYER met2 ;
        RECT 445.270 400.250 445.550 404.000 ;
        RECT 444.060 400.110 445.550 400.250 ;
        RECT 444.060 386.230 444.200 400.110 ;
        RECT 445.270 400.000 445.550 400.110 ;
        RECT 441.700 385.910 441.960 386.230 ;
        RECT 444.000 385.910 444.260 386.230 ;
        RECT 441.760 33.650 441.900 385.910 ;
        RECT 441.700 33.330 441.960 33.650 ;
        RECT 559.460 33.330 559.720 33.650 ;
        RECT 559.520 18.690 559.660 33.330 ;
        RECT 559.460 18.370 559.720 18.690 ;
        RECT 800.500 18.370 800.760 18.690 ;
        RECT 800.560 2.400 800.700 18.370 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1083.370 376.280 1083.690 376.340 ;
        RECT 1088.430 376.280 1088.750 376.340 ;
        RECT 1083.370 376.140 1088.750 376.280 ;
        RECT 1083.370 376.080 1083.690 376.140 ;
        RECT 1088.430 376.080 1088.750 376.140 ;
      LAYER via ;
        RECT 1083.400 376.080 1083.660 376.340 ;
        RECT 1088.460 376.080 1088.720 376.340 ;
      LAYER met2 ;
        RECT 1089.730 400.250 1090.010 404.000 ;
        RECT 1088.520 400.110 1090.010 400.250 ;
        RECT 1088.520 376.370 1088.660 400.110 ;
        RECT 1089.730 400.000 1090.010 400.110 ;
        RECT 1083.400 376.050 1083.660 376.370 ;
        RECT 1088.460 376.050 1088.720 376.370 ;
        RECT 1083.460 106.605 1083.600 376.050 ;
        RECT 1083.390 106.235 1083.670 106.605 ;
        RECT 2898.090 106.235 2898.370 106.605 ;
        RECT 2898.160 1.770 2898.300 106.235 ;
        RECT 2898.870 1.770 2899.430 2.400 ;
        RECT 2898.160 1.630 2899.430 1.770 ;
        RECT 2898.870 -4.800 2899.430 1.630 ;
      LAYER via2 ;
        RECT 1083.390 106.280 1083.670 106.560 ;
        RECT 2898.090 106.280 2898.370 106.560 ;
      LAYER met3 ;
        RECT 1083.365 106.570 1083.695 106.585 ;
        RECT 2898.065 106.570 2898.395 106.585 ;
        RECT 1083.365 106.270 2898.395 106.570 ;
        RECT 1083.365 106.255 1083.695 106.270 ;
        RECT 2898.065 106.255 2898.395 106.270 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.190 17.240 1114.510 17.300 ;
        RECT 2904.970 17.240 2905.290 17.300 ;
        RECT 1114.190 17.100 2905.290 17.240 ;
        RECT 1114.190 17.040 1114.510 17.100 ;
        RECT 2904.970 17.040 2905.290 17.100 ;
      LAYER via ;
        RECT 1114.220 17.040 1114.480 17.300 ;
        RECT 2905.000 17.040 2905.260 17.300 ;
      LAYER met2 ;
        RECT 1114.210 462.555 1114.490 462.925 ;
        RECT 1114.280 17.330 1114.420 462.555 ;
        RECT 1114.220 17.010 1114.480 17.330 ;
        RECT 2905.000 17.010 2905.260 17.330 ;
        RECT 2905.060 2.400 2905.200 17.010 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 1114.210 462.600 1114.490 462.880 ;
      LAYER met3 ;
        RECT 1096.000 463.960 1100.000 464.560 ;
        RECT 1098.790 462.890 1099.090 463.960 ;
        RECT 1114.185 462.890 1114.515 462.905 ;
        RECT 1098.790 462.590 1114.515 462.890 ;
        RECT 1114.185 462.575 1114.515 462.590 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1091.650 389.540 1091.970 389.600 ;
        RECT 1127.990 389.540 1128.310 389.600 ;
        RECT 1091.650 389.400 1128.310 389.540 ;
        RECT 1091.650 389.340 1091.970 389.400 ;
        RECT 1127.990 389.340 1128.310 389.400 ;
        RECT 1127.990 31.860 1128.310 31.920 ;
        RECT 2910.950 31.860 2911.270 31.920 ;
        RECT 1127.990 31.720 2911.270 31.860 ;
        RECT 1127.990 31.660 1128.310 31.720 ;
        RECT 2910.950 31.660 2911.270 31.720 ;
      LAYER via ;
        RECT 1091.680 389.340 1091.940 389.600 ;
        RECT 1128.020 389.340 1128.280 389.600 ;
        RECT 1128.020 31.660 1128.280 31.920 ;
        RECT 2910.980 31.660 2911.240 31.920 ;
      LAYER met2 ;
        RECT 1091.570 400.180 1091.850 404.000 ;
        RECT 1091.570 400.000 1091.880 400.180 ;
        RECT 1091.740 389.630 1091.880 400.000 ;
        RECT 1091.680 389.310 1091.940 389.630 ;
        RECT 1128.020 389.310 1128.280 389.630 ;
        RECT 1128.080 31.950 1128.220 389.310 ;
        RECT 1128.020 31.630 1128.280 31.950 ;
        RECT 2910.980 31.630 2911.240 31.950 ;
        RECT 2911.040 2.400 2911.180 31.630 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1060.370 1007.660 1060.690 1007.720 ;
        RECT 2197.490 1007.660 2197.810 1007.720 ;
        RECT 1060.370 1007.520 2197.810 1007.660 ;
        RECT 1060.370 1007.460 1060.690 1007.520 ;
        RECT 2197.490 1007.460 2197.810 1007.520 ;
        RECT 2197.490 16.220 2197.810 16.280 ;
        RECT 2916.930 16.220 2917.250 16.280 ;
        RECT 2197.490 16.080 2917.250 16.220 ;
        RECT 2197.490 16.020 2197.810 16.080 ;
        RECT 2916.930 16.020 2917.250 16.080 ;
      LAYER via ;
        RECT 1060.400 1007.460 1060.660 1007.720 ;
        RECT 2197.520 1007.460 2197.780 1007.720 ;
        RECT 2197.520 16.020 2197.780 16.280 ;
        RECT 2916.960 16.020 2917.220 16.280 ;
      LAYER met2 ;
        RECT 1060.400 1007.430 1060.660 1007.750 ;
        RECT 2197.520 1007.430 2197.780 1007.750 ;
        RECT 1058.910 999.330 1059.190 1000.000 ;
        RECT 1060.460 999.330 1060.600 1007.430 ;
        RECT 1058.910 999.190 1060.600 999.330 ;
        RECT 1058.910 996.000 1059.190 999.190 ;
        RECT 2197.580 16.310 2197.720 1007.430 ;
        RECT 2197.520 15.990 2197.780 16.310 ;
        RECT 2916.960 15.990 2917.220 16.310 ;
        RECT 2917.020 2.400 2917.160 15.990 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
        RECT 188.970 1010.000 192.070 3529.150 ;
        RECT 368.970 1010.000 372.070 3529.150 ;
        RECT 548.970 1010.000 552.070 3529.150 ;
        RECT 728.970 1010.000 732.070 3529.150 ;
        RECT 908.970 1010.000 912.070 3529.150 ;
        RECT 1088.970 1010.000 1092.070 3529.150 ;
        RECT 221.040 410.640 222.640 987.760 ;
        RECT 374.640 410.640 376.240 987.760 ;
        RECT 528.240 410.640 529.840 987.760 ;
        RECT 681.840 410.640 683.440 987.760 ;
        RECT 835.440 410.640 837.040 987.760 ;
        RECT 989.040 410.640 990.640 987.760 ;
        RECT 188.970 -9.470 192.070 390.000 ;
        RECT 368.970 -9.470 372.070 390.000 ;
        RECT 548.970 -9.470 552.070 390.000 ;
        RECT 728.970 -9.470 732.070 390.000 ;
        RECT 908.970 -9.470 912.070 390.000 ;
        RECT 1088.970 -9.470 1092.070 390.000 ;
        RECT 1268.970 -9.470 1272.070 3529.150 ;
        RECT 1448.970 -9.470 1452.070 3529.150 ;
        RECT 1628.970 -9.470 1632.070 3529.150 ;
        RECT 1808.970 -9.470 1812.070 3529.150 ;
        RECT 1988.970 -9.470 1992.070 3529.150 ;
        RECT 2168.970 -9.470 2172.070 3529.150 ;
        RECT 2348.970 -9.470 2352.070 3529.150 ;
        RECT 2528.970 -9.470 2532.070 3529.150 ;
        RECT 2708.970 -9.470 2712.070 3529.150 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
      LAYER via4 ;
        RECT -9.870 3523.010 -8.690 3524.190 ;
        RECT -8.270 3523.010 -7.090 3524.190 ;
        RECT -9.870 3521.410 -8.690 3522.590 ;
        RECT -8.270 3521.410 -7.090 3522.590 ;
        RECT -9.870 3436.090 -8.690 3437.270 ;
        RECT -8.270 3436.090 -7.090 3437.270 ;
        RECT -9.870 3434.490 -8.690 3435.670 ;
        RECT -8.270 3434.490 -7.090 3435.670 ;
        RECT -9.870 3256.090 -8.690 3257.270 ;
        RECT -8.270 3256.090 -7.090 3257.270 ;
        RECT -9.870 3254.490 -8.690 3255.670 ;
        RECT -8.270 3254.490 -7.090 3255.670 ;
        RECT -9.870 3076.090 -8.690 3077.270 ;
        RECT -8.270 3076.090 -7.090 3077.270 ;
        RECT -9.870 3074.490 -8.690 3075.670 ;
        RECT -8.270 3074.490 -7.090 3075.670 ;
        RECT -9.870 2896.090 -8.690 2897.270 ;
        RECT -8.270 2896.090 -7.090 2897.270 ;
        RECT -9.870 2894.490 -8.690 2895.670 ;
        RECT -8.270 2894.490 -7.090 2895.670 ;
        RECT -9.870 2716.090 -8.690 2717.270 ;
        RECT -8.270 2716.090 -7.090 2717.270 ;
        RECT -9.870 2714.490 -8.690 2715.670 ;
        RECT -8.270 2714.490 -7.090 2715.670 ;
        RECT -9.870 2536.090 -8.690 2537.270 ;
        RECT -8.270 2536.090 -7.090 2537.270 ;
        RECT -9.870 2534.490 -8.690 2535.670 ;
        RECT -8.270 2534.490 -7.090 2535.670 ;
        RECT -9.870 2356.090 -8.690 2357.270 ;
        RECT -8.270 2356.090 -7.090 2357.270 ;
        RECT -9.870 2354.490 -8.690 2355.670 ;
        RECT -8.270 2354.490 -7.090 2355.670 ;
        RECT -9.870 2176.090 -8.690 2177.270 ;
        RECT -8.270 2176.090 -7.090 2177.270 ;
        RECT -9.870 2174.490 -8.690 2175.670 ;
        RECT -8.270 2174.490 -7.090 2175.670 ;
        RECT -9.870 1996.090 -8.690 1997.270 ;
        RECT -8.270 1996.090 -7.090 1997.270 ;
        RECT -9.870 1994.490 -8.690 1995.670 ;
        RECT -8.270 1994.490 -7.090 1995.670 ;
        RECT -9.870 1816.090 -8.690 1817.270 ;
        RECT -8.270 1816.090 -7.090 1817.270 ;
        RECT -9.870 1814.490 -8.690 1815.670 ;
        RECT -8.270 1814.490 -7.090 1815.670 ;
        RECT -9.870 1636.090 -8.690 1637.270 ;
        RECT -8.270 1636.090 -7.090 1637.270 ;
        RECT -9.870 1634.490 -8.690 1635.670 ;
        RECT -8.270 1634.490 -7.090 1635.670 ;
        RECT -9.870 1456.090 -8.690 1457.270 ;
        RECT -8.270 1456.090 -7.090 1457.270 ;
        RECT -9.870 1454.490 -8.690 1455.670 ;
        RECT -8.270 1454.490 -7.090 1455.670 ;
        RECT -9.870 1276.090 -8.690 1277.270 ;
        RECT -8.270 1276.090 -7.090 1277.270 ;
        RECT -9.870 1274.490 -8.690 1275.670 ;
        RECT -8.270 1274.490 -7.090 1275.670 ;
        RECT -9.870 1096.090 -8.690 1097.270 ;
        RECT -8.270 1096.090 -7.090 1097.270 ;
        RECT -9.870 1094.490 -8.690 1095.670 ;
        RECT -8.270 1094.490 -7.090 1095.670 ;
        RECT -9.870 916.090 -8.690 917.270 ;
        RECT -8.270 916.090 -7.090 917.270 ;
        RECT -9.870 914.490 -8.690 915.670 ;
        RECT -8.270 914.490 -7.090 915.670 ;
        RECT -9.870 736.090 -8.690 737.270 ;
        RECT -8.270 736.090 -7.090 737.270 ;
        RECT -9.870 734.490 -8.690 735.670 ;
        RECT -8.270 734.490 -7.090 735.670 ;
        RECT -9.870 556.090 -8.690 557.270 ;
        RECT -8.270 556.090 -7.090 557.270 ;
        RECT -9.870 554.490 -8.690 555.670 ;
        RECT -8.270 554.490 -7.090 555.670 ;
        RECT -9.870 376.090 -8.690 377.270 ;
        RECT -8.270 376.090 -7.090 377.270 ;
        RECT -9.870 374.490 -8.690 375.670 ;
        RECT -8.270 374.490 -7.090 375.670 ;
        RECT -9.870 196.090 -8.690 197.270 ;
        RECT -8.270 196.090 -7.090 197.270 ;
        RECT -9.870 194.490 -8.690 195.670 ;
        RECT -8.270 194.490 -7.090 195.670 ;
        RECT -9.870 16.090 -8.690 17.270 ;
        RECT -8.270 16.090 -7.090 17.270 ;
        RECT -9.870 14.490 -8.690 15.670 ;
        RECT -8.270 14.490 -7.090 15.670 ;
        RECT -9.870 -2.910 -8.690 -1.730 ;
        RECT -8.270 -2.910 -7.090 -1.730 ;
        RECT -9.870 -4.510 -8.690 -3.330 ;
        RECT -8.270 -4.510 -7.090 -3.330 ;
        RECT 9.130 3523.010 10.310 3524.190 ;
        RECT 10.730 3523.010 11.910 3524.190 ;
        RECT 9.130 3521.410 10.310 3522.590 ;
        RECT 10.730 3521.410 11.910 3522.590 ;
        RECT 9.130 3436.090 10.310 3437.270 ;
        RECT 10.730 3436.090 11.910 3437.270 ;
        RECT 9.130 3434.490 10.310 3435.670 ;
        RECT 10.730 3434.490 11.910 3435.670 ;
        RECT 9.130 3256.090 10.310 3257.270 ;
        RECT 10.730 3256.090 11.910 3257.270 ;
        RECT 9.130 3254.490 10.310 3255.670 ;
        RECT 10.730 3254.490 11.910 3255.670 ;
        RECT 9.130 3076.090 10.310 3077.270 ;
        RECT 10.730 3076.090 11.910 3077.270 ;
        RECT 9.130 3074.490 10.310 3075.670 ;
        RECT 10.730 3074.490 11.910 3075.670 ;
        RECT 9.130 2896.090 10.310 2897.270 ;
        RECT 10.730 2896.090 11.910 2897.270 ;
        RECT 9.130 2894.490 10.310 2895.670 ;
        RECT 10.730 2894.490 11.910 2895.670 ;
        RECT 9.130 2716.090 10.310 2717.270 ;
        RECT 10.730 2716.090 11.910 2717.270 ;
        RECT 9.130 2714.490 10.310 2715.670 ;
        RECT 10.730 2714.490 11.910 2715.670 ;
        RECT 9.130 2536.090 10.310 2537.270 ;
        RECT 10.730 2536.090 11.910 2537.270 ;
        RECT 9.130 2534.490 10.310 2535.670 ;
        RECT 10.730 2534.490 11.910 2535.670 ;
        RECT 9.130 2356.090 10.310 2357.270 ;
        RECT 10.730 2356.090 11.910 2357.270 ;
        RECT 9.130 2354.490 10.310 2355.670 ;
        RECT 10.730 2354.490 11.910 2355.670 ;
        RECT 9.130 2176.090 10.310 2177.270 ;
        RECT 10.730 2176.090 11.910 2177.270 ;
        RECT 9.130 2174.490 10.310 2175.670 ;
        RECT 10.730 2174.490 11.910 2175.670 ;
        RECT 9.130 1996.090 10.310 1997.270 ;
        RECT 10.730 1996.090 11.910 1997.270 ;
        RECT 9.130 1994.490 10.310 1995.670 ;
        RECT 10.730 1994.490 11.910 1995.670 ;
        RECT 9.130 1816.090 10.310 1817.270 ;
        RECT 10.730 1816.090 11.910 1817.270 ;
        RECT 9.130 1814.490 10.310 1815.670 ;
        RECT 10.730 1814.490 11.910 1815.670 ;
        RECT 9.130 1636.090 10.310 1637.270 ;
        RECT 10.730 1636.090 11.910 1637.270 ;
        RECT 9.130 1634.490 10.310 1635.670 ;
        RECT 10.730 1634.490 11.910 1635.670 ;
        RECT 9.130 1456.090 10.310 1457.270 ;
        RECT 10.730 1456.090 11.910 1457.270 ;
        RECT 9.130 1454.490 10.310 1455.670 ;
        RECT 10.730 1454.490 11.910 1455.670 ;
        RECT 9.130 1276.090 10.310 1277.270 ;
        RECT 10.730 1276.090 11.910 1277.270 ;
        RECT 9.130 1274.490 10.310 1275.670 ;
        RECT 10.730 1274.490 11.910 1275.670 ;
        RECT 9.130 1096.090 10.310 1097.270 ;
        RECT 10.730 1096.090 11.910 1097.270 ;
        RECT 9.130 1094.490 10.310 1095.670 ;
        RECT 10.730 1094.490 11.910 1095.670 ;
        RECT 189.130 3523.010 190.310 3524.190 ;
        RECT 190.730 3523.010 191.910 3524.190 ;
        RECT 189.130 3521.410 190.310 3522.590 ;
        RECT 190.730 3521.410 191.910 3522.590 ;
        RECT 189.130 3436.090 190.310 3437.270 ;
        RECT 190.730 3436.090 191.910 3437.270 ;
        RECT 189.130 3434.490 190.310 3435.670 ;
        RECT 190.730 3434.490 191.910 3435.670 ;
        RECT 189.130 3256.090 190.310 3257.270 ;
        RECT 190.730 3256.090 191.910 3257.270 ;
        RECT 189.130 3254.490 190.310 3255.670 ;
        RECT 190.730 3254.490 191.910 3255.670 ;
        RECT 189.130 3076.090 190.310 3077.270 ;
        RECT 190.730 3076.090 191.910 3077.270 ;
        RECT 189.130 3074.490 190.310 3075.670 ;
        RECT 190.730 3074.490 191.910 3075.670 ;
        RECT 189.130 2896.090 190.310 2897.270 ;
        RECT 190.730 2896.090 191.910 2897.270 ;
        RECT 189.130 2894.490 190.310 2895.670 ;
        RECT 190.730 2894.490 191.910 2895.670 ;
        RECT 189.130 2716.090 190.310 2717.270 ;
        RECT 190.730 2716.090 191.910 2717.270 ;
        RECT 189.130 2714.490 190.310 2715.670 ;
        RECT 190.730 2714.490 191.910 2715.670 ;
        RECT 189.130 2536.090 190.310 2537.270 ;
        RECT 190.730 2536.090 191.910 2537.270 ;
        RECT 189.130 2534.490 190.310 2535.670 ;
        RECT 190.730 2534.490 191.910 2535.670 ;
        RECT 189.130 2356.090 190.310 2357.270 ;
        RECT 190.730 2356.090 191.910 2357.270 ;
        RECT 189.130 2354.490 190.310 2355.670 ;
        RECT 190.730 2354.490 191.910 2355.670 ;
        RECT 189.130 2176.090 190.310 2177.270 ;
        RECT 190.730 2176.090 191.910 2177.270 ;
        RECT 189.130 2174.490 190.310 2175.670 ;
        RECT 190.730 2174.490 191.910 2175.670 ;
        RECT 189.130 1996.090 190.310 1997.270 ;
        RECT 190.730 1996.090 191.910 1997.270 ;
        RECT 189.130 1994.490 190.310 1995.670 ;
        RECT 190.730 1994.490 191.910 1995.670 ;
        RECT 189.130 1816.090 190.310 1817.270 ;
        RECT 190.730 1816.090 191.910 1817.270 ;
        RECT 189.130 1814.490 190.310 1815.670 ;
        RECT 190.730 1814.490 191.910 1815.670 ;
        RECT 189.130 1636.090 190.310 1637.270 ;
        RECT 190.730 1636.090 191.910 1637.270 ;
        RECT 189.130 1634.490 190.310 1635.670 ;
        RECT 190.730 1634.490 191.910 1635.670 ;
        RECT 189.130 1456.090 190.310 1457.270 ;
        RECT 190.730 1456.090 191.910 1457.270 ;
        RECT 189.130 1454.490 190.310 1455.670 ;
        RECT 190.730 1454.490 191.910 1455.670 ;
        RECT 189.130 1276.090 190.310 1277.270 ;
        RECT 190.730 1276.090 191.910 1277.270 ;
        RECT 189.130 1274.490 190.310 1275.670 ;
        RECT 190.730 1274.490 191.910 1275.670 ;
        RECT 189.130 1096.090 190.310 1097.270 ;
        RECT 190.730 1096.090 191.910 1097.270 ;
        RECT 189.130 1094.490 190.310 1095.670 ;
        RECT 190.730 1094.490 191.910 1095.670 ;
        RECT 369.130 3523.010 370.310 3524.190 ;
        RECT 370.730 3523.010 371.910 3524.190 ;
        RECT 369.130 3521.410 370.310 3522.590 ;
        RECT 370.730 3521.410 371.910 3522.590 ;
        RECT 369.130 3436.090 370.310 3437.270 ;
        RECT 370.730 3436.090 371.910 3437.270 ;
        RECT 369.130 3434.490 370.310 3435.670 ;
        RECT 370.730 3434.490 371.910 3435.670 ;
        RECT 369.130 3256.090 370.310 3257.270 ;
        RECT 370.730 3256.090 371.910 3257.270 ;
        RECT 369.130 3254.490 370.310 3255.670 ;
        RECT 370.730 3254.490 371.910 3255.670 ;
        RECT 369.130 3076.090 370.310 3077.270 ;
        RECT 370.730 3076.090 371.910 3077.270 ;
        RECT 369.130 3074.490 370.310 3075.670 ;
        RECT 370.730 3074.490 371.910 3075.670 ;
        RECT 369.130 2896.090 370.310 2897.270 ;
        RECT 370.730 2896.090 371.910 2897.270 ;
        RECT 369.130 2894.490 370.310 2895.670 ;
        RECT 370.730 2894.490 371.910 2895.670 ;
        RECT 369.130 2716.090 370.310 2717.270 ;
        RECT 370.730 2716.090 371.910 2717.270 ;
        RECT 369.130 2714.490 370.310 2715.670 ;
        RECT 370.730 2714.490 371.910 2715.670 ;
        RECT 369.130 2536.090 370.310 2537.270 ;
        RECT 370.730 2536.090 371.910 2537.270 ;
        RECT 369.130 2534.490 370.310 2535.670 ;
        RECT 370.730 2534.490 371.910 2535.670 ;
        RECT 369.130 2356.090 370.310 2357.270 ;
        RECT 370.730 2356.090 371.910 2357.270 ;
        RECT 369.130 2354.490 370.310 2355.670 ;
        RECT 370.730 2354.490 371.910 2355.670 ;
        RECT 369.130 2176.090 370.310 2177.270 ;
        RECT 370.730 2176.090 371.910 2177.270 ;
        RECT 369.130 2174.490 370.310 2175.670 ;
        RECT 370.730 2174.490 371.910 2175.670 ;
        RECT 369.130 1996.090 370.310 1997.270 ;
        RECT 370.730 1996.090 371.910 1997.270 ;
        RECT 369.130 1994.490 370.310 1995.670 ;
        RECT 370.730 1994.490 371.910 1995.670 ;
        RECT 369.130 1816.090 370.310 1817.270 ;
        RECT 370.730 1816.090 371.910 1817.270 ;
        RECT 369.130 1814.490 370.310 1815.670 ;
        RECT 370.730 1814.490 371.910 1815.670 ;
        RECT 369.130 1636.090 370.310 1637.270 ;
        RECT 370.730 1636.090 371.910 1637.270 ;
        RECT 369.130 1634.490 370.310 1635.670 ;
        RECT 370.730 1634.490 371.910 1635.670 ;
        RECT 369.130 1456.090 370.310 1457.270 ;
        RECT 370.730 1456.090 371.910 1457.270 ;
        RECT 369.130 1454.490 370.310 1455.670 ;
        RECT 370.730 1454.490 371.910 1455.670 ;
        RECT 369.130 1276.090 370.310 1277.270 ;
        RECT 370.730 1276.090 371.910 1277.270 ;
        RECT 369.130 1274.490 370.310 1275.670 ;
        RECT 370.730 1274.490 371.910 1275.670 ;
        RECT 369.130 1096.090 370.310 1097.270 ;
        RECT 370.730 1096.090 371.910 1097.270 ;
        RECT 369.130 1094.490 370.310 1095.670 ;
        RECT 370.730 1094.490 371.910 1095.670 ;
        RECT 549.130 3523.010 550.310 3524.190 ;
        RECT 550.730 3523.010 551.910 3524.190 ;
        RECT 549.130 3521.410 550.310 3522.590 ;
        RECT 550.730 3521.410 551.910 3522.590 ;
        RECT 549.130 3436.090 550.310 3437.270 ;
        RECT 550.730 3436.090 551.910 3437.270 ;
        RECT 549.130 3434.490 550.310 3435.670 ;
        RECT 550.730 3434.490 551.910 3435.670 ;
        RECT 549.130 3256.090 550.310 3257.270 ;
        RECT 550.730 3256.090 551.910 3257.270 ;
        RECT 549.130 3254.490 550.310 3255.670 ;
        RECT 550.730 3254.490 551.910 3255.670 ;
        RECT 549.130 3076.090 550.310 3077.270 ;
        RECT 550.730 3076.090 551.910 3077.270 ;
        RECT 549.130 3074.490 550.310 3075.670 ;
        RECT 550.730 3074.490 551.910 3075.670 ;
        RECT 549.130 2896.090 550.310 2897.270 ;
        RECT 550.730 2896.090 551.910 2897.270 ;
        RECT 549.130 2894.490 550.310 2895.670 ;
        RECT 550.730 2894.490 551.910 2895.670 ;
        RECT 549.130 2716.090 550.310 2717.270 ;
        RECT 550.730 2716.090 551.910 2717.270 ;
        RECT 549.130 2714.490 550.310 2715.670 ;
        RECT 550.730 2714.490 551.910 2715.670 ;
        RECT 549.130 2536.090 550.310 2537.270 ;
        RECT 550.730 2536.090 551.910 2537.270 ;
        RECT 549.130 2534.490 550.310 2535.670 ;
        RECT 550.730 2534.490 551.910 2535.670 ;
        RECT 549.130 2356.090 550.310 2357.270 ;
        RECT 550.730 2356.090 551.910 2357.270 ;
        RECT 549.130 2354.490 550.310 2355.670 ;
        RECT 550.730 2354.490 551.910 2355.670 ;
        RECT 549.130 2176.090 550.310 2177.270 ;
        RECT 550.730 2176.090 551.910 2177.270 ;
        RECT 549.130 2174.490 550.310 2175.670 ;
        RECT 550.730 2174.490 551.910 2175.670 ;
        RECT 549.130 1996.090 550.310 1997.270 ;
        RECT 550.730 1996.090 551.910 1997.270 ;
        RECT 549.130 1994.490 550.310 1995.670 ;
        RECT 550.730 1994.490 551.910 1995.670 ;
        RECT 549.130 1816.090 550.310 1817.270 ;
        RECT 550.730 1816.090 551.910 1817.270 ;
        RECT 549.130 1814.490 550.310 1815.670 ;
        RECT 550.730 1814.490 551.910 1815.670 ;
        RECT 549.130 1636.090 550.310 1637.270 ;
        RECT 550.730 1636.090 551.910 1637.270 ;
        RECT 549.130 1634.490 550.310 1635.670 ;
        RECT 550.730 1634.490 551.910 1635.670 ;
        RECT 549.130 1456.090 550.310 1457.270 ;
        RECT 550.730 1456.090 551.910 1457.270 ;
        RECT 549.130 1454.490 550.310 1455.670 ;
        RECT 550.730 1454.490 551.910 1455.670 ;
        RECT 549.130 1276.090 550.310 1277.270 ;
        RECT 550.730 1276.090 551.910 1277.270 ;
        RECT 549.130 1274.490 550.310 1275.670 ;
        RECT 550.730 1274.490 551.910 1275.670 ;
        RECT 549.130 1096.090 550.310 1097.270 ;
        RECT 550.730 1096.090 551.910 1097.270 ;
        RECT 549.130 1094.490 550.310 1095.670 ;
        RECT 550.730 1094.490 551.910 1095.670 ;
        RECT 729.130 3523.010 730.310 3524.190 ;
        RECT 730.730 3523.010 731.910 3524.190 ;
        RECT 729.130 3521.410 730.310 3522.590 ;
        RECT 730.730 3521.410 731.910 3522.590 ;
        RECT 729.130 3436.090 730.310 3437.270 ;
        RECT 730.730 3436.090 731.910 3437.270 ;
        RECT 729.130 3434.490 730.310 3435.670 ;
        RECT 730.730 3434.490 731.910 3435.670 ;
        RECT 729.130 3256.090 730.310 3257.270 ;
        RECT 730.730 3256.090 731.910 3257.270 ;
        RECT 729.130 3254.490 730.310 3255.670 ;
        RECT 730.730 3254.490 731.910 3255.670 ;
        RECT 729.130 3076.090 730.310 3077.270 ;
        RECT 730.730 3076.090 731.910 3077.270 ;
        RECT 729.130 3074.490 730.310 3075.670 ;
        RECT 730.730 3074.490 731.910 3075.670 ;
        RECT 729.130 2896.090 730.310 2897.270 ;
        RECT 730.730 2896.090 731.910 2897.270 ;
        RECT 729.130 2894.490 730.310 2895.670 ;
        RECT 730.730 2894.490 731.910 2895.670 ;
        RECT 729.130 2716.090 730.310 2717.270 ;
        RECT 730.730 2716.090 731.910 2717.270 ;
        RECT 729.130 2714.490 730.310 2715.670 ;
        RECT 730.730 2714.490 731.910 2715.670 ;
        RECT 729.130 2536.090 730.310 2537.270 ;
        RECT 730.730 2536.090 731.910 2537.270 ;
        RECT 729.130 2534.490 730.310 2535.670 ;
        RECT 730.730 2534.490 731.910 2535.670 ;
        RECT 729.130 2356.090 730.310 2357.270 ;
        RECT 730.730 2356.090 731.910 2357.270 ;
        RECT 729.130 2354.490 730.310 2355.670 ;
        RECT 730.730 2354.490 731.910 2355.670 ;
        RECT 729.130 2176.090 730.310 2177.270 ;
        RECT 730.730 2176.090 731.910 2177.270 ;
        RECT 729.130 2174.490 730.310 2175.670 ;
        RECT 730.730 2174.490 731.910 2175.670 ;
        RECT 729.130 1996.090 730.310 1997.270 ;
        RECT 730.730 1996.090 731.910 1997.270 ;
        RECT 729.130 1994.490 730.310 1995.670 ;
        RECT 730.730 1994.490 731.910 1995.670 ;
        RECT 729.130 1816.090 730.310 1817.270 ;
        RECT 730.730 1816.090 731.910 1817.270 ;
        RECT 729.130 1814.490 730.310 1815.670 ;
        RECT 730.730 1814.490 731.910 1815.670 ;
        RECT 729.130 1636.090 730.310 1637.270 ;
        RECT 730.730 1636.090 731.910 1637.270 ;
        RECT 729.130 1634.490 730.310 1635.670 ;
        RECT 730.730 1634.490 731.910 1635.670 ;
        RECT 729.130 1456.090 730.310 1457.270 ;
        RECT 730.730 1456.090 731.910 1457.270 ;
        RECT 729.130 1454.490 730.310 1455.670 ;
        RECT 730.730 1454.490 731.910 1455.670 ;
        RECT 729.130 1276.090 730.310 1277.270 ;
        RECT 730.730 1276.090 731.910 1277.270 ;
        RECT 729.130 1274.490 730.310 1275.670 ;
        RECT 730.730 1274.490 731.910 1275.670 ;
        RECT 729.130 1096.090 730.310 1097.270 ;
        RECT 730.730 1096.090 731.910 1097.270 ;
        RECT 729.130 1094.490 730.310 1095.670 ;
        RECT 730.730 1094.490 731.910 1095.670 ;
        RECT 909.130 3523.010 910.310 3524.190 ;
        RECT 910.730 3523.010 911.910 3524.190 ;
        RECT 909.130 3521.410 910.310 3522.590 ;
        RECT 910.730 3521.410 911.910 3522.590 ;
        RECT 909.130 3436.090 910.310 3437.270 ;
        RECT 910.730 3436.090 911.910 3437.270 ;
        RECT 909.130 3434.490 910.310 3435.670 ;
        RECT 910.730 3434.490 911.910 3435.670 ;
        RECT 909.130 3256.090 910.310 3257.270 ;
        RECT 910.730 3256.090 911.910 3257.270 ;
        RECT 909.130 3254.490 910.310 3255.670 ;
        RECT 910.730 3254.490 911.910 3255.670 ;
        RECT 909.130 3076.090 910.310 3077.270 ;
        RECT 910.730 3076.090 911.910 3077.270 ;
        RECT 909.130 3074.490 910.310 3075.670 ;
        RECT 910.730 3074.490 911.910 3075.670 ;
        RECT 909.130 2896.090 910.310 2897.270 ;
        RECT 910.730 2896.090 911.910 2897.270 ;
        RECT 909.130 2894.490 910.310 2895.670 ;
        RECT 910.730 2894.490 911.910 2895.670 ;
        RECT 909.130 2716.090 910.310 2717.270 ;
        RECT 910.730 2716.090 911.910 2717.270 ;
        RECT 909.130 2714.490 910.310 2715.670 ;
        RECT 910.730 2714.490 911.910 2715.670 ;
        RECT 909.130 2536.090 910.310 2537.270 ;
        RECT 910.730 2536.090 911.910 2537.270 ;
        RECT 909.130 2534.490 910.310 2535.670 ;
        RECT 910.730 2534.490 911.910 2535.670 ;
        RECT 909.130 2356.090 910.310 2357.270 ;
        RECT 910.730 2356.090 911.910 2357.270 ;
        RECT 909.130 2354.490 910.310 2355.670 ;
        RECT 910.730 2354.490 911.910 2355.670 ;
        RECT 909.130 2176.090 910.310 2177.270 ;
        RECT 910.730 2176.090 911.910 2177.270 ;
        RECT 909.130 2174.490 910.310 2175.670 ;
        RECT 910.730 2174.490 911.910 2175.670 ;
        RECT 909.130 1996.090 910.310 1997.270 ;
        RECT 910.730 1996.090 911.910 1997.270 ;
        RECT 909.130 1994.490 910.310 1995.670 ;
        RECT 910.730 1994.490 911.910 1995.670 ;
        RECT 909.130 1816.090 910.310 1817.270 ;
        RECT 910.730 1816.090 911.910 1817.270 ;
        RECT 909.130 1814.490 910.310 1815.670 ;
        RECT 910.730 1814.490 911.910 1815.670 ;
        RECT 909.130 1636.090 910.310 1637.270 ;
        RECT 910.730 1636.090 911.910 1637.270 ;
        RECT 909.130 1634.490 910.310 1635.670 ;
        RECT 910.730 1634.490 911.910 1635.670 ;
        RECT 909.130 1456.090 910.310 1457.270 ;
        RECT 910.730 1456.090 911.910 1457.270 ;
        RECT 909.130 1454.490 910.310 1455.670 ;
        RECT 910.730 1454.490 911.910 1455.670 ;
        RECT 909.130 1276.090 910.310 1277.270 ;
        RECT 910.730 1276.090 911.910 1277.270 ;
        RECT 909.130 1274.490 910.310 1275.670 ;
        RECT 910.730 1274.490 911.910 1275.670 ;
        RECT 909.130 1096.090 910.310 1097.270 ;
        RECT 910.730 1096.090 911.910 1097.270 ;
        RECT 909.130 1094.490 910.310 1095.670 ;
        RECT 910.730 1094.490 911.910 1095.670 ;
        RECT 1089.130 3523.010 1090.310 3524.190 ;
        RECT 1090.730 3523.010 1091.910 3524.190 ;
        RECT 1089.130 3521.410 1090.310 3522.590 ;
        RECT 1090.730 3521.410 1091.910 3522.590 ;
        RECT 1089.130 3436.090 1090.310 3437.270 ;
        RECT 1090.730 3436.090 1091.910 3437.270 ;
        RECT 1089.130 3434.490 1090.310 3435.670 ;
        RECT 1090.730 3434.490 1091.910 3435.670 ;
        RECT 1089.130 3256.090 1090.310 3257.270 ;
        RECT 1090.730 3256.090 1091.910 3257.270 ;
        RECT 1089.130 3254.490 1090.310 3255.670 ;
        RECT 1090.730 3254.490 1091.910 3255.670 ;
        RECT 1089.130 3076.090 1090.310 3077.270 ;
        RECT 1090.730 3076.090 1091.910 3077.270 ;
        RECT 1089.130 3074.490 1090.310 3075.670 ;
        RECT 1090.730 3074.490 1091.910 3075.670 ;
        RECT 1089.130 2896.090 1090.310 2897.270 ;
        RECT 1090.730 2896.090 1091.910 2897.270 ;
        RECT 1089.130 2894.490 1090.310 2895.670 ;
        RECT 1090.730 2894.490 1091.910 2895.670 ;
        RECT 1089.130 2716.090 1090.310 2717.270 ;
        RECT 1090.730 2716.090 1091.910 2717.270 ;
        RECT 1089.130 2714.490 1090.310 2715.670 ;
        RECT 1090.730 2714.490 1091.910 2715.670 ;
        RECT 1089.130 2536.090 1090.310 2537.270 ;
        RECT 1090.730 2536.090 1091.910 2537.270 ;
        RECT 1089.130 2534.490 1090.310 2535.670 ;
        RECT 1090.730 2534.490 1091.910 2535.670 ;
        RECT 1089.130 2356.090 1090.310 2357.270 ;
        RECT 1090.730 2356.090 1091.910 2357.270 ;
        RECT 1089.130 2354.490 1090.310 2355.670 ;
        RECT 1090.730 2354.490 1091.910 2355.670 ;
        RECT 1089.130 2176.090 1090.310 2177.270 ;
        RECT 1090.730 2176.090 1091.910 2177.270 ;
        RECT 1089.130 2174.490 1090.310 2175.670 ;
        RECT 1090.730 2174.490 1091.910 2175.670 ;
        RECT 1089.130 1996.090 1090.310 1997.270 ;
        RECT 1090.730 1996.090 1091.910 1997.270 ;
        RECT 1089.130 1994.490 1090.310 1995.670 ;
        RECT 1090.730 1994.490 1091.910 1995.670 ;
        RECT 1089.130 1816.090 1090.310 1817.270 ;
        RECT 1090.730 1816.090 1091.910 1817.270 ;
        RECT 1089.130 1814.490 1090.310 1815.670 ;
        RECT 1090.730 1814.490 1091.910 1815.670 ;
        RECT 1089.130 1636.090 1090.310 1637.270 ;
        RECT 1090.730 1636.090 1091.910 1637.270 ;
        RECT 1089.130 1634.490 1090.310 1635.670 ;
        RECT 1090.730 1634.490 1091.910 1635.670 ;
        RECT 1089.130 1456.090 1090.310 1457.270 ;
        RECT 1090.730 1456.090 1091.910 1457.270 ;
        RECT 1089.130 1454.490 1090.310 1455.670 ;
        RECT 1090.730 1454.490 1091.910 1455.670 ;
        RECT 1089.130 1276.090 1090.310 1277.270 ;
        RECT 1090.730 1276.090 1091.910 1277.270 ;
        RECT 1089.130 1274.490 1090.310 1275.670 ;
        RECT 1090.730 1274.490 1091.910 1275.670 ;
        RECT 1089.130 1096.090 1090.310 1097.270 ;
        RECT 1090.730 1096.090 1091.910 1097.270 ;
        RECT 1089.130 1094.490 1090.310 1095.670 ;
        RECT 1090.730 1094.490 1091.910 1095.670 ;
        RECT 1269.130 3523.010 1270.310 3524.190 ;
        RECT 1270.730 3523.010 1271.910 3524.190 ;
        RECT 1269.130 3521.410 1270.310 3522.590 ;
        RECT 1270.730 3521.410 1271.910 3522.590 ;
        RECT 1269.130 3436.090 1270.310 3437.270 ;
        RECT 1270.730 3436.090 1271.910 3437.270 ;
        RECT 1269.130 3434.490 1270.310 3435.670 ;
        RECT 1270.730 3434.490 1271.910 3435.670 ;
        RECT 1269.130 3256.090 1270.310 3257.270 ;
        RECT 1270.730 3256.090 1271.910 3257.270 ;
        RECT 1269.130 3254.490 1270.310 3255.670 ;
        RECT 1270.730 3254.490 1271.910 3255.670 ;
        RECT 1269.130 3076.090 1270.310 3077.270 ;
        RECT 1270.730 3076.090 1271.910 3077.270 ;
        RECT 1269.130 3074.490 1270.310 3075.670 ;
        RECT 1270.730 3074.490 1271.910 3075.670 ;
        RECT 1269.130 2896.090 1270.310 2897.270 ;
        RECT 1270.730 2896.090 1271.910 2897.270 ;
        RECT 1269.130 2894.490 1270.310 2895.670 ;
        RECT 1270.730 2894.490 1271.910 2895.670 ;
        RECT 1269.130 2716.090 1270.310 2717.270 ;
        RECT 1270.730 2716.090 1271.910 2717.270 ;
        RECT 1269.130 2714.490 1270.310 2715.670 ;
        RECT 1270.730 2714.490 1271.910 2715.670 ;
        RECT 1269.130 2536.090 1270.310 2537.270 ;
        RECT 1270.730 2536.090 1271.910 2537.270 ;
        RECT 1269.130 2534.490 1270.310 2535.670 ;
        RECT 1270.730 2534.490 1271.910 2535.670 ;
        RECT 1269.130 2356.090 1270.310 2357.270 ;
        RECT 1270.730 2356.090 1271.910 2357.270 ;
        RECT 1269.130 2354.490 1270.310 2355.670 ;
        RECT 1270.730 2354.490 1271.910 2355.670 ;
        RECT 1269.130 2176.090 1270.310 2177.270 ;
        RECT 1270.730 2176.090 1271.910 2177.270 ;
        RECT 1269.130 2174.490 1270.310 2175.670 ;
        RECT 1270.730 2174.490 1271.910 2175.670 ;
        RECT 1269.130 1996.090 1270.310 1997.270 ;
        RECT 1270.730 1996.090 1271.910 1997.270 ;
        RECT 1269.130 1994.490 1270.310 1995.670 ;
        RECT 1270.730 1994.490 1271.910 1995.670 ;
        RECT 1269.130 1816.090 1270.310 1817.270 ;
        RECT 1270.730 1816.090 1271.910 1817.270 ;
        RECT 1269.130 1814.490 1270.310 1815.670 ;
        RECT 1270.730 1814.490 1271.910 1815.670 ;
        RECT 1269.130 1636.090 1270.310 1637.270 ;
        RECT 1270.730 1636.090 1271.910 1637.270 ;
        RECT 1269.130 1634.490 1270.310 1635.670 ;
        RECT 1270.730 1634.490 1271.910 1635.670 ;
        RECT 1269.130 1456.090 1270.310 1457.270 ;
        RECT 1270.730 1456.090 1271.910 1457.270 ;
        RECT 1269.130 1454.490 1270.310 1455.670 ;
        RECT 1270.730 1454.490 1271.910 1455.670 ;
        RECT 1269.130 1276.090 1270.310 1277.270 ;
        RECT 1270.730 1276.090 1271.910 1277.270 ;
        RECT 1269.130 1274.490 1270.310 1275.670 ;
        RECT 1270.730 1274.490 1271.910 1275.670 ;
        RECT 1269.130 1096.090 1270.310 1097.270 ;
        RECT 1270.730 1096.090 1271.910 1097.270 ;
        RECT 1269.130 1094.490 1270.310 1095.670 ;
        RECT 1270.730 1094.490 1271.910 1095.670 ;
        RECT 9.130 916.090 10.310 917.270 ;
        RECT 10.730 916.090 11.910 917.270 ;
        RECT 9.130 914.490 10.310 915.670 ;
        RECT 10.730 914.490 11.910 915.670 ;
        RECT 9.130 736.090 10.310 737.270 ;
        RECT 10.730 736.090 11.910 737.270 ;
        RECT 9.130 734.490 10.310 735.670 ;
        RECT 10.730 734.490 11.910 735.670 ;
        RECT 9.130 556.090 10.310 557.270 ;
        RECT 10.730 556.090 11.910 557.270 ;
        RECT 9.130 554.490 10.310 555.670 ;
        RECT 10.730 554.490 11.910 555.670 ;
        RECT 221.250 916.090 222.430 917.270 ;
        RECT 221.250 914.490 222.430 915.670 ;
        RECT 221.250 736.090 222.430 737.270 ;
        RECT 221.250 734.490 222.430 735.670 ;
        RECT 221.250 556.090 222.430 557.270 ;
        RECT 221.250 554.490 222.430 555.670 ;
        RECT 374.850 916.090 376.030 917.270 ;
        RECT 374.850 914.490 376.030 915.670 ;
        RECT 374.850 736.090 376.030 737.270 ;
        RECT 374.850 734.490 376.030 735.670 ;
        RECT 374.850 556.090 376.030 557.270 ;
        RECT 374.850 554.490 376.030 555.670 ;
        RECT 528.450 916.090 529.630 917.270 ;
        RECT 528.450 914.490 529.630 915.670 ;
        RECT 528.450 736.090 529.630 737.270 ;
        RECT 528.450 734.490 529.630 735.670 ;
        RECT 528.450 556.090 529.630 557.270 ;
        RECT 528.450 554.490 529.630 555.670 ;
        RECT 682.050 916.090 683.230 917.270 ;
        RECT 682.050 914.490 683.230 915.670 ;
        RECT 682.050 736.090 683.230 737.270 ;
        RECT 682.050 734.490 683.230 735.670 ;
        RECT 682.050 556.090 683.230 557.270 ;
        RECT 682.050 554.490 683.230 555.670 ;
        RECT 835.650 916.090 836.830 917.270 ;
        RECT 835.650 914.490 836.830 915.670 ;
        RECT 835.650 736.090 836.830 737.270 ;
        RECT 835.650 734.490 836.830 735.670 ;
        RECT 835.650 556.090 836.830 557.270 ;
        RECT 835.650 554.490 836.830 555.670 ;
        RECT 989.250 916.090 990.430 917.270 ;
        RECT 989.250 914.490 990.430 915.670 ;
        RECT 989.250 736.090 990.430 737.270 ;
        RECT 989.250 734.490 990.430 735.670 ;
        RECT 989.250 556.090 990.430 557.270 ;
        RECT 989.250 554.490 990.430 555.670 ;
        RECT 1269.130 916.090 1270.310 917.270 ;
        RECT 1270.730 916.090 1271.910 917.270 ;
        RECT 1269.130 914.490 1270.310 915.670 ;
        RECT 1270.730 914.490 1271.910 915.670 ;
        RECT 1269.130 736.090 1270.310 737.270 ;
        RECT 1270.730 736.090 1271.910 737.270 ;
        RECT 1269.130 734.490 1270.310 735.670 ;
        RECT 1270.730 734.490 1271.910 735.670 ;
        RECT 1269.130 556.090 1270.310 557.270 ;
        RECT 1270.730 556.090 1271.910 557.270 ;
        RECT 1269.130 554.490 1270.310 555.670 ;
        RECT 1270.730 554.490 1271.910 555.670 ;
        RECT 9.130 376.090 10.310 377.270 ;
        RECT 10.730 376.090 11.910 377.270 ;
        RECT 9.130 374.490 10.310 375.670 ;
        RECT 10.730 374.490 11.910 375.670 ;
        RECT 9.130 196.090 10.310 197.270 ;
        RECT 10.730 196.090 11.910 197.270 ;
        RECT 9.130 194.490 10.310 195.670 ;
        RECT 10.730 194.490 11.910 195.670 ;
        RECT 9.130 16.090 10.310 17.270 ;
        RECT 10.730 16.090 11.910 17.270 ;
        RECT 9.130 14.490 10.310 15.670 ;
        RECT 10.730 14.490 11.910 15.670 ;
        RECT 9.130 -2.910 10.310 -1.730 ;
        RECT 10.730 -2.910 11.910 -1.730 ;
        RECT 9.130 -4.510 10.310 -3.330 ;
        RECT 10.730 -4.510 11.910 -3.330 ;
        RECT 189.130 376.090 190.310 377.270 ;
        RECT 190.730 376.090 191.910 377.270 ;
        RECT 189.130 374.490 190.310 375.670 ;
        RECT 190.730 374.490 191.910 375.670 ;
        RECT 189.130 196.090 190.310 197.270 ;
        RECT 190.730 196.090 191.910 197.270 ;
        RECT 189.130 194.490 190.310 195.670 ;
        RECT 190.730 194.490 191.910 195.670 ;
        RECT 189.130 16.090 190.310 17.270 ;
        RECT 190.730 16.090 191.910 17.270 ;
        RECT 189.130 14.490 190.310 15.670 ;
        RECT 190.730 14.490 191.910 15.670 ;
        RECT 189.130 -2.910 190.310 -1.730 ;
        RECT 190.730 -2.910 191.910 -1.730 ;
        RECT 189.130 -4.510 190.310 -3.330 ;
        RECT 190.730 -4.510 191.910 -3.330 ;
        RECT 369.130 376.090 370.310 377.270 ;
        RECT 370.730 376.090 371.910 377.270 ;
        RECT 369.130 374.490 370.310 375.670 ;
        RECT 370.730 374.490 371.910 375.670 ;
        RECT 369.130 196.090 370.310 197.270 ;
        RECT 370.730 196.090 371.910 197.270 ;
        RECT 369.130 194.490 370.310 195.670 ;
        RECT 370.730 194.490 371.910 195.670 ;
        RECT 369.130 16.090 370.310 17.270 ;
        RECT 370.730 16.090 371.910 17.270 ;
        RECT 369.130 14.490 370.310 15.670 ;
        RECT 370.730 14.490 371.910 15.670 ;
        RECT 369.130 -2.910 370.310 -1.730 ;
        RECT 370.730 -2.910 371.910 -1.730 ;
        RECT 369.130 -4.510 370.310 -3.330 ;
        RECT 370.730 -4.510 371.910 -3.330 ;
        RECT 549.130 376.090 550.310 377.270 ;
        RECT 550.730 376.090 551.910 377.270 ;
        RECT 549.130 374.490 550.310 375.670 ;
        RECT 550.730 374.490 551.910 375.670 ;
        RECT 549.130 196.090 550.310 197.270 ;
        RECT 550.730 196.090 551.910 197.270 ;
        RECT 549.130 194.490 550.310 195.670 ;
        RECT 550.730 194.490 551.910 195.670 ;
        RECT 549.130 16.090 550.310 17.270 ;
        RECT 550.730 16.090 551.910 17.270 ;
        RECT 549.130 14.490 550.310 15.670 ;
        RECT 550.730 14.490 551.910 15.670 ;
        RECT 549.130 -2.910 550.310 -1.730 ;
        RECT 550.730 -2.910 551.910 -1.730 ;
        RECT 549.130 -4.510 550.310 -3.330 ;
        RECT 550.730 -4.510 551.910 -3.330 ;
        RECT 729.130 376.090 730.310 377.270 ;
        RECT 730.730 376.090 731.910 377.270 ;
        RECT 729.130 374.490 730.310 375.670 ;
        RECT 730.730 374.490 731.910 375.670 ;
        RECT 729.130 196.090 730.310 197.270 ;
        RECT 730.730 196.090 731.910 197.270 ;
        RECT 729.130 194.490 730.310 195.670 ;
        RECT 730.730 194.490 731.910 195.670 ;
        RECT 729.130 16.090 730.310 17.270 ;
        RECT 730.730 16.090 731.910 17.270 ;
        RECT 729.130 14.490 730.310 15.670 ;
        RECT 730.730 14.490 731.910 15.670 ;
        RECT 729.130 -2.910 730.310 -1.730 ;
        RECT 730.730 -2.910 731.910 -1.730 ;
        RECT 729.130 -4.510 730.310 -3.330 ;
        RECT 730.730 -4.510 731.910 -3.330 ;
        RECT 909.130 376.090 910.310 377.270 ;
        RECT 910.730 376.090 911.910 377.270 ;
        RECT 909.130 374.490 910.310 375.670 ;
        RECT 910.730 374.490 911.910 375.670 ;
        RECT 909.130 196.090 910.310 197.270 ;
        RECT 910.730 196.090 911.910 197.270 ;
        RECT 909.130 194.490 910.310 195.670 ;
        RECT 910.730 194.490 911.910 195.670 ;
        RECT 909.130 16.090 910.310 17.270 ;
        RECT 910.730 16.090 911.910 17.270 ;
        RECT 909.130 14.490 910.310 15.670 ;
        RECT 910.730 14.490 911.910 15.670 ;
        RECT 909.130 -2.910 910.310 -1.730 ;
        RECT 910.730 -2.910 911.910 -1.730 ;
        RECT 909.130 -4.510 910.310 -3.330 ;
        RECT 910.730 -4.510 911.910 -3.330 ;
        RECT 1089.130 376.090 1090.310 377.270 ;
        RECT 1090.730 376.090 1091.910 377.270 ;
        RECT 1089.130 374.490 1090.310 375.670 ;
        RECT 1090.730 374.490 1091.910 375.670 ;
        RECT 1089.130 196.090 1090.310 197.270 ;
        RECT 1090.730 196.090 1091.910 197.270 ;
        RECT 1089.130 194.490 1090.310 195.670 ;
        RECT 1090.730 194.490 1091.910 195.670 ;
        RECT 1089.130 16.090 1090.310 17.270 ;
        RECT 1090.730 16.090 1091.910 17.270 ;
        RECT 1089.130 14.490 1090.310 15.670 ;
        RECT 1090.730 14.490 1091.910 15.670 ;
        RECT 1089.130 -2.910 1090.310 -1.730 ;
        RECT 1090.730 -2.910 1091.910 -1.730 ;
        RECT 1089.130 -4.510 1090.310 -3.330 ;
        RECT 1090.730 -4.510 1091.910 -3.330 ;
        RECT 1269.130 376.090 1270.310 377.270 ;
        RECT 1270.730 376.090 1271.910 377.270 ;
        RECT 1269.130 374.490 1270.310 375.670 ;
        RECT 1270.730 374.490 1271.910 375.670 ;
        RECT 1269.130 196.090 1270.310 197.270 ;
        RECT 1270.730 196.090 1271.910 197.270 ;
        RECT 1269.130 194.490 1270.310 195.670 ;
        RECT 1270.730 194.490 1271.910 195.670 ;
        RECT 1269.130 16.090 1270.310 17.270 ;
        RECT 1270.730 16.090 1271.910 17.270 ;
        RECT 1269.130 14.490 1270.310 15.670 ;
        RECT 1270.730 14.490 1271.910 15.670 ;
        RECT 1269.130 -2.910 1270.310 -1.730 ;
        RECT 1270.730 -2.910 1271.910 -1.730 ;
        RECT 1269.130 -4.510 1270.310 -3.330 ;
        RECT 1270.730 -4.510 1271.910 -3.330 ;
        RECT 1449.130 3523.010 1450.310 3524.190 ;
        RECT 1450.730 3523.010 1451.910 3524.190 ;
        RECT 1449.130 3521.410 1450.310 3522.590 ;
        RECT 1450.730 3521.410 1451.910 3522.590 ;
        RECT 1449.130 3436.090 1450.310 3437.270 ;
        RECT 1450.730 3436.090 1451.910 3437.270 ;
        RECT 1449.130 3434.490 1450.310 3435.670 ;
        RECT 1450.730 3434.490 1451.910 3435.670 ;
        RECT 1449.130 3256.090 1450.310 3257.270 ;
        RECT 1450.730 3256.090 1451.910 3257.270 ;
        RECT 1449.130 3254.490 1450.310 3255.670 ;
        RECT 1450.730 3254.490 1451.910 3255.670 ;
        RECT 1449.130 3076.090 1450.310 3077.270 ;
        RECT 1450.730 3076.090 1451.910 3077.270 ;
        RECT 1449.130 3074.490 1450.310 3075.670 ;
        RECT 1450.730 3074.490 1451.910 3075.670 ;
        RECT 1449.130 2896.090 1450.310 2897.270 ;
        RECT 1450.730 2896.090 1451.910 2897.270 ;
        RECT 1449.130 2894.490 1450.310 2895.670 ;
        RECT 1450.730 2894.490 1451.910 2895.670 ;
        RECT 1449.130 2716.090 1450.310 2717.270 ;
        RECT 1450.730 2716.090 1451.910 2717.270 ;
        RECT 1449.130 2714.490 1450.310 2715.670 ;
        RECT 1450.730 2714.490 1451.910 2715.670 ;
        RECT 1449.130 2536.090 1450.310 2537.270 ;
        RECT 1450.730 2536.090 1451.910 2537.270 ;
        RECT 1449.130 2534.490 1450.310 2535.670 ;
        RECT 1450.730 2534.490 1451.910 2535.670 ;
        RECT 1449.130 2356.090 1450.310 2357.270 ;
        RECT 1450.730 2356.090 1451.910 2357.270 ;
        RECT 1449.130 2354.490 1450.310 2355.670 ;
        RECT 1450.730 2354.490 1451.910 2355.670 ;
        RECT 1449.130 2176.090 1450.310 2177.270 ;
        RECT 1450.730 2176.090 1451.910 2177.270 ;
        RECT 1449.130 2174.490 1450.310 2175.670 ;
        RECT 1450.730 2174.490 1451.910 2175.670 ;
        RECT 1449.130 1996.090 1450.310 1997.270 ;
        RECT 1450.730 1996.090 1451.910 1997.270 ;
        RECT 1449.130 1994.490 1450.310 1995.670 ;
        RECT 1450.730 1994.490 1451.910 1995.670 ;
        RECT 1449.130 1816.090 1450.310 1817.270 ;
        RECT 1450.730 1816.090 1451.910 1817.270 ;
        RECT 1449.130 1814.490 1450.310 1815.670 ;
        RECT 1450.730 1814.490 1451.910 1815.670 ;
        RECT 1449.130 1636.090 1450.310 1637.270 ;
        RECT 1450.730 1636.090 1451.910 1637.270 ;
        RECT 1449.130 1634.490 1450.310 1635.670 ;
        RECT 1450.730 1634.490 1451.910 1635.670 ;
        RECT 1449.130 1456.090 1450.310 1457.270 ;
        RECT 1450.730 1456.090 1451.910 1457.270 ;
        RECT 1449.130 1454.490 1450.310 1455.670 ;
        RECT 1450.730 1454.490 1451.910 1455.670 ;
        RECT 1449.130 1276.090 1450.310 1277.270 ;
        RECT 1450.730 1276.090 1451.910 1277.270 ;
        RECT 1449.130 1274.490 1450.310 1275.670 ;
        RECT 1450.730 1274.490 1451.910 1275.670 ;
        RECT 1449.130 1096.090 1450.310 1097.270 ;
        RECT 1450.730 1096.090 1451.910 1097.270 ;
        RECT 1449.130 1094.490 1450.310 1095.670 ;
        RECT 1450.730 1094.490 1451.910 1095.670 ;
        RECT 1449.130 916.090 1450.310 917.270 ;
        RECT 1450.730 916.090 1451.910 917.270 ;
        RECT 1449.130 914.490 1450.310 915.670 ;
        RECT 1450.730 914.490 1451.910 915.670 ;
        RECT 1449.130 736.090 1450.310 737.270 ;
        RECT 1450.730 736.090 1451.910 737.270 ;
        RECT 1449.130 734.490 1450.310 735.670 ;
        RECT 1450.730 734.490 1451.910 735.670 ;
        RECT 1449.130 556.090 1450.310 557.270 ;
        RECT 1450.730 556.090 1451.910 557.270 ;
        RECT 1449.130 554.490 1450.310 555.670 ;
        RECT 1450.730 554.490 1451.910 555.670 ;
        RECT 1449.130 376.090 1450.310 377.270 ;
        RECT 1450.730 376.090 1451.910 377.270 ;
        RECT 1449.130 374.490 1450.310 375.670 ;
        RECT 1450.730 374.490 1451.910 375.670 ;
        RECT 1449.130 196.090 1450.310 197.270 ;
        RECT 1450.730 196.090 1451.910 197.270 ;
        RECT 1449.130 194.490 1450.310 195.670 ;
        RECT 1450.730 194.490 1451.910 195.670 ;
        RECT 1449.130 16.090 1450.310 17.270 ;
        RECT 1450.730 16.090 1451.910 17.270 ;
        RECT 1449.130 14.490 1450.310 15.670 ;
        RECT 1450.730 14.490 1451.910 15.670 ;
        RECT 1449.130 -2.910 1450.310 -1.730 ;
        RECT 1450.730 -2.910 1451.910 -1.730 ;
        RECT 1449.130 -4.510 1450.310 -3.330 ;
        RECT 1450.730 -4.510 1451.910 -3.330 ;
        RECT 1629.130 3523.010 1630.310 3524.190 ;
        RECT 1630.730 3523.010 1631.910 3524.190 ;
        RECT 1629.130 3521.410 1630.310 3522.590 ;
        RECT 1630.730 3521.410 1631.910 3522.590 ;
        RECT 1629.130 3436.090 1630.310 3437.270 ;
        RECT 1630.730 3436.090 1631.910 3437.270 ;
        RECT 1629.130 3434.490 1630.310 3435.670 ;
        RECT 1630.730 3434.490 1631.910 3435.670 ;
        RECT 1629.130 3256.090 1630.310 3257.270 ;
        RECT 1630.730 3256.090 1631.910 3257.270 ;
        RECT 1629.130 3254.490 1630.310 3255.670 ;
        RECT 1630.730 3254.490 1631.910 3255.670 ;
        RECT 1629.130 3076.090 1630.310 3077.270 ;
        RECT 1630.730 3076.090 1631.910 3077.270 ;
        RECT 1629.130 3074.490 1630.310 3075.670 ;
        RECT 1630.730 3074.490 1631.910 3075.670 ;
        RECT 1629.130 2896.090 1630.310 2897.270 ;
        RECT 1630.730 2896.090 1631.910 2897.270 ;
        RECT 1629.130 2894.490 1630.310 2895.670 ;
        RECT 1630.730 2894.490 1631.910 2895.670 ;
        RECT 1629.130 2716.090 1630.310 2717.270 ;
        RECT 1630.730 2716.090 1631.910 2717.270 ;
        RECT 1629.130 2714.490 1630.310 2715.670 ;
        RECT 1630.730 2714.490 1631.910 2715.670 ;
        RECT 1629.130 2536.090 1630.310 2537.270 ;
        RECT 1630.730 2536.090 1631.910 2537.270 ;
        RECT 1629.130 2534.490 1630.310 2535.670 ;
        RECT 1630.730 2534.490 1631.910 2535.670 ;
        RECT 1629.130 2356.090 1630.310 2357.270 ;
        RECT 1630.730 2356.090 1631.910 2357.270 ;
        RECT 1629.130 2354.490 1630.310 2355.670 ;
        RECT 1630.730 2354.490 1631.910 2355.670 ;
        RECT 1629.130 2176.090 1630.310 2177.270 ;
        RECT 1630.730 2176.090 1631.910 2177.270 ;
        RECT 1629.130 2174.490 1630.310 2175.670 ;
        RECT 1630.730 2174.490 1631.910 2175.670 ;
        RECT 1629.130 1996.090 1630.310 1997.270 ;
        RECT 1630.730 1996.090 1631.910 1997.270 ;
        RECT 1629.130 1994.490 1630.310 1995.670 ;
        RECT 1630.730 1994.490 1631.910 1995.670 ;
        RECT 1629.130 1816.090 1630.310 1817.270 ;
        RECT 1630.730 1816.090 1631.910 1817.270 ;
        RECT 1629.130 1814.490 1630.310 1815.670 ;
        RECT 1630.730 1814.490 1631.910 1815.670 ;
        RECT 1629.130 1636.090 1630.310 1637.270 ;
        RECT 1630.730 1636.090 1631.910 1637.270 ;
        RECT 1629.130 1634.490 1630.310 1635.670 ;
        RECT 1630.730 1634.490 1631.910 1635.670 ;
        RECT 1629.130 1456.090 1630.310 1457.270 ;
        RECT 1630.730 1456.090 1631.910 1457.270 ;
        RECT 1629.130 1454.490 1630.310 1455.670 ;
        RECT 1630.730 1454.490 1631.910 1455.670 ;
        RECT 1629.130 1276.090 1630.310 1277.270 ;
        RECT 1630.730 1276.090 1631.910 1277.270 ;
        RECT 1629.130 1274.490 1630.310 1275.670 ;
        RECT 1630.730 1274.490 1631.910 1275.670 ;
        RECT 1629.130 1096.090 1630.310 1097.270 ;
        RECT 1630.730 1096.090 1631.910 1097.270 ;
        RECT 1629.130 1094.490 1630.310 1095.670 ;
        RECT 1630.730 1094.490 1631.910 1095.670 ;
        RECT 1629.130 916.090 1630.310 917.270 ;
        RECT 1630.730 916.090 1631.910 917.270 ;
        RECT 1629.130 914.490 1630.310 915.670 ;
        RECT 1630.730 914.490 1631.910 915.670 ;
        RECT 1629.130 736.090 1630.310 737.270 ;
        RECT 1630.730 736.090 1631.910 737.270 ;
        RECT 1629.130 734.490 1630.310 735.670 ;
        RECT 1630.730 734.490 1631.910 735.670 ;
        RECT 1629.130 556.090 1630.310 557.270 ;
        RECT 1630.730 556.090 1631.910 557.270 ;
        RECT 1629.130 554.490 1630.310 555.670 ;
        RECT 1630.730 554.490 1631.910 555.670 ;
        RECT 1629.130 376.090 1630.310 377.270 ;
        RECT 1630.730 376.090 1631.910 377.270 ;
        RECT 1629.130 374.490 1630.310 375.670 ;
        RECT 1630.730 374.490 1631.910 375.670 ;
        RECT 1629.130 196.090 1630.310 197.270 ;
        RECT 1630.730 196.090 1631.910 197.270 ;
        RECT 1629.130 194.490 1630.310 195.670 ;
        RECT 1630.730 194.490 1631.910 195.670 ;
        RECT 1629.130 16.090 1630.310 17.270 ;
        RECT 1630.730 16.090 1631.910 17.270 ;
        RECT 1629.130 14.490 1630.310 15.670 ;
        RECT 1630.730 14.490 1631.910 15.670 ;
        RECT 1629.130 -2.910 1630.310 -1.730 ;
        RECT 1630.730 -2.910 1631.910 -1.730 ;
        RECT 1629.130 -4.510 1630.310 -3.330 ;
        RECT 1630.730 -4.510 1631.910 -3.330 ;
        RECT 1809.130 3523.010 1810.310 3524.190 ;
        RECT 1810.730 3523.010 1811.910 3524.190 ;
        RECT 1809.130 3521.410 1810.310 3522.590 ;
        RECT 1810.730 3521.410 1811.910 3522.590 ;
        RECT 1809.130 3436.090 1810.310 3437.270 ;
        RECT 1810.730 3436.090 1811.910 3437.270 ;
        RECT 1809.130 3434.490 1810.310 3435.670 ;
        RECT 1810.730 3434.490 1811.910 3435.670 ;
        RECT 1809.130 3256.090 1810.310 3257.270 ;
        RECT 1810.730 3256.090 1811.910 3257.270 ;
        RECT 1809.130 3254.490 1810.310 3255.670 ;
        RECT 1810.730 3254.490 1811.910 3255.670 ;
        RECT 1809.130 3076.090 1810.310 3077.270 ;
        RECT 1810.730 3076.090 1811.910 3077.270 ;
        RECT 1809.130 3074.490 1810.310 3075.670 ;
        RECT 1810.730 3074.490 1811.910 3075.670 ;
        RECT 1809.130 2896.090 1810.310 2897.270 ;
        RECT 1810.730 2896.090 1811.910 2897.270 ;
        RECT 1809.130 2894.490 1810.310 2895.670 ;
        RECT 1810.730 2894.490 1811.910 2895.670 ;
        RECT 1809.130 2716.090 1810.310 2717.270 ;
        RECT 1810.730 2716.090 1811.910 2717.270 ;
        RECT 1809.130 2714.490 1810.310 2715.670 ;
        RECT 1810.730 2714.490 1811.910 2715.670 ;
        RECT 1809.130 2536.090 1810.310 2537.270 ;
        RECT 1810.730 2536.090 1811.910 2537.270 ;
        RECT 1809.130 2534.490 1810.310 2535.670 ;
        RECT 1810.730 2534.490 1811.910 2535.670 ;
        RECT 1809.130 2356.090 1810.310 2357.270 ;
        RECT 1810.730 2356.090 1811.910 2357.270 ;
        RECT 1809.130 2354.490 1810.310 2355.670 ;
        RECT 1810.730 2354.490 1811.910 2355.670 ;
        RECT 1809.130 2176.090 1810.310 2177.270 ;
        RECT 1810.730 2176.090 1811.910 2177.270 ;
        RECT 1809.130 2174.490 1810.310 2175.670 ;
        RECT 1810.730 2174.490 1811.910 2175.670 ;
        RECT 1809.130 1996.090 1810.310 1997.270 ;
        RECT 1810.730 1996.090 1811.910 1997.270 ;
        RECT 1809.130 1994.490 1810.310 1995.670 ;
        RECT 1810.730 1994.490 1811.910 1995.670 ;
        RECT 1809.130 1816.090 1810.310 1817.270 ;
        RECT 1810.730 1816.090 1811.910 1817.270 ;
        RECT 1809.130 1814.490 1810.310 1815.670 ;
        RECT 1810.730 1814.490 1811.910 1815.670 ;
        RECT 1809.130 1636.090 1810.310 1637.270 ;
        RECT 1810.730 1636.090 1811.910 1637.270 ;
        RECT 1809.130 1634.490 1810.310 1635.670 ;
        RECT 1810.730 1634.490 1811.910 1635.670 ;
        RECT 1809.130 1456.090 1810.310 1457.270 ;
        RECT 1810.730 1456.090 1811.910 1457.270 ;
        RECT 1809.130 1454.490 1810.310 1455.670 ;
        RECT 1810.730 1454.490 1811.910 1455.670 ;
        RECT 1809.130 1276.090 1810.310 1277.270 ;
        RECT 1810.730 1276.090 1811.910 1277.270 ;
        RECT 1809.130 1274.490 1810.310 1275.670 ;
        RECT 1810.730 1274.490 1811.910 1275.670 ;
        RECT 1809.130 1096.090 1810.310 1097.270 ;
        RECT 1810.730 1096.090 1811.910 1097.270 ;
        RECT 1809.130 1094.490 1810.310 1095.670 ;
        RECT 1810.730 1094.490 1811.910 1095.670 ;
        RECT 1809.130 916.090 1810.310 917.270 ;
        RECT 1810.730 916.090 1811.910 917.270 ;
        RECT 1809.130 914.490 1810.310 915.670 ;
        RECT 1810.730 914.490 1811.910 915.670 ;
        RECT 1809.130 736.090 1810.310 737.270 ;
        RECT 1810.730 736.090 1811.910 737.270 ;
        RECT 1809.130 734.490 1810.310 735.670 ;
        RECT 1810.730 734.490 1811.910 735.670 ;
        RECT 1809.130 556.090 1810.310 557.270 ;
        RECT 1810.730 556.090 1811.910 557.270 ;
        RECT 1809.130 554.490 1810.310 555.670 ;
        RECT 1810.730 554.490 1811.910 555.670 ;
        RECT 1809.130 376.090 1810.310 377.270 ;
        RECT 1810.730 376.090 1811.910 377.270 ;
        RECT 1809.130 374.490 1810.310 375.670 ;
        RECT 1810.730 374.490 1811.910 375.670 ;
        RECT 1809.130 196.090 1810.310 197.270 ;
        RECT 1810.730 196.090 1811.910 197.270 ;
        RECT 1809.130 194.490 1810.310 195.670 ;
        RECT 1810.730 194.490 1811.910 195.670 ;
        RECT 1809.130 16.090 1810.310 17.270 ;
        RECT 1810.730 16.090 1811.910 17.270 ;
        RECT 1809.130 14.490 1810.310 15.670 ;
        RECT 1810.730 14.490 1811.910 15.670 ;
        RECT 1809.130 -2.910 1810.310 -1.730 ;
        RECT 1810.730 -2.910 1811.910 -1.730 ;
        RECT 1809.130 -4.510 1810.310 -3.330 ;
        RECT 1810.730 -4.510 1811.910 -3.330 ;
        RECT 1989.130 3523.010 1990.310 3524.190 ;
        RECT 1990.730 3523.010 1991.910 3524.190 ;
        RECT 1989.130 3521.410 1990.310 3522.590 ;
        RECT 1990.730 3521.410 1991.910 3522.590 ;
        RECT 1989.130 3436.090 1990.310 3437.270 ;
        RECT 1990.730 3436.090 1991.910 3437.270 ;
        RECT 1989.130 3434.490 1990.310 3435.670 ;
        RECT 1990.730 3434.490 1991.910 3435.670 ;
        RECT 1989.130 3256.090 1990.310 3257.270 ;
        RECT 1990.730 3256.090 1991.910 3257.270 ;
        RECT 1989.130 3254.490 1990.310 3255.670 ;
        RECT 1990.730 3254.490 1991.910 3255.670 ;
        RECT 1989.130 3076.090 1990.310 3077.270 ;
        RECT 1990.730 3076.090 1991.910 3077.270 ;
        RECT 1989.130 3074.490 1990.310 3075.670 ;
        RECT 1990.730 3074.490 1991.910 3075.670 ;
        RECT 1989.130 2896.090 1990.310 2897.270 ;
        RECT 1990.730 2896.090 1991.910 2897.270 ;
        RECT 1989.130 2894.490 1990.310 2895.670 ;
        RECT 1990.730 2894.490 1991.910 2895.670 ;
        RECT 1989.130 2716.090 1990.310 2717.270 ;
        RECT 1990.730 2716.090 1991.910 2717.270 ;
        RECT 1989.130 2714.490 1990.310 2715.670 ;
        RECT 1990.730 2714.490 1991.910 2715.670 ;
        RECT 1989.130 2536.090 1990.310 2537.270 ;
        RECT 1990.730 2536.090 1991.910 2537.270 ;
        RECT 1989.130 2534.490 1990.310 2535.670 ;
        RECT 1990.730 2534.490 1991.910 2535.670 ;
        RECT 1989.130 2356.090 1990.310 2357.270 ;
        RECT 1990.730 2356.090 1991.910 2357.270 ;
        RECT 1989.130 2354.490 1990.310 2355.670 ;
        RECT 1990.730 2354.490 1991.910 2355.670 ;
        RECT 1989.130 2176.090 1990.310 2177.270 ;
        RECT 1990.730 2176.090 1991.910 2177.270 ;
        RECT 1989.130 2174.490 1990.310 2175.670 ;
        RECT 1990.730 2174.490 1991.910 2175.670 ;
        RECT 1989.130 1996.090 1990.310 1997.270 ;
        RECT 1990.730 1996.090 1991.910 1997.270 ;
        RECT 1989.130 1994.490 1990.310 1995.670 ;
        RECT 1990.730 1994.490 1991.910 1995.670 ;
        RECT 1989.130 1816.090 1990.310 1817.270 ;
        RECT 1990.730 1816.090 1991.910 1817.270 ;
        RECT 1989.130 1814.490 1990.310 1815.670 ;
        RECT 1990.730 1814.490 1991.910 1815.670 ;
        RECT 1989.130 1636.090 1990.310 1637.270 ;
        RECT 1990.730 1636.090 1991.910 1637.270 ;
        RECT 1989.130 1634.490 1990.310 1635.670 ;
        RECT 1990.730 1634.490 1991.910 1635.670 ;
        RECT 1989.130 1456.090 1990.310 1457.270 ;
        RECT 1990.730 1456.090 1991.910 1457.270 ;
        RECT 1989.130 1454.490 1990.310 1455.670 ;
        RECT 1990.730 1454.490 1991.910 1455.670 ;
        RECT 1989.130 1276.090 1990.310 1277.270 ;
        RECT 1990.730 1276.090 1991.910 1277.270 ;
        RECT 1989.130 1274.490 1990.310 1275.670 ;
        RECT 1990.730 1274.490 1991.910 1275.670 ;
        RECT 1989.130 1096.090 1990.310 1097.270 ;
        RECT 1990.730 1096.090 1991.910 1097.270 ;
        RECT 1989.130 1094.490 1990.310 1095.670 ;
        RECT 1990.730 1094.490 1991.910 1095.670 ;
        RECT 1989.130 916.090 1990.310 917.270 ;
        RECT 1990.730 916.090 1991.910 917.270 ;
        RECT 1989.130 914.490 1990.310 915.670 ;
        RECT 1990.730 914.490 1991.910 915.670 ;
        RECT 1989.130 736.090 1990.310 737.270 ;
        RECT 1990.730 736.090 1991.910 737.270 ;
        RECT 1989.130 734.490 1990.310 735.670 ;
        RECT 1990.730 734.490 1991.910 735.670 ;
        RECT 1989.130 556.090 1990.310 557.270 ;
        RECT 1990.730 556.090 1991.910 557.270 ;
        RECT 1989.130 554.490 1990.310 555.670 ;
        RECT 1990.730 554.490 1991.910 555.670 ;
        RECT 1989.130 376.090 1990.310 377.270 ;
        RECT 1990.730 376.090 1991.910 377.270 ;
        RECT 1989.130 374.490 1990.310 375.670 ;
        RECT 1990.730 374.490 1991.910 375.670 ;
        RECT 1989.130 196.090 1990.310 197.270 ;
        RECT 1990.730 196.090 1991.910 197.270 ;
        RECT 1989.130 194.490 1990.310 195.670 ;
        RECT 1990.730 194.490 1991.910 195.670 ;
        RECT 1989.130 16.090 1990.310 17.270 ;
        RECT 1990.730 16.090 1991.910 17.270 ;
        RECT 1989.130 14.490 1990.310 15.670 ;
        RECT 1990.730 14.490 1991.910 15.670 ;
        RECT 1989.130 -2.910 1990.310 -1.730 ;
        RECT 1990.730 -2.910 1991.910 -1.730 ;
        RECT 1989.130 -4.510 1990.310 -3.330 ;
        RECT 1990.730 -4.510 1991.910 -3.330 ;
        RECT 2169.130 3523.010 2170.310 3524.190 ;
        RECT 2170.730 3523.010 2171.910 3524.190 ;
        RECT 2169.130 3521.410 2170.310 3522.590 ;
        RECT 2170.730 3521.410 2171.910 3522.590 ;
        RECT 2169.130 3436.090 2170.310 3437.270 ;
        RECT 2170.730 3436.090 2171.910 3437.270 ;
        RECT 2169.130 3434.490 2170.310 3435.670 ;
        RECT 2170.730 3434.490 2171.910 3435.670 ;
        RECT 2169.130 3256.090 2170.310 3257.270 ;
        RECT 2170.730 3256.090 2171.910 3257.270 ;
        RECT 2169.130 3254.490 2170.310 3255.670 ;
        RECT 2170.730 3254.490 2171.910 3255.670 ;
        RECT 2169.130 3076.090 2170.310 3077.270 ;
        RECT 2170.730 3076.090 2171.910 3077.270 ;
        RECT 2169.130 3074.490 2170.310 3075.670 ;
        RECT 2170.730 3074.490 2171.910 3075.670 ;
        RECT 2169.130 2896.090 2170.310 2897.270 ;
        RECT 2170.730 2896.090 2171.910 2897.270 ;
        RECT 2169.130 2894.490 2170.310 2895.670 ;
        RECT 2170.730 2894.490 2171.910 2895.670 ;
        RECT 2169.130 2716.090 2170.310 2717.270 ;
        RECT 2170.730 2716.090 2171.910 2717.270 ;
        RECT 2169.130 2714.490 2170.310 2715.670 ;
        RECT 2170.730 2714.490 2171.910 2715.670 ;
        RECT 2169.130 2536.090 2170.310 2537.270 ;
        RECT 2170.730 2536.090 2171.910 2537.270 ;
        RECT 2169.130 2534.490 2170.310 2535.670 ;
        RECT 2170.730 2534.490 2171.910 2535.670 ;
        RECT 2169.130 2356.090 2170.310 2357.270 ;
        RECT 2170.730 2356.090 2171.910 2357.270 ;
        RECT 2169.130 2354.490 2170.310 2355.670 ;
        RECT 2170.730 2354.490 2171.910 2355.670 ;
        RECT 2169.130 2176.090 2170.310 2177.270 ;
        RECT 2170.730 2176.090 2171.910 2177.270 ;
        RECT 2169.130 2174.490 2170.310 2175.670 ;
        RECT 2170.730 2174.490 2171.910 2175.670 ;
        RECT 2169.130 1996.090 2170.310 1997.270 ;
        RECT 2170.730 1996.090 2171.910 1997.270 ;
        RECT 2169.130 1994.490 2170.310 1995.670 ;
        RECT 2170.730 1994.490 2171.910 1995.670 ;
        RECT 2169.130 1816.090 2170.310 1817.270 ;
        RECT 2170.730 1816.090 2171.910 1817.270 ;
        RECT 2169.130 1814.490 2170.310 1815.670 ;
        RECT 2170.730 1814.490 2171.910 1815.670 ;
        RECT 2169.130 1636.090 2170.310 1637.270 ;
        RECT 2170.730 1636.090 2171.910 1637.270 ;
        RECT 2169.130 1634.490 2170.310 1635.670 ;
        RECT 2170.730 1634.490 2171.910 1635.670 ;
        RECT 2169.130 1456.090 2170.310 1457.270 ;
        RECT 2170.730 1456.090 2171.910 1457.270 ;
        RECT 2169.130 1454.490 2170.310 1455.670 ;
        RECT 2170.730 1454.490 2171.910 1455.670 ;
        RECT 2169.130 1276.090 2170.310 1277.270 ;
        RECT 2170.730 1276.090 2171.910 1277.270 ;
        RECT 2169.130 1274.490 2170.310 1275.670 ;
        RECT 2170.730 1274.490 2171.910 1275.670 ;
        RECT 2169.130 1096.090 2170.310 1097.270 ;
        RECT 2170.730 1096.090 2171.910 1097.270 ;
        RECT 2169.130 1094.490 2170.310 1095.670 ;
        RECT 2170.730 1094.490 2171.910 1095.670 ;
        RECT 2169.130 916.090 2170.310 917.270 ;
        RECT 2170.730 916.090 2171.910 917.270 ;
        RECT 2169.130 914.490 2170.310 915.670 ;
        RECT 2170.730 914.490 2171.910 915.670 ;
        RECT 2169.130 736.090 2170.310 737.270 ;
        RECT 2170.730 736.090 2171.910 737.270 ;
        RECT 2169.130 734.490 2170.310 735.670 ;
        RECT 2170.730 734.490 2171.910 735.670 ;
        RECT 2169.130 556.090 2170.310 557.270 ;
        RECT 2170.730 556.090 2171.910 557.270 ;
        RECT 2169.130 554.490 2170.310 555.670 ;
        RECT 2170.730 554.490 2171.910 555.670 ;
        RECT 2169.130 376.090 2170.310 377.270 ;
        RECT 2170.730 376.090 2171.910 377.270 ;
        RECT 2169.130 374.490 2170.310 375.670 ;
        RECT 2170.730 374.490 2171.910 375.670 ;
        RECT 2169.130 196.090 2170.310 197.270 ;
        RECT 2170.730 196.090 2171.910 197.270 ;
        RECT 2169.130 194.490 2170.310 195.670 ;
        RECT 2170.730 194.490 2171.910 195.670 ;
        RECT 2169.130 16.090 2170.310 17.270 ;
        RECT 2170.730 16.090 2171.910 17.270 ;
        RECT 2169.130 14.490 2170.310 15.670 ;
        RECT 2170.730 14.490 2171.910 15.670 ;
        RECT 2169.130 -2.910 2170.310 -1.730 ;
        RECT 2170.730 -2.910 2171.910 -1.730 ;
        RECT 2169.130 -4.510 2170.310 -3.330 ;
        RECT 2170.730 -4.510 2171.910 -3.330 ;
        RECT 2349.130 3523.010 2350.310 3524.190 ;
        RECT 2350.730 3523.010 2351.910 3524.190 ;
        RECT 2349.130 3521.410 2350.310 3522.590 ;
        RECT 2350.730 3521.410 2351.910 3522.590 ;
        RECT 2349.130 3436.090 2350.310 3437.270 ;
        RECT 2350.730 3436.090 2351.910 3437.270 ;
        RECT 2349.130 3434.490 2350.310 3435.670 ;
        RECT 2350.730 3434.490 2351.910 3435.670 ;
        RECT 2349.130 3256.090 2350.310 3257.270 ;
        RECT 2350.730 3256.090 2351.910 3257.270 ;
        RECT 2349.130 3254.490 2350.310 3255.670 ;
        RECT 2350.730 3254.490 2351.910 3255.670 ;
        RECT 2349.130 3076.090 2350.310 3077.270 ;
        RECT 2350.730 3076.090 2351.910 3077.270 ;
        RECT 2349.130 3074.490 2350.310 3075.670 ;
        RECT 2350.730 3074.490 2351.910 3075.670 ;
        RECT 2349.130 2896.090 2350.310 2897.270 ;
        RECT 2350.730 2896.090 2351.910 2897.270 ;
        RECT 2349.130 2894.490 2350.310 2895.670 ;
        RECT 2350.730 2894.490 2351.910 2895.670 ;
        RECT 2349.130 2716.090 2350.310 2717.270 ;
        RECT 2350.730 2716.090 2351.910 2717.270 ;
        RECT 2349.130 2714.490 2350.310 2715.670 ;
        RECT 2350.730 2714.490 2351.910 2715.670 ;
        RECT 2349.130 2536.090 2350.310 2537.270 ;
        RECT 2350.730 2536.090 2351.910 2537.270 ;
        RECT 2349.130 2534.490 2350.310 2535.670 ;
        RECT 2350.730 2534.490 2351.910 2535.670 ;
        RECT 2349.130 2356.090 2350.310 2357.270 ;
        RECT 2350.730 2356.090 2351.910 2357.270 ;
        RECT 2349.130 2354.490 2350.310 2355.670 ;
        RECT 2350.730 2354.490 2351.910 2355.670 ;
        RECT 2349.130 2176.090 2350.310 2177.270 ;
        RECT 2350.730 2176.090 2351.910 2177.270 ;
        RECT 2349.130 2174.490 2350.310 2175.670 ;
        RECT 2350.730 2174.490 2351.910 2175.670 ;
        RECT 2349.130 1996.090 2350.310 1997.270 ;
        RECT 2350.730 1996.090 2351.910 1997.270 ;
        RECT 2349.130 1994.490 2350.310 1995.670 ;
        RECT 2350.730 1994.490 2351.910 1995.670 ;
        RECT 2349.130 1816.090 2350.310 1817.270 ;
        RECT 2350.730 1816.090 2351.910 1817.270 ;
        RECT 2349.130 1814.490 2350.310 1815.670 ;
        RECT 2350.730 1814.490 2351.910 1815.670 ;
        RECT 2349.130 1636.090 2350.310 1637.270 ;
        RECT 2350.730 1636.090 2351.910 1637.270 ;
        RECT 2349.130 1634.490 2350.310 1635.670 ;
        RECT 2350.730 1634.490 2351.910 1635.670 ;
        RECT 2349.130 1456.090 2350.310 1457.270 ;
        RECT 2350.730 1456.090 2351.910 1457.270 ;
        RECT 2349.130 1454.490 2350.310 1455.670 ;
        RECT 2350.730 1454.490 2351.910 1455.670 ;
        RECT 2349.130 1276.090 2350.310 1277.270 ;
        RECT 2350.730 1276.090 2351.910 1277.270 ;
        RECT 2349.130 1274.490 2350.310 1275.670 ;
        RECT 2350.730 1274.490 2351.910 1275.670 ;
        RECT 2349.130 1096.090 2350.310 1097.270 ;
        RECT 2350.730 1096.090 2351.910 1097.270 ;
        RECT 2349.130 1094.490 2350.310 1095.670 ;
        RECT 2350.730 1094.490 2351.910 1095.670 ;
        RECT 2349.130 916.090 2350.310 917.270 ;
        RECT 2350.730 916.090 2351.910 917.270 ;
        RECT 2349.130 914.490 2350.310 915.670 ;
        RECT 2350.730 914.490 2351.910 915.670 ;
        RECT 2349.130 736.090 2350.310 737.270 ;
        RECT 2350.730 736.090 2351.910 737.270 ;
        RECT 2349.130 734.490 2350.310 735.670 ;
        RECT 2350.730 734.490 2351.910 735.670 ;
        RECT 2349.130 556.090 2350.310 557.270 ;
        RECT 2350.730 556.090 2351.910 557.270 ;
        RECT 2349.130 554.490 2350.310 555.670 ;
        RECT 2350.730 554.490 2351.910 555.670 ;
        RECT 2349.130 376.090 2350.310 377.270 ;
        RECT 2350.730 376.090 2351.910 377.270 ;
        RECT 2349.130 374.490 2350.310 375.670 ;
        RECT 2350.730 374.490 2351.910 375.670 ;
        RECT 2349.130 196.090 2350.310 197.270 ;
        RECT 2350.730 196.090 2351.910 197.270 ;
        RECT 2349.130 194.490 2350.310 195.670 ;
        RECT 2350.730 194.490 2351.910 195.670 ;
        RECT 2349.130 16.090 2350.310 17.270 ;
        RECT 2350.730 16.090 2351.910 17.270 ;
        RECT 2349.130 14.490 2350.310 15.670 ;
        RECT 2350.730 14.490 2351.910 15.670 ;
        RECT 2349.130 -2.910 2350.310 -1.730 ;
        RECT 2350.730 -2.910 2351.910 -1.730 ;
        RECT 2349.130 -4.510 2350.310 -3.330 ;
        RECT 2350.730 -4.510 2351.910 -3.330 ;
        RECT 2529.130 3523.010 2530.310 3524.190 ;
        RECT 2530.730 3523.010 2531.910 3524.190 ;
        RECT 2529.130 3521.410 2530.310 3522.590 ;
        RECT 2530.730 3521.410 2531.910 3522.590 ;
        RECT 2529.130 3436.090 2530.310 3437.270 ;
        RECT 2530.730 3436.090 2531.910 3437.270 ;
        RECT 2529.130 3434.490 2530.310 3435.670 ;
        RECT 2530.730 3434.490 2531.910 3435.670 ;
        RECT 2529.130 3256.090 2530.310 3257.270 ;
        RECT 2530.730 3256.090 2531.910 3257.270 ;
        RECT 2529.130 3254.490 2530.310 3255.670 ;
        RECT 2530.730 3254.490 2531.910 3255.670 ;
        RECT 2529.130 3076.090 2530.310 3077.270 ;
        RECT 2530.730 3076.090 2531.910 3077.270 ;
        RECT 2529.130 3074.490 2530.310 3075.670 ;
        RECT 2530.730 3074.490 2531.910 3075.670 ;
        RECT 2529.130 2896.090 2530.310 2897.270 ;
        RECT 2530.730 2896.090 2531.910 2897.270 ;
        RECT 2529.130 2894.490 2530.310 2895.670 ;
        RECT 2530.730 2894.490 2531.910 2895.670 ;
        RECT 2529.130 2716.090 2530.310 2717.270 ;
        RECT 2530.730 2716.090 2531.910 2717.270 ;
        RECT 2529.130 2714.490 2530.310 2715.670 ;
        RECT 2530.730 2714.490 2531.910 2715.670 ;
        RECT 2529.130 2536.090 2530.310 2537.270 ;
        RECT 2530.730 2536.090 2531.910 2537.270 ;
        RECT 2529.130 2534.490 2530.310 2535.670 ;
        RECT 2530.730 2534.490 2531.910 2535.670 ;
        RECT 2529.130 2356.090 2530.310 2357.270 ;
        RECT 2530.730 2356.090 2531.910 2357.270 ;
        RECT 2529.130 2354.490 2530.310 2355.670 ;
        RECT 2530.730 2354.490 2531.910 2355.670 ;
        RECT 2529.130 2176.090 2530.310 2177.270 ;
        RECT 2530.730 2176.090 2531.910 2177.270 ;
        RECT 2529.130 2174.490 2530.310 2175.670 ;
        RECT 2530.730 2174.490 2531.910 2175.670 ;
        RECT 2529.130 1996.090 2530.310 1997.270 ;
        RECT 2530.730 1996.090 2531.910 1997.270 ;
        RECT 2529.130 1994.490 2530.310 1995.670 ;
        RECT 2530.730 1994.490 2531.910 1995.670 ;
        RECT 2529.130 1816.090 2530.310 1817.270 ;
        RECT 2530.730 1816.090 2531.910 1817.270 ;
        RECT 2529.130 1814.490 2530.310 1815.670 ;
        RECT 2530.730 1814.490 2531.910 1815.670 ;
        RECT 2529.130 1636.090 2530.310 1637.270 ;
        RECT 2530.730 1636.090 2531.910 1637.270 ;
        RECT 2529.130 1634.490 2530.310 1635.670 ;
        RECT 2530.730 1634.490 2531.910 1635.670 ;
        RECT 2529.130 1456.090 2530.310 1457.270 ;
        RECT 2530.730 1456.090 2531.910 1457.270 ;
        RECT 2529.130 1454.490 2530.310 1455.670 ;
        RECT 2530.730 1454.490 2531.910 1455.670 ;
        RECT 2529.130 1276.090 2530.310 1277.270 ;
        RECT 2530.730 1276.090 2531.910 1277.270 ;
        RECT 2529.130 1274.490 2530.310 1275.670 ;
        RECT 2530.730 1274.490 2531.910 1275.670 ;
        RECT 2529.130 1096.090 2530.310 1097.270 ;
        RECT 2530.730 1096.090 2531.910 1097.270 ;
        RECT 2529.130 1094.490 2530.310 1095.670 ;
        RECT 2530.730 1094.490 2531.910 1095.670 ;
        RECT 2529.130 916.090 2530.310 917.270 ;
        RECT 2530.730 916.090 2531.910 917.270 ;
        RECT 2529.130 914.490 2530.310 915.670 ;
        RECT 2530.730 914.490 2531.910 915.670 ;
        RECT 2529.130 736.090 2530.310 737.270 ;
        RECT 2530.730 736.090 2531.910 737.270 ;
        RECT 2529.130 734.490 2530.310 735.670 ;
        RECT 2530.730 734.490 2531.910 735.670 ;
        RECT 2529.130 556.090 2530.310 557.270 ;
        RECT 2530.730 556.090 2531.910 557.270 ;
        RECT 2529.130 554.490 2530.310 555.670 ;
        RECT 2530.730 554.490 2531.910 555.670 ;
        RECT 2529.130 376.090 2530.310 377.270 ;
        RECT 2530.730 376.090 2531.910 377.270 ;
        RECT 2529.130 374.490 2530.310 375.670 ;
        RECT 2530.730 374.490 2531.910 375.670 ;
        RECT 2529.130 196.090 2530.310 197.270 ;
        RECT 2530.730 196.090 2531.910 197.270 ;
        RECT 2529.130 194.490 2530.310 195.670 ;
        RECT 2530.730 194.490 2531.910 195.670 ;
        RECT 2529.130 16.090 2530.310 17.270 ;
        RECT 2530.730 16.090 2531.910 17.270 ;
        RECT 2529.130 14.490 2530.310 15.670 ;
        RECT 2530.730 14.490 2531.910 15.670 ;
        RECT 2529.130 -2.910 2530.310 -1.730 ;
        RECT 2530.730 -2.910 2531.910 -1.730 ;
        RECT 2529.130 -4.510 2530.310 -3.330 ;
        RECT 2530.730 -4.510 2531.910 -3.330 ;
        RECT 2709.130 3523.010 2710.310 3524.190 ;
        RECT 2710.730 3523.010 2711.910 3524.190 ;
        RECT 2709.130 3521.410 2710.310 3522.590 ;
        RECT 2710.730 3521.410 2711.910 3522.590 ;
        RECT 2709.130 3436.090 2710.310 3437.270 ;
        RECT 2710.730 3436.090 2711.910 3437.270 ;
        RECT 2709.130 3434.490 2710.310 3435.670 ;
        RECT 2710.730 3434.490 2711.910 3435.670 ;
        RECT 2709.130 3256.090 2710.310 3257.270 ;
        RECT 2710.730 3256.090 2711.910 3257.270 ;
        RECT 2709.130 3254.490 2710.310 3255.670 ;
        RECT 2710.730 3254.490 2711.910 3255.670 ;
        RECT 2709.130 3076.090 2710.310 3077.270 ;
        RECT 2710.730 3076.090 2711.910 3077.270 ;
        RECT 2709.130 3074.490 2710.310 3075.670 ;
        RECT 2710.730 3074.490 2711.910 3075.670 ;
        RECT 2709.130 2896.090 2710.310 2897.270 ;
        RECT 2710.730 2896.090 2711.910 2897.270 ;
        RECT 2709.130 2894.490 2710.310 2895.670 ;
        RECT 2710.730 2894.490 2711.910 2895.670 ;
        RECT 2709.130 2716.090 2710.310 2717.270 ;
        RECT 2710.730 2716.090 2711.910 2717.270 ;
        RECT 2709.130 2714.490 2710.310 2715.670 ;
        RECT 2710.730 2714.490 2711.910 2715.670 ;
        RECT 2709.130 2536.090 2710.310 2537.270 ;
        RECT 2710.730 2536.090 2711.910 2537.270 ;
        RECT 2709.130 2534.490 2710.310 2535.670 ;
        RECT 2710.730 2534.490 2711.910 2535.670 ;
        RECT 2709.130 2356.090 2710.310 2357.270 ;
        RECT 2710.730 2356.090 2711.910 2357.270 ;
        RECT 2709.130 2354.490 2710.310 2355.670 ;
        RECT 2710.730 2354.490 2711.910 2355.670 ;
        RECT 2709.130 2176.090 2710.310 2177.270 ;
        RECT 2710.730 2176.090 2711.910 2177.270 ;
        RECT 2709.130 2174.490 2710.310 2175.670 ;
        RECT 2710.730 2174.490 2711.910 2175.670 ;
        RECT 2709.130 1996.090 2710.310 1997.270 ;
        RECT 2710.730 1996.090 2711.910 1997.270 ;
        RECT 2709.130 1994.490 2710.310 1995.670 ;
        RECT 2710.730 1994.490 2711.910 1995.670 ;
        RECT 2709.130 1816.090 2710.310 1817.270 ;
        RECT 2710.730 1816.090 2711.910 1817.270 ;
        RECT 2709.130 1814.490 2710.310 1815.670 ;
        RECT 2710.730 1814.490 2711.910 1815.670 ;
        RECT 2709.130 1636.090 2710.310 1637.270 ;
        RECT 2710.730 1636.090 2711.910 1637.270 ;
        RECT 2709.130 1634.490 2710.310 1635.670 ;
        RECT 2710.730 1634.490 2711.910 1635.670 ;
        RECT 2709.130 1456.090 2710.310 1457.270 ;
        RECT 2710.730 1456.090 2711.910 1457.270 ;
        RECT 2709.130 1454.490 2710.310 1455.670 ;
        RECT 2710.730 1454.490 2711.910 1455.670 ;
        RECT 2709.130 1276.090 2710.310 1277.270 ;
        RECT 2710.730 1276.090 2711.910 1277.270 ;
        RECT 2709.130 1274.490 2710.310 1275.670 ;
        RECT 2710.730 1274.490 2711.910 1275.670 ;
        RECT 2709.130 1096.090 2710.310 1097.270 ;
        RECT 2710.730 1096.090 2711.910 1097.270 ;
        RECT 2709.130 1094.490 2710.310 1095.670 ;
        RECT 2710.730 1094.490 2711.910 1095.670 ;
        RECT 2709.130 916.090 2710.310 917.270 ;
        RECT 2710.730 916.090 2711.910 917.270 ;
        RECT 2709.130 914.490 2710.310 915.670 ;
        RECT 2710.730 914.490 2711.910 915.670 ;
        RECT 2709.130 736.090 2710.310 737.270 ;
        RECT 2710.730 736.090 2711.910 737.270 ;
        RECT 2709.130 734.490 2710.310 735.670 ;
        RECT 2710.730 734.490 2711.910 735.670 ;
        RECT 2709.130 556.090 2710.310 557.270 ;
        RECT 2710.730 556.090 2711.910 557.270 ;
        RECT 2709.130 554.490 2710.310 555.670 ;
        RECT 2710.730 554.490 2711.910 555.670 ;
        RECT 2709.130 376.090 2710.310 377.270 ;
        RECT 2710.730 376.090 2711.910 377.270 ;
        RECT 2709.130 374.490 2710.310 375.670 ;
        RECT 2710.730 374.490 2711.910 375.670 ;
        RECT 2709.130 196.090 2710.310 197.270 ;
        RECT 2710.730 196.090 2711.910 197.270 ;
        RECT 2709.130 194.490 2710.310 195.670 ;
        RECT 2710.730 194.490 2711.910 195.670 ;
        RECT 2709.130 16.090 2710.310 17.270 ;
        RECT 2710.730 16.090 2711.910 17.270 ;
        RECT 2709.130 14.490 2710.310 15.670 ;
        RECT 2710.730 14.490 2711.910 15.670 ;
        RECT 2709.130 -2.910 2710.310 -1.730 ;
        RECT 2710.730 -2.910 2711.910 -1.730 ;
        RECT 2709.130 -4.510 2710.310 -3.330 ;
        RECT 2710.730 -4.510 2711.910 -3.330 ;
        RECT 2889.130 3523.010 2890.310 3524.190 ;
        RECT 2890.730 3523.010 2891.910 3524.190 ;
        RECT 2889.130 3521.410 2890.310 3522.590 ;
        RECT 2890.730 3521.410 2891.910 3522.590 ;
        RECT 2889.130 3436.090 2890.310 3437.270 ;
        RECT 2890.730 3436.090 2891.910 3437.270 ;
        RECT 2889.130 3434.490 2890.310 3435.670 ;
        RECT 2890.730 3434.490 2891.910 3435.670 ;
        RECT 2889.130 3256.090 2890.310 3257.270 ;
        RECT 2890.730 3256.090 2891.910 3257.270 ;
        RECT 2889.130 3254.490 2890.310 3255.670 ;
        RECT 2890.730 3254.490 2891.910 3255.670 ;
        RECT 2889.130 3076.090 2890.310 3077.270 ;
        RECT 2890.730 3076.090 2891.910 3077.270 ;
        RECT 2889.130 3074.490 2890.310 3075.670 ;
        RECT 2890.730 3074.490 2891.910 3075.670 ;
        RECT 2889.130 2896.090 2890.310 2897.270 ;
        RECT 2890.730 2896.090 2891.910 2897.270 ;
        RECT 2889.130 2894.490 2890.310 2895.670 ;
        RECT 2890.730 2894.490 2891.910 2895.670 ;
        RECT 2889.130 2716.090 2890.310 2717.270 ;
        RECT 2890.730 2716.090 2891.910 2717.270 ;
        RECT 2889.130 2714.490 2890.310 2715.670 ;
        RECT 2890.730 2714.490 2891.910 2715.670 ;
        RECT 2889.130 2536.090 2890.310 2537.270 ;
        RECT 2890.730 2536.090 2891.910 2537.270 ;
        RECT 2889.130 2534.490 2890.310 2535.670 ;
        RECT 2890.730 2534.490 2891.910 2535.670 ;
        RECT 2889.130 2356.090 2890.310 2357.270 ;
        RECT 2890.730 2356.090 2891.910 2357.270 ;
        RECT 2889.130 2354.490 2890.310 2355.670 ;
        RECT 2890.730 2354.490 2891.910 2355.670 ;
        RECT 2889.130 2176.090 2890.310 2177.270 ;
        RECT 2890.730 2176.090 2891.910 2177.270 ;
        RECT 2889.130 2174.490 2890.310 2175.670 ;
        RECT 2890.730 2174.490 2891.910 2175.670 ;
        RECT 2889.130 1996.090 2890.310 1997.270 ;
        RECT 2890.730 1996.090 2891.910 1997.270 ;
        RECT 2889.130 1994.490 2890.310 1995.670 ;
        RECT 2890.730 1994.490 2891.910 1995.670 ;
        RECT 2889.130 1816.090 2890.310 1817.270 ;
        RECT 2890.730 1816.090 2891.910 1817.270 ;
        RECT 2889.130 1814.490 2890.310 1815.670 ;
        RECT 2890.730 1814.490 2891.910 1815.670 ;
        RECT 2889.130 1636.090 2890.310 1637.270 ;
        RECT 2890.730 1636.090 2891.910 1637.270 ;
        RECT 2889.130 1634.490 2890.310 1635.670 ;
        RECT 2890.730 1634.490 2891.910 1635.670 ;
        RECT 2889.130 1456.090 2890.310 1457.270 ;
        RECT 2890.730 1456.090 2891.910 1457.270 ;
        RECT 2889.130 1454.490 2890.310 1455.670 ;
        RECT 2890.730 1454.490 2891.910 1455.670 ;
        RECT 2889.130 1276.090 2890.310 1277.270 ;
        RECT 2890.730 1276.090 2891.910 1277.270 ;
        RECT 2889.130 1274.490 2890.310 1275.670 ;
        RECT 2890.730 1274.490 2891.910 1275.670 ;
        RECT 2889.130 1096.090 2890.310 1097.270 ;
        RECT 2890.730 1096.090 2891.910 1097.270 ;
        RECT 2889.130 1094.490 2890.310 1095.670 ;
        RECT 2890.730 1094.490 2891.910 1095.670 ;
        RECT 2889.130 916.090 2890.310 917.270 ;
        RECT 2890.730 916.090 2891.910 917.270 ;
        RECT 2889.130 914.490 2890.310 915.670 ;
        RECT 2890.730 914.490 2891.910 915.670 ;
        RECT 2889.130 736.090 2890.310 737.270 ;
        RECT 2890.730 736.090 2891.910 737.270 ;
        RECT 2889.130 734.490 2890.310 735.670 ;
        RECT 2890.730 734.490 2891.910 735.670 ;
        RECT 2889.130 556.090 2890.310 557.270 ;
        RECT 2890.730 556.090 2891.910 557.270 ;
        RECT 2889.130 554.490 2890.310 555.670 ;
        RECT 2890.730 554.490 2891.910 555.670 ;
        RECT 2889.130 376.090 2890.310 377.270 ;
        RECT 2890.730 376.090 2891.910 377.270 ;
        RECT 2889.130 374.490 2890.310 375.670 ;
        RECT 2890.730 374.490 2891.910 375.670 ;
        RECT 2889.130 196.090 2890.310 197.270 ;
        RECT 2890.730 196.090 2891.910 197.270 ;
        RECT 2889.130 194.490 2890.310 195.670 ;
        RECT 2890.730 194.490 2891.910 195.670 ;
        RECT 2889.130 16.090 2890.310 17.270 ;
        RECT 2890.730 16.090 2891.910 17.270 ;
        RECT 2889.130 14.490 2890.310 15.670 ;
        RECT 2890.730 14.490 2891.910 15.670 ;
        RECT 2889.130 -2.910 2890.310 -1.730 ;
        RECT 2890.730 -2.910 2891.910 -1.730 ;
        RECT 2889.130 -4.510 2890.310 -3.330 ;
        RECT 2890.730 -4.510 2891.910 -3.330 ;
        RECT 2926.710 3523.010 2927.890 3524.190 ;
        RECT 2928.310 3523.010 2929.490 3524.190 ;
        RECT 2926.710 3521.410 2927.890 3522.590 ;
        RECT 2928.310 3521.410 2929.490 3522.590 ;
        RECT 2926.710 3436.090 2927.890 3437.270 ;
        RECT 2928.310 3436.090 2929.490 3437.270 ;
        RECT 2926.710 3434.490 2927.890 3435.670 ;
        RECT 2928.310 3434.490 2929.490 3435.670 ;
        RECT 2926.710 3256.090 2927.890 3257.270 ;
        RECT 2928.310 3256.090 2929.490 3257.270 ;
        RECT 2926.710 3254.490 2927.890 3255.670 ;
        RECT 2928.310 3254.490 2929.490 3255.670 ;
        RECT 2926.710 3076.090 2927.890 3077.270 ;
        RECT 2928.310 3076.090 2929.490 3077.270 ;
        RECT 2926.710 3074.490 2927.890 3075.670 ;
        RECT 2928.310 3074.490 2929.490 3075.670 ;
        RECT 2926.710 2896.090 2927.890 2897.270 ;
        RECT 2928.310 2896.090 2929.490 2897.270 ;
        RECT 2926.710 2894.490 2927.890 2895.670 ;
        RECT 2928.310 2894.490 2929.490 2895.670 ;
        RECT 2926.710 2716.090 2927.890 2717.270 ;
        RECT 2928.310 2716.090 2929.490 2717.270 ;
        RECT 2926.710 2714.490 2927.890 2715.670 ;
        RECT 2928.310 2714.490 2929.490 2715.670 ;
        RECT 2926.710 2536.090 2927.890 2537.270 ;
        RECT 2928.310 2536.090 2929.490 2537.270 ;
        RECT 2926.710 2534.490 2927.890 2535.670 ;
        RECT 2928.310 2534.490 2929.490 2535.670 ;
        RECT 2926.710 2356.090 2927.890 2357.270 ;
        RECT 2928.310 2356.090 2929.490 2357.270 ;
        RECT 2926.710 2354.490 2927.890 2355.670 ;
        RECT 2928.310 2354.490 2929.490 2355.670 ;
        RECT 2926.710 2176.090 2927.890 2177.270 ;
        RECT 2928.310 2176.090 2929.490 2177.270 ;
        RECT 2926.710 2174.490 2927.890 2175.670 ;
        RECT 2928.310 2174.490 2929.490 2175.670 ;
        RECT 2926.710 1996.090 2927.890 1997.270 ;
        RECT 2928.310 1996.090 2929.490 1997.270 ;
        RECT 2926.710 1994.490 2927.890 1995.670 ;
        RECT 2928.310 1994.490 2929.490 1995.670 ;
        RECT 2926.710 1816.090 2927.890 1817.270 ;
        RECT 2928.310 1816.090 2929.490 1817.270 ;
        RECT 2926.710 1814.490 2927.890 1815.670 ;
        RECT 2928.310 1814.490 2929.490 1815.670 ;
        RECT 2926.710 1636.090 2927.890 1637.270 ;
        RECT 2928.310 1636.090 2929.490 1637.270 ;
        RECT 2926.710 1634.490 2927.890 1635.670 ;
        RECT 2928.310 1634.490 2929.490 1635.670 ;
        RECT 2926.710 1456.090 2927.890 1457.270 ;
        RECT 2928.310 1456.090 2929.490 1457.270 ;
        RECT 2926.710 1454.490 2927.890 1455.670 ;
        RECT 2928.310 1454.490 2929.490 1455.670 ;
        RECT 2926.710 1276.090 2927.890 1277.270 ;
        RECT 2928.310 1276.090 2929.490 1277.270 ;
        RECT 2926.710 1274.490 2927.890 1275.670 ;
        RECT 2928.310 1274.490 2929.490 1275.670 ;
        RECT 2926.710 1096.090 2927.890 1097.270 ;
        RECT 2928.310 1096.090 2929.490 1097.270 ;
        RECT 2926.710 1094.490 2927.890 1095.670 ;
        RECT 2928.310 1094.490 2929.490 1095.670 ;
        RECT 2926.710 916.090 2927.890 917.270 ;
        RECT 2928.310 916.090 2929.490 917.270 ;
        RECT 2926.710 914.490 2927.890 915.670 ;
        RECT 2928.310 914.490 2929.490 915.670 ;
        RECT 2926.710 736.090 2927.890 737.270 ;
        RECT 2928.310 736.090 2929.490 737.270 ;
        RECT 2926.710 734.490 2927.890 735.670 ;
        RECT 2928.310 734.490 2929.490 735.670 ;
        RECT 2926.710 556.090 2927.890 557.270 ;
        RECT 2928.310 556.090 2929.490 557.270 ;
        RECT 2926.710 554.490 2927.890 555.670 ;
        RECT 2928.310 554.490 2929.490 555.670 ;
        RECT 2926.710 376.090 2927.890 377.270 ;
        RECT 2928.310 376.090 2929.490 377.270 ;
        RECT 2926.710 374.490 2927.890 375.670 ;
        RECT 2928.310 374.490 2929.490 375.670 ;
        RECT 2926.710 196.090 2927.890 197.270 ;
        RECT 2928.310 196.090 2929.490 197.270 ;
        RECT 2926.710 194.490 2927.890 195.670 ;
        RECT 2928.310 194.490 2929.490 195.670 ;
        RECT 2926.710 16.090 2927.890 17.270 ;
        RECT 2928.310 16.090 2929.490 17.270 ;
        RECT 2926.710 14.490 2927.890 15.670 ;
        RECT 2928.310 14.490 2929.490 15.670 ;
        RECT 2926.710 -2.910 2927.890 -1.730 ;
        RECT 2928.310 -2.910 2929.490 -1.730 ;
        RECT 2926.710 -4.510 2927.890 -3.330 ;
        RECT 2928.310 -4.510 2929.490 -3.330 ;
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
        RECT -14.830 3434.330 2934.450 3437.430 ;
        RECT -14.830 3254.330 2934.450 3257.430 ;
        RECT -14.830 3074.330 2934.450 3077.430 ;
        RECT -14.830 2894.330 2934.450 2897.430 ;
        RECT -14.830 2714.330 2934.450 2717.430 ;
        RECT -14.830 2534.330 2934.450 2537.430 ;
        RECT -14.830 2354.330 2934.450 2357.430 ;
        RECT -14.830 2174.330 2934.450 2177.430 ;
        RECT -14.830 1994.330 2934.450 1997.430 ;
        RECT -14.830 1814.330 2934.450 1817.430 ;
        RECT -14.830 1634.330 2934.450 1637.430 ;
        RECT -14.830 1454.330 2934.450 1457.430 ;
        RECT -14.830 1274.330 2934.450 1277.430 ;
        RECT -14.830 1094.330 2934.450 1097.430 ;
        RECT -14.830 914.330 2934.450 917.430 ;
        RECT -14.830 734.330 2934.450 737.430 ;
        RECT -14.830 554.330 2934.450 557.430 ;
        RECT -14.830 374.330 2934.450 377.430 ;
        RECT -14.830 194.330 2934.450 197.430 ;
        RECT -14.830 14.330 2934.450 17.430 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
        RECT 207.570 1010.000 210.670 3538.750 ;
        RECT 387.570 1010.000 390.670 3538.750 ;
        RECT 567.570 1010.000 570.670 3538.750 ;
        RECT 747.570 1010.000 750.670 3538.750 ;
        RECT 927.570 1010.000 930.670 3538.750 ;
        RECT 1107.570 1010.000 1110.670 3538.750 ;
        RECT 207.570 -19.070 210.670 390.000 ;
        RECT 387.570 -19.070 390.670 390.000 ;
        RECT 567.570 -19.070 570.670 390.000 ;
        RECT 747.570 -19.070 750.670 390.000 ;
        RECT 927.570 -19.070 930.670 390.000 ;
        RECT 1107.570 -19.070 1110.670 390.000 ;
        RECT 1287.570 -19.070 1290.670 3538.750 ;
        RECT 1467.570 -19.070 1470.670 3538.750 ;
        RECT 1647.570 -19.070 1650.670 3538.750 ;
        RECT 1827.570 -19.070 1830.670 3538.750 ;
        RECT 2007.570 -19.070 2010.670 3538.750 ;
        RECT 2187.570 -19.070 2190.670 3538.750 ;
        RECT 2367.570 -19.070 2370.670 3538.750 ;
        RECT 2547.570 -19.070 2550.670 3538.750 ;
        RECT 2727.570 -19.070 2730.670 3538.750 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
      LAYER via4 ;
        RECT -19.470 3532.610 -18.290 3533.790 ;
        RECT -17.870 3532.610 -16.690 3533.790 ;
        RECT -19.470 3531.010 -18.290 3532.190 ;
        RECT -17.870 3531.010 -16.690 3532.190 ;
        RECT -19.470 3454.690 -18.290 3455.870 ;
        RECT -17.870 3454.690 -16.690 3455.870 ;
        RECT -19.470 3453.090 -18.290 3454.270 ;
        RECT -17.870 3453.090 -16.690 3454.270 ;
        RECT -19.470 3274.690 -18.290 3275.870 ;
        RECT -17.870 3274.690 -16.690 3275.870 ;
        RECT -19.470 3273.090 -18.290 3274.270 ;
        RECT -17.870 3273.090 -16.690 3274.270 ;
        RECT -19.470 3094.690 -18.290 3095.870 ;
        RECT -17.870 3094.690 -16.690 3095.870 ;
        RECT -19.470 3093.090 -18.290 3094.270 ;
        RECT -17.870 3093.090 -16.690 3094.270 ;
        RECT -19.470 2914.690 -18.290 2915.870 ;
        RECT -17.870 2914.690 -16.690 2915.870 ;
        RECT -19.470 2913.090 -18.290 2914.270 ;
        RECT -17.870 2913.090 -16.690 2914.270 ;
        RECT -19.470 2734.690 -18.290 2735.870 ;
        RECT -17.870 2734.690 -16.690 2735.870 ;
        RECT -19.470 2733.090 -18.290 2734.270 ;
        RECT -17.870 2733.090 -16.690 2734.270 ;
        RECT -19.470 2554.690 -18.290 2555.870 ;
        RECT -17.870 2554.690 -16.690 2555.870 ;
        RECT -19.470 2553.090 -18.290 2554.270 ;
        RECT -17.870 2553.090 -16.690 2554.270 ;
        RECT -19.470 2374.690 -18.290 2375.870 ;
        RECT -17.870 2374.690 -16.690 2375.870 ;
        RECT -19.470 2373.090 -18.290 2374.270 ;
        RECT -17.870 2373.090 -16.690 2374.270 ;
        RECT -19.470 2194.690 -18.290 2195.870 ;
        RECT -17.870 2194.690 -16.690 2195.870 ;
        RECT -19.470 2193.090 -18.290 2194.270 ;
        RECT -17.870 2193.090 -16.690 2194.270 ;
        RECT -19.470 2014.690 -18.290 2015.870 ;
        RECT -17.870 2014.690 -16.690 2015.870 ;
        RECT -19.470 2013.090 -18.290 2014.270 ;
        RECT -17.870 2013.090 -16.690 2014.270 ;
        RECT -19.470 1834.690 -18.290 1835.870 ;
        RECT -17.870 1834.690 -16.690 1835.870 ;
        RECT -19.470 1833.090 -18.290 1834.270 ;
        RECT -17.870 1833.090 -16.690 1834.270 ;
        RECT -19.470 1654.690 -18.290 1655.870 ;
        RECT -17.870 1654.690 -16.690 1655.870 ;
        RECT -19.470 1653.090 -18.290 1654.270 ;
        RECT -17.870 1653.090 -16.690 1654.270 ;
        RECT -19.470 1474.690 -18.290 1475.870 ;
        RECT -17.870 1474.690 -16.690 1475.870 ;
        RECT -19.470 1473.090 -18.290 1474.270 ;
        RECT -17.870 1473.090 -16.690 1474.270 ;
        RECT -19.470 1294.690 -18.290 1295.870 ;
        RECT -17.870 1294.690 -16.690 1295.870 ;
        RECT -19.470 1293.090 -18.290 1294.270 ;
        RECT -17.870 1293.090 -16.690 1294.270 ;
        RECT -19.470 1114.690 -18.290 1115.870 ;
        RECT -17.870 1114.690 -16.690 1115.870 ;
        RECT -19.470 1113.090 -18.290 1114.270 ;
        RECT -17.870 1113.090 -16.690 1114.270 ;
        RECT -19.470 934.690 -18.290 935.870 ;
        RECT -17.870 934.690 -16.690 935.870 ;
        RECT -19.470 933.090 -18.290 934.270 ;
        RECT -17.870 933.090 -16.690 934.270 ;
        RECT -19.470 754.690 -18.290 755.870 ;
        RECT -17.870 754.690 -16.690 755.870 ;
        RECT -19.470 753.090 -18.290 754.270 ;
        RECT -17.870 753.090 -16.690 754.270 ;
        RECT -19.470 574.690 -18.290 575.870 ;
        RECT -17.870 574.690 -16.690 575.870 ;
        RECT -19.470 573.090 -18.290 574.270 ;
        RECT -17.870 573.090 -16.690 574.270 ;
        RECT -19.470 394.690 -18.290 395.870 ;
        RECT -17.870 394.690 -16.690 395.870 ;
        RECT -19.470 393.090 -18.290 394.270 ;
        RECT -17.870 393.090 -16.690 394.270 ;
        RECT -19.470 214.690 -18.290 215.870 ;
        RECT -17.870 214.690 -16.690 215.870 ;
        RECT -19.470 213.090 -18.290 214.270 ;
        RECT -17.870 213.090 -16.690 214.270 ;
        RECT -19.470 34.690 -18.290 35.870 ;
        RECT -17.870 34.690 -16.690 35.870 ;
        RECT -19.470 33.090 -18.290 34.270 ;
        RECT -17.870 33.090 -16.690 34.270 ;
        RECT -19.470 -12.510 -18.290 -11.330 ;
        RECT -17.870 -12.510 -16.690 -11.330 ;
        RECT -19.470 -14.110 -18.290 -12.930 ;
        RECT -17.870 -14.110 -16.690 -12.930 ;
        RECT 27.730 3532.610 28.910 3533.790 ;
        RECT 29.330 3532.610 30.510 3533.790 ;
        RECT 27.730 3531.010 28.910 3532.190 ;
        RECT 29.330 3531.010 30.510 3532.190 ;
        RECT 27.730 3454.690 28.910 3455.870 ;
        RECT 29.330 3454.690 30.510 3455.870 ;
        RECT 27.730 3453.090 28.910 3454.270 ;
        RECT 29.330 3453.090 30.510 3454.270 ;
        RECT 27.730 3274.690 28.910 3275.870 ;
        RECT 29.330 3274.690 30.510 3275.870 ;
        RECT 27.730 3273.090 28.910 3274.270 ;
        RECT 29.330 3273.090 30.510 3274.270 ;
        RECT 27.730 3094.690 28.910 3095.870 ;
        RECT 29.330 3094.690 30.510 3095.870 ;
        RECT 27.730 3093.090 28.910 3094.270 ;
        RECT 29.330 3093.090 30.510 3094.270 ;
        RECT 27.730 2914.690 28.910 2915.870 ;
        RECT 29.330 2914.690 30.510 2915.870 ;
        RECT 27.730 2913.090 28.910 2914.270 ;
        RECT 29.330 2913.090 30.510 2914.270 ;
        RECT 27.730 2734.690 28.910 2735.870 ;
        RECT 29.330 2734.690 30.510 2735.870 ;
        RECT 27.730 2733.090 28.910 2734.270 ;
        RECT 29.330 2733.090 30.510 2734.270 ;
        RECT 27.730 2554.690 28.910 2555.870 ;
        RECT 29.330 2554.690 30.510 2555.870 ;
        RECT 27.730 2553.090 28.910 2554.270 ;
        RECT 29.330 2553.090 30.510 2554.270 ;
        RECT 27.730 2374.690 28.910 2375.870 ;
        RECT 29.330 2374.690 30.510 2375.870 ;
        RECT 27.730 2373.090 28.910 2374.270 ;
        RECT 29.330 2373.090 30.510 2374.270 ;
        RECT 27.730 2194.690 28.910 2195.870 ;
        RECT 29.330 2194.690 30.510 2195.870 ;
        RECT 27.730 2193.090 28.910 2194.270 ;
        RECT 29.330 2193.090 30.510 2194.270 ;
        RECT 27.730 2014.690 28.910 2015.870 ;
        RECT 29.330 2014.690 30.510 2015.870 ;
        RECT 27.730 2013.090 28.910 2014.270 ;
        RECT 29.330 2013.090 30.510 2014.270 ;
        RECT 27.730 1834.690 28.910 1835.870 ;
        RECT 29.330 1834.690 30.510 1835.870 ;
        RECT 27.730 1833.090 28.910 1834.270 ;
        RECT 29.330 1833.090 30.510 1834.270 ;
        RECT 27.730 1654.690 28.910 1655.870 ;
        RECT 29.330 1654.690 30.510 1655.870 ;
        RECT 27.730 1653.090 28.910 1654.270 ;
        RECT 29.330 1653.090 30.510 1654.270 ;
        RECT 27.730 1474.690 28.910 1475.870 ;
        RECT 29.330 1474.690 30.510 1475.870 ;
        RECT 27.730 1473.090 28.910 1474.270 ;
        RECT 29.330 1473.090 30.510 1474.270 ;
        RECT 27.730 1294.690 28.910 1295.870 ;
        RECT 29.330 1294.690 30.510 1295.870 ;
        RECT 27.730 1293.090 28.910 1294.270 ;
        RECT 29.330 1293.090 30.510 1294.270 ;
        RECT 27.730 1114.690 28.910 1115.870 ;
        RECT 29.330 1114.690 30.510 1115.870 ;
        RECT 27.730 1113.090 28.910 1114.270 ;
        RECT 29.330 1113.090 30.510 1114.270 ;
        RECT 207.730 3532.610 208.910 3533.790 ;
        RECT 209.330 3532.610 210.510 3533.790 ;
        RECT 207.730 3531.010 208.910 3532.190 ;
        RECT 209.330 3531.010 210.510 3532.190 ;
        RECT 207.730 3454.690 208.910 3455.870 ;
        RECT 209.330 3454.690 210.510 3455.870 ;
        RECT 207.730 3453.090 208.910 3454.270 ;
        RECT 209.330 3453.090 210.510 3454.270 ;
        RECT 207.730 3274.690 208.910 3275.870 ;
        RECT 209.330 3274.690 210.510 3275.870 ;
        RECT 207.730 3273.090 208.910 3274.270 ;
        RECT 209.330 3273.090 210.510 3274.270 ;
        RECT 207.730 3094.690 208.910 3095.870 ;
        RECT 209.330 3094.690 210.510 3095.870 ;
        RECT 207.730 3093.090 208.910 3094.270 ;
        RECT 209.330 3093.090 210.510 3094.270 ;
        RECT 207.730 2914.690 208.910 2915.870 ;
        RECT 209.330 2914.690 210.510 2915.870 ;
        RECT 207.730 2913.090 208.910 2914.270 ;
        RECT 209.330 2913.090 210.510 2914.270 ;
        RECT 207.730 2734.690 208.910 2735.870 ;
        RECT 209.330 2734.690 210.510 2735.870 ;
        RECT 207.730 2733.090 208.910 2734.270 ;
        RECT 209.330 2733.090 210.510 2734.270 ;
        RECT 207.730 2554.690 208.910 2555.870 ;
        RECT 209.330 2554.690 210.510 2555.870 ;
        RECT 207.730 2553.090 208.910 2554.270 ;
        RECT 209.330 2553.090 210.510 2554.270 ;
        RECT 207.730 2374.690 208.910 2375.870 ;
        RECT 209.330 2374.690 210.510 2375.870 ;
        RECT 207.730 2373.090 208.910 2374.270 ;
        RECT 209.330 2373.090 210.510 2374.270 ;
        RECT 207.730 2194.690 208.910 2195.870 ;
        RECT 209.330 2194.690 210.510 2195.870 ;
        RECT 207.730 2193.090 208.910 2194.270 ;
        RECT 209.330 2193.090 210.510 2194.270 ;
        RECT 207.730 2014.690 208.910 2015.870 ;
        RECT 209.330 2014.690 210.510 2015.870 ;
        RECT 207.730 2013.090 208.910 2014.270 ;
        RECT 209.330 2013.090 210.510 2014.270 ;
        RECT 207.730 1834.690 208.910 1835.870 ;
        RECT 209.330 1834.690 210.510 1835.870 ;
        RECT 207.730 1833.090 208.910 1834.270 ;
        RECT 209.330 1833.090 210.510 1834.270 ;
        RECT 207.730 1654.690 208.910 1655.870 ;
        RECT 209.330 1654.690 210.510 1655.870 ;
        RECT 207.730 1653.090 208.910 1654.270 ;
        RECT 209.330 1653.090 210.510 1654.270 ;
        RECT 207.730 1474.690 208.910 1475.870 ;
        RECT 209.330 1474.690 210.510 1475.870 ;
        RECT 207.730 1473.090 208.910 1474.270 ;
        RECT 209.330 1473.090 210.510 1474.270 ;
        RECT 207.730 1294.690 208.910 1295.870 ;
        RECT 209.330 1294.690 210.510 1295.870 ;
        RECT 207.730 1293.090 208.910 1294.270 ;
        RECT 209.330 1293.090 210.510 1294.270 ;
        RECT 207.730 1114.690 208.910 1115.870 ;
        RECT 209.330 1114.690 210.510 1115.870 ;
        RECT 207.730 1113.090 208.910 1114.270 ;
        RECT 209.330 1113.090 210.510 1114.270 ;
        RECT 387.730 3532.610 388.910 3533.790 ;
        RECT 389.330 3532.610 390.510 3533.790 ;
        RECT 387.730 3531.010 388.910 3532.190 ;
        RECT 389.330 3531.010 390.510 3532.190 ;
        RECT 387.730 3454.690 388.910 3455.870 ;
        RECT 389.330 3454.690 390.510 3455.870 ;
        RECT 387.730 3453.090 388.910 3454.270 ;
        RECT 389.330 3453.090 390.510 3454.270 ;
        RECT 387.730 3274.690 388.910 3275.870 ;
        RECT 389.330 3274.690 390.510 3275.870 ;
        RECT 387.730 3273.090 388.910 3274.270 ;
        RECT 389.330 3273.090 390.510 3274.270 ;
        RECT 387.730 3094.690 388.910 3095.870 ;
        RECT 389.330 3094.690 390.510 3095.870 ;
        RECT 387.730 3093.090 388.910 3094.270 ;
        RECT 389.330 3093.090 390.510 3094.270 ;
        RECT 387.730 2914.690 388.910 2915.870 ;
        RECT 389.330 2914.690 390.510 2915.870 ;
        RECT 387.730 2913.090 388.910 2914.270 ;
        RECT 389.330 2913.090 390.510 2914.270 ;
        RECT 387.730 2734.690 388.910 2735.870 ;
        RECT 389.330 2734.690 390.510 2735.870 ;
        RECT 387.730 2733.090 388.910 2734.270 ;
        RECT 389.330 2733.090 390.510 2734.270 ;
        RECT 387.730 2554.690 388.910 2555.870 ;
        RECT 389.330 2554.690 390.510 2555.870 ;
        RECT 387.730 2553.090 388.910 2554.270 ;
        RECT 389.330 2553.090 390.510 2554.270 ;
        RECT 387.730 2374.690 388.910 2375.870 ;
        RECT 389.330 2374.690 390.510 2375.870 ;
        RECT 387.730 2373.090 388.910 2374.270 ;
        RECT 389.330 2373.090 390.510 2374.270 ;
        RECT 387.730 2194.690 388.910 2195.870 ;
        RECT 389.330 2194.690 390.510 2195.870 ;
        RECT 387.730 2193.090 388.910 2194.270 ;
        RECT 389.330 2193.090 390.510 2194.270 ;
        RECT 387.730 2014.690 388.910 2015.870 ;
        RECT 389.330 2014.690 390.510 2015.870 ;
        RECT 387.730 2013.090 388.910 2014.270 ;
        RECT 389.330 2013.090 390.510 2014.270 ;
        RECT 387.730 1834.690 388.910 1835.870 ;
        RECT 389.330 1834.690 390.510 1835.870 ;
        RECT 387.730 1833.090 388.910 1834.270 ;
        RECT 389.330 1833.090 390.510 1834.270 ;
        RECT 387.730 1654.690 388.910 1655.870 ;
        RECT 389.330 1654.690 390.510 1655.870 ;
        RECT 387.730 1653.090 388.910 1654.270 ;
        RECT 389.330 1653.090 390.510 1654.270 ;
        RECT 387.730 1474.690 388.910 1475.870 ;
        RECT 389.330 1474.690 390.510 1475.870 ;
        RECT 387.730 1473.090 388.910 1474.270 ;
        RECT 389.330 1473.090 390.510 1474.270 ;
        RECT 387.730 1294.690 388.910 1295.870 ;
        RECT 389.330 1294.690 390.510 1295.870 ;
        RECT 387.730 1293.090 388.910 1294.270 ;
        RECT 389.330 1293.090 390.510 1294.270 ;
        RECT 387.730 1114.690 388.910 1115.870 ;
        RECT 389.330 1114.690 390.510 1115.870 ;
        RECT 387.730 1113.090 388.910 1114.270 ;
        RECT 389.330 1113.090 390.510 1114.270 ;
        RECT 567.730 3532.610 568.910 3533.790 ;
        RECT 569.330 3532.610 570.510 3533.790 ;
        RECT 567.730 3531.010 568.910 3532.190 ;
        RECT 569.330 3531.010 570.510 3532.190 ;
        RECT 567.730 3454.690 568.910 3455.870 ;
        RECT 569.330 3454.690 570.510 3455.870 ;
        RECT 567.730 3453.090 568.910 3454.270 ;
        RECT 569.330 3453.090 570.510 3454.270 ;
        RECT 567.730 3274.690 568.910 3275.870 ;
        RECT 569.330 3274.690 570.510 3275.870 ;
        RECT 567.730 3273.090 568.910 3274.270 ;
        RECT 569.330 3273.090 570.510 3274.270 ;
        RECT 567.730 3094.690 568.910 3095.870 ;
        RECT 569.330 3094.690 570.510 3095.870 ;
        RECT 567.730 3093.090 568.910 3094.270 ;
        RECT 569.330 3093.090 570.510 3094.270 ;
        RECT 567.730 2914.690 568.910 2915.870 ;
        RECT 569.330 2914.690 570.510 2915.870 ;
        RECT 567.730 2913.090 568.910 2914.270 ;
        RECT 569.330 2913.090 570.510 2914.270 ;
        RECT 567.730 2734.690 568.910 2735.870 ;
        RECT 569.330 2734.690 570.510 2735.870 ;
        RECT 567.730 2733.090 568.910 2734.270 ;
        RECT 569.330 2733.090 570.510 2734.270 ;
        RECT 567.730 2554.690 568.910 2555.870 ;
        RECT 569.330 2554.690 570.510 2555.870 ;
        RECT 567.730 2553.090 568.910 2554.270 ;
        RECT 569.330 2553.090 570.510 2554.270 ;
        RECT 567.730 2374.690 568.910 2375.870 ;
        RECT 569.330 2374.690 570.510 2375.870 ;
        RECT 567.730 2373.090 568.910 2374.270 ;
        RECT 569.330 2373.090 570.510 2374.270 ;
        RECT 567.730 2194.690 568.910 2195.870 ;
        RECT 569.330 2194.690 570.510 2195.870 ;
        RECT 567.730 2193.090 568.910 2194.270 ;
        RECT 569.330 2193.090 570.510 2194.270 ;
        RECT 567.730 2014.690 568.910 2015.870 ;
        RECT 569.330 2014.690 570.510 2015.870 ;
        RECT 567.730 2013.090 568.910 2014.270 ;
        RECT 569.330 2013.090 570.510 2014.270 ;
        RECT 567.730 1834.690 568.910 1835.870 ;
        RECT 569.330 1834.690 570.510 1835.870 ;
        RECT 567.730 1833.090 568.910 1834.270 ;
        RECT 569.330 1833.090 570.510 1834.270 ;
        RECT 567.730 1654.690 568.910 1655.870 ;
        RECT 569.330 1654.690 570.510 1655.870 ;
        RECT 567.730 1653.090 568.910 1654.270 ;
        RECT 569.330 1653.090 570.510 1654.270 ;
        RECT 567.730 1474.690 568.910 1475.870 ;
        RECT 569.330 1474.690 570.510 1475.870 ;
        RECT 567.730 1473.090 568.910 1474.270 ;
        RECT 569.330 1473.090 570.510 1474.270 ;
        RECT 567.730 1294.690 568.910 1295.870 ;
        RECT 569.330 1294.690 570.510 1295.870 ;
        RECT 567.730 1293.090 568.910 1294.270 ;
        RECT 569.330 1293.090 570.510 1294.270 ;
        RECT 567.730 1114.690 568.910 1115.870 ;
        RECT 569.330 1114.690 570.510 1115.870 ;
        RECT 567.730 1113.090 568.910 1114.270 ;
        RECT 569.330 1113.090 570.510 1114.270 ;
        RECT 747.730 3532.610 748.910 3533.790 ;
        RECT 749.330 3532.610 750.510 3533.790 ;
        RECT 747.730 3531.010 748.910 3532.190 ;
        RECT 749.330 3531.010 750.510 3532.190 ;
        RECT 747.730 3454.690 748.910 3455.870 ;
        RECT 749.330 3454.690 750.510 3455.870 ;
        RECT 747.730 3453.090 748.910 3454.270 ;
        RECT 749.330 3453.090 750.510 3454.270 ;
        RECT 747.730 3274.690 748.910 3275.870 ;
        RECT 749.330 3274.690 750.510 3275.870 ;
        RECT 747.730 3273.090 748.910 3274.270 ;
        RECT 749.330 3273.090 750.510 3274.270 ;
        RECT 747.730 3094.690 748.910 3095.870 ;
        RECT 749.330 3094.690 750.510 3095.870 ;
        RECT 747.730 3093.090 748.910 3094.270 ;
        RECT 749.330 3093.090 750.510 3094.270 ;
        RECT 747.730 2914.690 748.910 2915.870 ;
        RECT 749.330 2914.690 750.510 2915.870 ;
        RECT 747.730 2913.090 748.910 2914.270 ;
        RECT 749.330 2913.090 750.510 2914.270 ;
        RECT 747.730 2734.690 748.910 2735.870 ;
        RECT 749.330 2734.690 750.510 2735.870 ;
        RECT 747.730 2733.090 748.910 2734.270 ;
        RECT 749.330 2733.090 750.510 2734.270 ;
        RECT 747.730 2554.690 748.910 2555.870 ;
        RECT 749.330 2554.690 750.510 2555.870 ;
        RECT 747.730 2553.090 748.910 2554.270 ;
        RECT 749.330 2553.090 750.510 2554.270 ;
        RECT 747.730 2374.690 748.910 2375.870 ;
        RECT 749.330 2374.690 750.510 2375.870 ;
        RECT 747.730 2373.090 748.910 2374.270 ;
        RECT 749.330 2373.090 750.510 2374.270 ;
        RECT 747.730 2194.690 748.910 2195.870 ;
        RECT 749.330 2194.690 750.510 2195.870 ;
        RECT 747.730 2193.090 748.910 2194.270 ;
        RECT 749.330 2193.090 750.510 2194.270 ;
        RECT 747.730 2014.690 748.910 2015.870 ;
        RECT 749.330 2014.690 750.510 2015.870 ;
        RECT 747.730 2013.090 748.910 2014.270 ;
        RECT 749.330 2013.090 750.510 2014.270 ;
        RECT 747.730 1834.690 748.910 1835.870 ;
        RECT 749.330 1834.690 750.510 1835.870 ;
        RECT 747.730 1833.090 748.910 1834.270 ;
        RECT 749.330 1833.090 750.510 1834.270 ;
        RECT 747.730 1654.690 748.910 1655.870 ;
        RECT 749.330 1654.690 750.510 1655.870 ;
        RECT 747.730 1653.090 748.910 1654.270 ;
        RECT 749.330 1653.090 750.510 1654.270 ;
        RECT 747.730 1474.690 748.910 1475.870 ;
        RECT 749.330 1474.690 750.510 1475.870 ;
        RECT 747.730 1473.090 748.910 1474.270 ;
        RECT 749.330 1473.090 750.510 1474.270 ;
        RECT 747.730 1294.690 748.910 1295.870 ;
        RECT 749.330 1294.690 750.510 1295.870 ;
        RECT 747.730 1293.090 748.910 1294.270 ;
        RECT 749.330 1293.090 750.510 1294.270 ;
        RECT 747.730 1114.690 748.910 1115.870 ;
        RECT 749.330 1114.690 750.510 1115.870 ;
        RECT 747.730 1113.090 748.910 1114.270 ;
        RECT 749.330 1113.090 750.510 1114.270 ;
        RECT 927.730 3532.610 928.910 3533.790 ;
        RECT 929.330 3532.610 930.510 3533.790 ;
        RECT 927.730 3531.010 928.910 3532.190 ;
        RECT 929.330 3531.010 930.510 3532.190 ;
        RECT 927.730 3454.690 928.910 3455.870 ;
        RECT 929.330 3454.690 930.510 3455.870 ;
        RECT 927.730 3453.090 928.910 3454.270 ;
        RECT 929.330 3453.090 930.510 3454.270 ;
        RECT 927.730 3274.690 928.910 3275.870 ;
        RECT 929.330 3274.690 930.510 3275.870 ;
        RECT 927.730 3273.090 928.910 3274.270 ;
        RECT 929.330 3273.090 930.510 3274.270 ;
        RECT 927.730 3094.690 928.910 3095.870 ;
        RECT 929.330 3094.690 930.510 3095.870 ;
        RECT 927.730 3093.090 928.910 3094.270 ;
        RECT 929.330 3093.090 930.510 3094.270 ;
        RECT 927.730 2914.690 928.910 2915.870 ;
        RECT 929.330 2914.690 930.510 2915.870 ;
        RECT 927.730 2913.090 928.910 2914.270 ;
        RECT 929.330 2913.090 930.510 2914.270 ;
        RECT 927.730 2734.690 928.910 2735.870 ;
        RECT 929.330 2734.690 930.510 2735.870 ;
        RECT 927.730 2733.090 928.910 2734.270 ;
        RECT 929.330 2733.090 930.510 2734.270 ;
        RECT 927.730 2554.690 928.910 2555.870 ;
        RECT 929.330 2554.690 930.510 2555.870 ;
        RECT 927.730 2553.090 928.910 2554.270 ;
        RECT 929.330 2553.090 930.510 2554.270 ;
        RECT 927.730 2374.690 928.910 2375.870 ;
        RECT 929.330 2374.690 930.510 2375.870 ;
        RECT 927.730 2373.090 928.910 2374.270 ;
        RECT 929.330 2373.090 930.510 2374.270 ;
        RECT 927.730 2194.690 928.910 2195.870 ;
        RECT 929.330 2194.690 930.510 2195.870 ;
        RECT 927.730 2193.090 928.910 2194.270 ;
        RECT 929.330 2193.090 930.510 2194.270 ;
        RECT 927.730 2014.690 928.910 2015.870 ;
        RECT 929.330 2014.690 930.510 2015.870 ;
        RECT 927.730 2013.090 928.910 2014.270 ;
        RECT 929.330 2013.090 930.510 2014.270 ;
        RECT 927.730 1834.690 928.910 1835.870 ;
        RECT 929.330 1834.690 930.510 1835.870 ;
        RECT 927.730 1833.090 928.910 1834.270 ;
        RECT 929.330 1833.090 930.510 1834.270 ;
        RECT 927.730 1654.690 928.910 1655.870 ;
        RECT 929.330 1654.690 930.510 1655.870 ;
        RECT 927.730 1653.090 928.910 1654.270 ;
        RECT 929.330 1653.090 930.510 1654.270 ;
        RECT 927.730 1474.690 928.910 1475.870 ;
        RECT 929.330 1474.690 930.510 1475.870 ;
        RECT 927.730 1473.090 928.910 1474.270 ;
        RECT 929.330 1473.090 930.510 1474.270 ;
        RECT 927.730 1294.690 928.910 1295.870 ;
        RECT 929.330 1294.690 930.510 1295.870 ;
        RECT 927.730 1293.090 928.910 1294.270 ;
        RECT 929.330 1293.090 930.510 1294.270 ;
        RECT 927.730 1114.690 928.910 1115.870 ;
        RECT 929.330 1114.690 930.510 1115.870 ;
        RECT 927.730 1113.090 928.910 1114.270 ;
        RECT 929.330 1113.090 930.510 1114.270 ;
        RECT 1107.730 3532.610 1108.910 3533.790 ;
        RECT 1109.330 3532.610 1110.510 3533.790 ;
        RECT 1107.730 3531.010 1108.910 3532.190 ;
        RECT 1109.330 3531.010 1110.510 3532.190 ;
        RECT 1107.730 3454.690 1108.910 3455.870 ;
        RECT 1109.330 3454.690 1110.510 3455.870 ;
        RECT 1107.730 3453.090 1108.910 3454.270 ;
        RECT 1109.330 3453.090 1110.510 3454.270 ;
        RECT 1107.730 3274.690 1108.910 3275.870 ;
        RECT 1109.330 3274.690 1110.510 3275.870 ;
        RECT 1107.730 3273.090 1108.910 3274.270 ;
        RECT 1109.330 3273.090 1110.510 3274.270 ;
        RECT 1107.730 3094.690 1108.910 3095.870 ;
        RECT 1109.330 3094.690 1110.510 3095.870 ;
        RECT 1107.730 3093.090 1108.910 3094.270 ;
        RECT 1109.330 3093.090 1110.510 3094.270 ;
        RECT 1107.730 2914.690 1108.910 2915.870 ;
        RECT 1109.330 2914.690 1110.510 2915.870 ;
        RECT 1107.730 2913.090 1108.910 2914.270 ;
        RECT 1109.330 2913.090 1110.510 2914.270 ;
        RECT 1107.730 2734.690 1108.910 2735.870 ;
        RECT 1109.330 2734.690 1110.510 2735.870 ;
        RECT 1107.730 2733.090 1108.910 2734.270 ;
        RECT 1109.330 2733.090 1110.510 2734.270 ;
        RECT 1107.730 2554.690 1108.910 2555.870 ;
        RECT 1109.330 2554.690 1110.510 2555.870 ;
        RECT 1107.730 2553.090 1108.910 2554.270 ;
        RECT 1109.330 2553.090 1110.510 2554.270 ;
        RECT 1107.730 2374.690 1108.910 2375.870 ;
        RECT 1109.330 2374.690 1110.510 2375.870 ;
        RECT 1107.730 2373.090 1108.910 2374.270 ;
        RECT 1109.330 2373.090 1110.510 2374.270 ;
        RECT 1107.730 2194.690 1108.910 2195.870 ;
        RECT 1109.330 2194.690 1110.510 2195.870 ;
        RECT 1107.730 2193.090 1108.910 2194.270 ;
        RECT 1109.330 2193.090 1110.510 2194.270 ;
        RECT 1107.730 2014.690 1108.910 2015.870 ;
        RECT 1109.330 2014.690 1110.510 2015.870 ;
        RECT 1107.730 2013.090 1108.910 2014.270 ;
        RECT 1109.330 2013.090 1110.510 2014.270 ;
        RECT 1107.730 1834.690 1108.910 1835.870 ;
        RECT 1109.330 1834.690 1110.510 1835.870 ;
        RECT 1107.730 1833.090 1108.910 1834.270 ;
        RECT 1109.330 1833.090 1110.510 1834.270 ;
        RECT 1107.730 1654.690 1108.910 1655.870 ;
        RECT 1109.330 1654.690 1110.510 1655.870 ;
        RECT 1107.730 1653.090 1108.910 1654.270 ;
        RECT 1109.330 1653.090 1110.510 1654.270 ;
        RECT 1107.730 1474.690 1108.910 1475.870 ;
        RECT 1109.330 1474.690 1110.510 1475.870 ;
        RECT 1107.730 1473.090 1108.910 1474.270 ;
        RECT 1109.330 1473.090 1110.510 1474.270 ;
        RECT 1107.730 1294.690 1108.910 1295.870 ;
        RECT 1109.330 1294.690 1110.510 1295.870 ;
        RECT 1107.730 1293.090 1108.910 1294.270 ;
        RECT 1109.330 1293.090 1110.510 1294.270 ;
        RECT 1107.730 1114.690 1108.910 1115.870 ;
        RECT 1109.330 1114.690 1110.510 1115.870 ;
        RECT 1107.730 1113.090 1108.910 1114.270 ;
        RECT 1109.330 1113.090 1110.510 1114.270 ;
        RECT 1287.730 3532.610 1288.910 3533.790 ;
        RECT 1289.330 3532.610 1290.510 3533.790 ;
        RECT 1287.730 3531.010 1288.910 3532.190 ;
        RECT 1289.330 3531.010 1290.510 3532.190 ;
        RECT 1287.730 3454.690 1288.910 3455.870 ;
        RECT 1289.330 3454.690 1290.510 3455.870 ;
        RECT 1287.730 3453.090 1288.910 3454.270 ;
        RECT 1289.330 3453.090 1290.510 3454.270 ;
        RECT 1287.730 3274.690 1288.910 3275.870 ;
        RECT 1289.330 3274.690 1290.510 3275.870 ;
        RECT 1287.730 3273.090 1288.910 3274.270 ;
        RECT 1289.330 3273.090 1290.510 3274.270 ;
        RECT 1287.730 3094.690 1288.910 3095.870 ;
        RECT 1289.330 3094.690 1290.510 3095.870 ;
        RECT 1287.730 3093.090 1288.910 3094.270 ;
        RECT 1289.330 3093.090 1290.510 3094.270 ;
        RECT 1287.730 2914.690 1288.910 2915.870 ;
        RECT 1289.330 2914.690 1290.510 2915.870 ;
        RECT 1287.730 2913.090 1288.910 2914.270 ;
        RECT 1289.330 2913.090 1290.510 2914.270 ;
        RECT 1287.730 2734.690 1288.910 2735.870 ;
        RECT 1289.330 2734.690 1290.510 2735.870 ;
        RECT 1287.730 2733.090 1288.910 2734.270 ;
        RECT 1289.330 2733.090 1290.510 2734.270 ;
        RECT 1287.730 2554.690 1288.910 2555.870 ;
        RECT 1289.330 2554.690 1290.510 2555.870 ;
        RECT 1287.730 2553.090 1288.910 2554.270 ;
        RECT 1289.330 2553.090 1290.510 2554.270 ;
        RECT 1287.730 2374.690 1288.910 2375.870 ;
        RECT 1289.330 2374.690 1290.510 2375.870 ;
        RECT 1287.730 2373.090 1288.910 2374.270 ;
        RECT 1289.330 2373.090 1290.510 2374.270 ;
        RECT 1287.730 2194.690 1288.910 2195.870 ;
        RECT 1289.330 2194.690 1290.510 2195.870 ;
        RECT 1287.730 2193.090 1288.910 2194.270 ;
        RECT 1289.330 2193.090 1290.510 2194.270 ;
        RECT 1287.730 2014.690 1288.910 2015.870 ;
        RECT 1289.330 2014.690 1290.510 2015.870 ;
        RECT 1287.730 2013.090 1288.910 2014.270 ;
        RECT 1289.330 2013.090 1290.510 2014.270 ;
        RECT 1287.730 1834.690 1288.910 1835.870 ;
        RECT 1289.330 1834.690 1290.510 1835.870 ;
        RECT 1287.730 1833.090 1288.910 1834.270 ;
        RECT 1289.330 1833.090 1290.510 1834.270 ;
        RECT 1287.730 1654.690 1288.910 1655.870 ;
        RECT 1289.330 1654.690 1290.510 1655.870 ;
        RECT 1287.730 1653.090 1288.910 1654.270 ;
        RECT 1289.330 1653.090 1290.510 1654.270 ;
        RECT 1287.730 1474.690 1288.910 1475.870 ;
        RECT 1289.330 1474.690 1290.510 1475.870 ;
        RECT 1287.730 1473.090 1288.910 1474.270 ;
        RECT 1289.330 1473.090 1290.510 1474.270 ;
        RECT 1287.730 1294.690 1288.910 1295.870 ;
        RECT 1289.330 1294.690 1290.510 1295.870 ;
        RECT 1287.730 1293.090 1288.910 1294.270 ;
        RECT 1289.330 1293.090 1290.510 1294.270 ;
        RECT 1287.730 1114.690 1288.910 1115.870 ;
        RECT 1289.330 1114.690 1290.510 1115.870 ;
        RECT 1287.730 1113.090 1288.910 1114.270 ;
        RECT 1289.330 1113.090 1290.510 1114.270 ;
        RECT 27.730 934.690 28.910 935.870 ;
        RECT 29.330 934.690 30.510 935.870 ;
        RECT 27.730 933.090 28.910 934.270 ;
        RECT 29.330 933.090 30.510 934.270 ;
        RECT 27.730 754.690 28.910 755.870 ;
        RECT 29.330 754.690 30.510 755.870 ;
        RECT 27.730 753.090 28.910 754.270 ;
        RECT 29.330 753.090 30.510 754.270 ;
        RECT 27.730 574.690 28.910 575.870 ;
        RECT 29.330 574.690 30.510 575.870 ;
        RECT 27.730 573.090 28.910 574.270 ;
        RECT 29.330 573.090 30.510 574.270 ;
        RECT 27.730 394.690 28.910 395.870 ;
        RECT 29.330 394.690 30.510 395.870 ;
        RECT 27.730 393.090 28.910 394.270 ;
        RECT 29.330 393.090 30.510 394.270 ;
        RECT 1287.730 934.690 1288.910 935.870 ;
        RECT 1289.330 934.690 1290.510 935.870 ;
        RECT 1287.730 933.090 1288.910 934.270 ;
        RECT 1289.330 933.090 1290.510 934.270 ;
        RECT 1287.730 754.690 1288.910 755.870 ;
        RECT 1289.330 754.690 1290.510 755.870 ;
        RECT 1287.730 753.090 1288.910 754.270 ;
        RECT 1289.330 753.090 1290.510 754.270 ;
        RECT 1287.730 574.690 1288.910 575.870 ;
        RECT 1289.330 574.690 1290.510 575.870 ;
        RECT 1287.730 573.090 1288.910 574.270 ;
        RECT 1289.330 573.090 1290.510 574.270 ;
        RECT 1287.730 394.690 1288.910 395.870 ;
        RECT 1289.330 394.690 1290.510 395.870 ;
        RECT 1287.730 393.090 1288.910 394.270 ;
        RECT 1289.330 393.090 1290.510 394.270 ;
        RECT 27.730 214.690 28.910 215.870 ;
        RECT 29.330 214.690 30.510 215.870 ;
        RECT 27.730 213.090 28.910 214.270 ;
        RECT 29.330 213.090 30.510 214.270 ;
        RECT 27.730 34.690 28.910 35.870 ;
        RECT 29.330 34.690 30.510 35.870 ;
        RECT 27.730 33.090 28.910 34.270 ;
        RECT 29.330 33.090 30.510 34.270 ;
        RECT 27.730 -12.510 28.910 -11.330 ;
        RECT 29.330 -12.510 30.510 -11.330 ;
        RECT 27.730 -14.110 28.910 -12.930 ;
        RECT 29.330 -14.110 30.510 -12.930 ;
        RECT 207.730 214.690 208.910 215.870 ;
        RECT 209.330 214.690 210.510 215.870 ;
        RECT 207.730 213.090 208.910 214.270 ;
        RECT 209.330 213.090 210.510 214.270 ;
        RECT 207.730 34.690 208.910 35.870 ;
        RECT 209.330 34.690 210.510 35.870 ;
        RECT 207.730 33.090 208.910 34.270 ;
        RECT 209.330 33.090 210.510 34.270 ;
        RECT 207.730 -12.510 208.910 -11.330 ;
        RECT 209.330 -12.510 210.510 -11.330 ;
        RECT 207.730 -14.110 208.910 -12.930 ;
        RECT 209.330 -14.110 210.510 -12.930 ;
        RECT 387.730 214.690 388.910 215.870 ;
        RECT 389.330 214.690 390.510 215.870 ;
        RECT 387.730 213.090 388.910 214.270 ;
        RECT 389.330 213.090 390.510 214.270 ;
        RECT 387.730 34.690 388.910 35.870 ;
        RECT 389.330 34.690 390.510 35.870 ;
        RECT 387.730 33.090 388.910 34.270 ;
        RECT 389.330 33.090 390.510 34.270 ;
        RECT 387.730 -12.510 388.910 -11.330 ;
        RECT 389.330 -12.510 390.510 -11.330 ;
        RECT 387.730 -14.110 388.910 -12.930 ;
        RECT 389.330 -14.110 390.510 -12.930 ;
        RECT 567.730 214.690 568.910 215.870 ;
        RECT 569.330 214.690 570.510 215.870 ;
        RECT 567.730 213.090 568.910 214.270 ;
        RECT 569.330 213.090 570.510 214.270 ;
        RECT 567.730 34.690 568.910 35.870 ;
        RECT 569.330 34.690 570.510 35.870 ;
        RECT 567.730 33.090 568.910 34.270 ;
        RECT 569.330 33.090 570.510 34.270 ;
        RECT 567.730 -12.510 568.910 -11.330 ;
        RECT 569.330 -12.510 570.510 -11.330 ;
        RECT 567.730 -14.110 568.910 -12.930 ;
        RECT 569.330 -14.110 570.510 -12.930 ;
        RECT 747.730 214.690 748.910 215.870 ;
        RECT 749.330 214.690 750.510 215.870 ;
        RECT 747.730 213.090 748.910 214.270 ;
        RECT 749.330 213.090 750.510 214.270 ;
        RECT 747.730 34.690 748.910 35.870 ;
        RECT 749.330 34.690 750.510 35.870 ;
        RECT 747.730 33.090 748.910 34.270 ;
        RECT 749.330 33.090 750.510 34.270 ;
        RECT 747.730 -12.510 748.910 -11.330 ;
        RECT 749.330 -12.510 750.510 -11.330 ;
        RECT 747.730 -14.110 748.910 -12.930 ;
        RECT 749.330 -14.110 750.510 -12.930 ;
        RECT 927.730 214.690 928.910 215.870 ;
        RECT 929.330 214.690 930.510 215.870 ;
        RECT 927.730 213.090 928.910 214.270 ;
        RECT 929.330 213.090 930.510 214.270 ;
        RECT 927.730 34.690 928.910 35.870 ;
        RECT 929.330 34.690 930.510 35.870 ;
        RECT 927.730 33.090 928.910 34.270 ;
        RECT 929.330 33.090 930.510 34.270 ;
        RECT 927.730 -12.510 928.910 -11.330 ;
        RECT 929.330 -12.510 930.510 -11.330 ;
        RECT 927.730 -14.110 928.910 -12.930 ;
        RECT 929.330 -14.110 930.510 -12.930 ;
        RECT 1107.730 214.690 1108.910 215.870 ;
        RECT 1109.330 214.690 1110.510 215.870 ;
        RECT 1107.730 213.090 1108.910 214.270 ;
        RECT 1109.330 213.090 1110.510 214.270 ;
        RECT 1107.730 34.690 1108.910 35.870 ;
        RECT 1109.330 34.690 1110.510 35.870 ;
        RECT 1107.730 33.090 1108.910 34.270 ;
        RECT 1109.330 33.090 1110.510 34.270 ;
        RECT 1107.730 -12.510 1108.910 -11.330 ;
        RECT 1109.330 -12.510 1110.510 -11.330 ;
        RECT 1107.730 -14.110 1108.910 -12.930 ;
        RECT 1109.330 -14.110 1110.510 -12.930 ;
        RECT 1287.730 214.690 1288.910 215.870 ;
        RECT 1289.330 214.690 1290.510 215.870 ;
        RECT 1287.730 213.090 1288.910 214.270 ;
        RECT 1289.330 213.090 1290.510 214.270 ;
        RECT 1287.730 34.690 1288.910 35.870 ;
        RECT 1289.330 34.690 1290.510 35.870 ;
        RECT 1287.730 33.090 1288.910 34.270 ;
        RECT 1289.330 33.090 1290.510 34.270 ;
        RECT 1287.730 -12.510 1288.910 -11.330 ;
        RECT 1289.330 -12.510 1290.510 -11.330 ;
        RECT 1287.730 -14.110 1288.910 -12.930 ;
        RECT 1289.330 -14.110 1290.510 -12.930 ;
        RECT 1467.730 3532.610 1468.910 3533.790 ;
        RECT 1469.330 3532.610 1470.510 3533.790 ;
        RECT 1467.730 3531.010 1468.910 3532.190 ;
        RECT 1469.330 3531.010 1470.510 3532.190 ;
        RECT 1467.730 3454.690 1468.910 3455.870 ;
        RECT 1469.330 3454.690 1470.510 3455.870 ;
        RECT 1467.730 3453.090 1468.910 3454.270 ;
        RECT 1469.330 3453.090 1470.510 3454.270 ;
        RECT 1467.730 3274.690 1468.910 3275.870 ;
        RECT 1469.330 3274.690 1470.510 3275.870 ;
        RECT 1467.730 3273.090 1468.910 3274.270 ;
        RECT 1469.330 3273.090 1470.510 3274.270 ;
        RECT 1467.730 3094.690 1468.910 3095.870 ;
        RECT 1469.330 3094.690 1470.510 3095.870 ;
        RECT 1467.730 3093.090 1468.910 3094.270 ;
        RECT 1469.330 3093.090 1470.510 3094.270 ;
        RECT 1467.730 2914.690 1468.910 2915.870 ;
        RECT 1469.330 2914.690 1470.510 2915.870 ;
        RECT 1467.730 2913.090 1468.910 2914.270 ;
        RECT 1469.330 2913.090 1470.510 2914.270 ;
        RECT 1467.730 2734.690 1468.910 2735.870 ;
        RECT 1469.330 2734.690 1470.510 2735.870 ;
        RECT 1467.730 2733.090 1468.910 2734.270 ;
        RECT 1469.330 2733.090 1470.510 2734.270 ;
        RECT 1467.730 2554.690 1468.910 2555.870 ;
        RECT 1469.330 2554.690 1470.510 2555.870 ;
        RECT 1467.730 2553.090 1468.910 2554.270 ;
        RECT 1469.330 2553.090 1470.510 2554.270 ;
        RECT 1467.730 2374.690 1468.910 2375.870 ;
        RECT 1469.330 2374.690 1470.510 2375.870 ;
        RECT 1467.730 2373.090 1468.910 2374.270 ;
        RECT 1469.330 2373.090 1470.510 2374.270 ;
        RECT 1467.730 2194.690 1468.910 2195.870 ;
        RECT 1469.330 2194.690 1470.510 2195.870 ;
        RECT 1467.730 2193.090 1468.910 2194.270 ;
        RECT 1469.330 2193.090 1470.510 2194.270 ;
        RECT 1467.730 2014.690 1468.910 2015.870 ;
        RECT 1469.330 2014.690 1470.510 2015.870 ;
        RECT 1467.730 2013.090 1468.910 2014.270 ;
        RECT 1469.330 2013.090 1470.510 2014.270 ;
        RECT 1467.730 1834.690 1468.910 1835.870 ;
        RECT 1469.330 1834.690 1470.510 1835.870 ;
        RECT 1467.730 1833.090 1468.910 1834.270 ;
        RECT 1469.330 1833.090 1470.510 1834.270 ;
        RECT 1467.730 1654.690 1468.910 1655.870 ;
        RECT 1469.330 1654.690 1470.510 1655.870 ;
        RECT 1467.730 1653.090 1468.910 1654.270 ;
        RECT 1469.330 1653.090 1470.510 1654.270 ;
        RECT 1467.730 1474.690 1468.910 1475.870 ;
        RECT 1469.330 1474.690 1470.510 1475.870 ;
        RECT 1467.730 1473.090 1468.910 1474.270 ;
        RECT 1469.330 1473.090 1470.510 1474.270 ;
        RECT 1467.730 1294.690 1468.910 1295.870 ;
        RECT 1469.330 1294.690 1470.510 1295.870 ;
        RECT 1467.730 1293.090 1468.910 1294.270 ;
        RECT 1469.330 1293.090 1470.510 1294.270 ;
        RECT 1467.730 1114.690 1468.910 1115.870 ;
        RECT 1469.330 1114.690 1470.510 1115.870 ;
        RECT 1467.730 1113.090 1468.910 1114.270 ;
        RECT 1469.330 1113.090 1470.510 1114.270 ;
        RECT 1467.730 934.690 1468.910 935.870 ;
        RECT 1469.330 934.690 1470.510 935.870 ;
        RECT 1467.730 933.090 1468.910 934.270 ;
        RECT 1469.330 933.090 1470.510 934.270 ;
        RECT 1467.730 754.690 1468.910 755.870 ;
        RECT 1469.330 754.690 1470.510 755.870 ;
        RECT 1467.730 753.090 1468.910 754.270 ;
        RECT 1469.330 753.090 1470.510 754.270 ;
        RECT 1467.730 574.690 1468.910 575.870 ;
        RECT 1469.330 574.690 1470.510 575.870 ;
        RECT 1467.730 573.090 1468.910 574.270 ;
        RECT 1469.330 573.090 1470.510 574.270 ;
        RECT 1467.730 394.690 1468.910 395.870 ;
        RECT 1469.330 394.690 1470.510 395.870 ;
        RECT 1467.730 393.090 1468.910 394.270 ;
        RECT 1469.330 393.090 1470.510 394.270 ;
        RECT 1467.730 214.690 1468.910 215.870 ;
        RECT 1469.330 214.690 1470.510 215.870 ;
        RECT 1467.730 213.090 1468.910 214.270 ;
        RECT 1469.330 213.090 1470.510 214.270 ;
        RECT 1467.730 34.690 1468.910 35.870 ;
        RECT 1469.330 34.690 1470.510 35.870 ;
        RECT 1467.730 33.090 1468.910 34.270 ;
        RECT 1469.330 33.090 1470.510 34.270 ;
        RECT 1467.730 -12.510 1468.910 -11.330 ;
        RECT 1469.330 -12.510 1470.510 -11.330 ;
        RECT 1467.730 -14.110 1468.910 -12.930 ;
        RECT 1469.330 -14.110 1470.510 -12.930 ;
        RECT 1647.730 3532.610 1648.910 3533.790 ;
        RECT 1649.330 3532.610 1650.510 3533.790 ;
        RECT 1647.730 3531.010 1648.910 3532.190 ;
        RECT 1649.330 3531.010 1650.510 3532.190 ;
        RECT 1647.730 3454.690 1648.910 3455.870 ;
        RECT 1649.330 3454.690 1650.510 3455.870 ;
        RECT 1647.730 3453.090 1648.910 3454.270 ;
        RECT 1649.330 3453.090 1650.510 3454.270 ;
        RECT 1647.730 3274.690 1648.910 3275.870 ;
        RECT 1649.330 3274.690 1650.510 3275.870 ;
        RECT 1647.730 3273.090 1648.910 3274.270 ;
        RECT 1649.330 3273.090 1650.510 3274.270 ;
        RECT 1647.730 3094.690 1648.910 3095.870 ;
        RECT 1649.330 3094.690 1650.510 3095.870 ;
        RECT 1647.730 3093.090 1648.910 3094.270 ;
        RECT 1649.330 3093.090 1650.510 3094.270 ;
        RECT 1647.730 2914.690 1648.910 2915.870 ;
        RECT 1649.330 2914.690 1650.510 2915.870 ;
        RECT 1647.730 2913.090 1648.910 2914.270 ;
        RECT 1649.330 2913.090 1650.510 2914.270 ;
        RECT 1647.730 2734.690 1648.910 2735.870 ;
        RECT 1649.330 2734.690 1650.510 2735.870 ;
        RECT 1647.730 2733.090 1648.910 2734.270 ;
        RECT 1649.330 2733.090 1650.510 2734.270 ;
        RECT 1647.730 2554.690 1648.910 2555.870 ;
        RECT 1649.330 2554.690 1650.510 2555.870 ;
        RECT 1647.730 2553.090 1648.910 2554.270 ;
        RECT 1649.330 2553.090 1650.510 2554.270 ;
        RECT 1647.730 2374.690 1648.910 2375.870 ;
        RECT 1649.330 2374.690 1650.510 2375.870 ;
        RECT 1647.730 2373.090 1648.910 2374.270 ;
        RECT 1649.330 2373.090 1650.510 2374.270 ;
        RECT 1647.730 2194.690 1648.910 2195.870 ;
        RECT 1649.330 2194.690 1650.510 2195.870 ;
        RECT 1647.730 2193.090 1648.910 2194.270 ;
        RECT 1649.330 2193.090 1650.510 2194.270 ;
        RECT 1647.730 2014.690 1648.910 2015.870 ;
        RECT 1649.330 2014.690 1650.510 2015.870 ;
        RECT 1647.730 2013.090 1648.910 2014.270 ;
        RECT 1649.330 2013.090 1650.510 2014.270 ;
        RECT 1647.730 1834.690 1648.910 1835.870 ;
        RECT 1649.330 1834.690 1650.510 1835.870 ;
        RECT 1647.730 1833.090 1648.910 1834.270 ;
        RECT 1649.330 1833.090 1650.510 1834.270 ;
        RECT 1647.730 1654.690 1648.910 1655.870 ;
        RECT 1649.330 1654.690 1650.510 1655.870 ;
        RECT 1647.730 1653.090 1648.910 1654.270 ;
        RECT 1649.330 1653.090 1650.510 1654.270 ;
        RECT 1647.730 1474.690 1648.910 1475.870 ;
        RECT 1649.330 1474.690 1650.510 1475.870 ;
        RECT 1647.730 1473.090 1648.910 1474.270 ;
        RECT 1649.330 1473.090 1650.510 1474.270 ;
        RECT 1647.730 1294.690 1648.910 1295.870 ;
        RECT 1649.330 1294.690 1650.510 1295.870 ;
        RECT 1647.730 1293.090 1648.910 1294.270 ;
        RECT 1649.330 1293.090 1650.510 1294.270 ;
        RECT 1647.730 1114.690 1648.910 1115.870 ;
        RECT 1649.330 1114.690 1650.510 1115.870 ;
        RECT 1647.730 1113.090 1648.910 1114.270 ;
        RECT 1649.330 1113.090 1650.510 1114.270 ;
        RECT 1647.730 934.690 1648.910 935.870 ;
        RECT 1649.330 934.690 1650.510 935.870 ;
        RECT 1647.730 933.090 1648.910 934.270 ;
        RECT 1649.330 933.090 1650.510 934.270 ;
        RECT 1647.730 754.690 1648.910 755.870 ;
        RECT 1649.330 754.690 1650.510 755.870 ;
        RECT 1647.730 753.090 1648.910 754.270 ;
        RECT 1649.330 753.090 1650.510 754.270 ;
        RECT 1647.730 574.690 1648.910 575.870 ;
        RECT 1649.330 574.690 1650.510 575.870 ;
        RECT 1647.730 573.090 1648.910 574.270 ;
        RECT 1649.330 573.090 1650.510 574.270 ;
        RECT 1647.730 394.690 1648.910 395.870 ;
        RECT 1649.330 394.690 1650.510 395.870 ;
        RECT 1647.730 393.090 1648.910 394.270 ;
        RECT 1649.330 393.090 1650.510 394.270 ;
        RECT 1647.730 214.690 1648.910 215.870 ;
        RECT 1649.330 214.690 1650.510 215.870 ;
        RECT 1647.730 213.090 1648.910 214.270 ;
        RECT 1649.330 213.090 1650.510 214.270 ;
        RECT 1647.730 34.690 1648.910 35.870 ;
        RECT 1649.330 34.690 1650.510 35.870 ;
        RECT 1647.730 33.090 1648.910 34.270 ;
        RECT 1649.330 33.090 1650.510 34.270 ;
        RECT 1647.730 -12.510 1648.910 -11.330 ;
        RECT 1649.330 -12.510 1650.510 -11.330 ;
        RECT 1647.730 -14.110 1648.910 -12.930 ;
        RECT 1649.330 -14.110 1650.510 -12.930 ;
        RECT 1827.730 3532.610 1828.910 3533.790 ;
        RECT 1829.330 3532.610 1830.510 3533.790 ;
        RECT 1827.730 3531.010 1828.910 3532.190 ;
        RECT 1829.330 3531.010 1830.510 3532.190 ;
        RECT 1827.730 3454.690 1828.910 3455.870 ;
        RECT 1829.330 3454.690 1830.510 3455.870 ;
        RECT 1827.730 3453.090 1828.910 3454.270 ;
        RECT 1829.330 3453.090 1830.510 3454.270 ;
        RECT 1827.730 3274.690 1828.910 3275.870 ;
        RECT 1829.330 3274.690 1830.510 3275.870 ;
        RECT 1827.730 3273.090 1828.910 3274.270 ;
        RECT 1829.330 3273.090 1830.510 3274.270 ;
        RECT 1827.730 3094.690 1828.910 3095.870 ;
        RECT 1829.330 3094.690 1830.510 3095.870 ;
        RECT 1827.730 3093.090 1828.910 3094.270 ;
        RECT 1829.330 3093.090 1830.510 3094.270 ;
        RECT 1827.730 2914.690 1828.910 2915.870 ;
        RECT 1829.330 2914.690 1830.510 2915.870 ;
        RECT 1827.730 2913.090 1828.910 2914.270 ;
        RECT 1829.330 2913.090 1830.510 2914.270 ;
        RECT 1827.730 2734.690 1828.910 2735.870 ;
        RECT 1829.330 2734.690 1830.510 2735.870 ;
        RECT 1827.730 2733.090 1828.910 2734.270 ;
        RECT 1829.330 2733.090 1830.510 2734.270 ;
        RECT 1827.730 2554.690 1828.910 2555.870 ;
        RECT 1829.330 2554.690 1830.510 2555.870 ;
        RECT 1827.730 2553.090 1828.910 2554.270 ;
        RECT 1829.330 2553.090 1830.510 2554.270 ;
        RECT 1827.730 2374.690 1828.910 2375.870 ;
        RECT 1829.330 2374.690 1830.510 2375.870 ;
        RECT 1827.730 2373.090 1828.910 2374.270 ;
        RECT 1829.330 2373.090 1830.510 2374.270 ;
        RECT 1827.730 2194.690 1828.910 2195.870 ;
        RECT 1829.330 2194.690 1830.510 2195.870 ;
        RECT 1827.730 2193.090 1828.910 2194.270 ;
        RECT 1829.330 2193.090 1830.510 2194.270 ;
        RECT 1827.730 2014.690 1828.910 2015.870 ;
        RECT 1829.330 2014.690 1830.510 2015.870 ;
        RECT 1827.730 2013.090 1828.910 2014.270 ;
        RECT 1829.330 2013.090 1830.510 2014.270 ;
        RECT 1827.730 1834.690 1828.910 1835.870 ;
        RECT 1829.330 1834.690 1830.510 1835.870 ;
        RECT 1827.730 1833.090 1828.910 1834.270 ;
        RECT 1829.330 1833.090 1830.510 1834.270 ;
        RECT 1827.730 1654.690 1828.910 1655.870 ;
        RECT 1829.330 1654.690 1830.510 1655.870 ;
        RECT 1827.730 1653.090 1828.910 1654.270 ;
        RECT 1829.330 1653.090 1830.510 1654.270 ;
        RECT 1827.730 1474.690 1828.910 1475.870 ;
        RECT 1829.330 1474.690 1830.510 1475.870 ;
        RECT 1827.730 1473.090 1828.910 1474.270 ;
        RECT 1829.330 1473.090 1830.510 1474.270 ;
        RECT 1827.730 1294.690 1828.910 1295.870 ;
        RECT 1829.330 1294.690 1830.510 1295.870 ;
        RECT 1827.730 1293.090 1828.910 1294.270 ;
        RECT 1829.330 1293.090 1830.510 1294.270 ;
        RECT 1827.730 1114.690 1828.910 1115.870 ;
        RECT 1829.330 1114.690 1830.510 1115.870 ;
        RECT 1827.730 1113.090 1828.910 1114.270 ;
        RECT 1829.330 1113.090 1830.510 1114.270 ;
        RECT 1827.730 934.690 1828.910 935.870 ;
        RECT 1829.330 934.690 1830.510 935.870 ;
        RECT 1827.730 933.090 1828.910 934.270 ;
        RECT 1829.330 933.090 1830.510 934.270 ;
        RECT 1827.730 754.690 1828.910 755.870 ;
        RECT 1829.330 754.690 1830.510 755.870 ;
        RECT 1827.730 753.090 1828.910 754.270 ;
        RECT 1829.330 753.090 1830.510 754.270 ;
        RECT 1827.730 574.690 1828.910 575.870 ;
        RECT 1829.330 574.690 1830.510 575.870 ;
        RECT 1827.730 573.090 1828.910 574.270 ;
        RECT 1829.330 573.090 1830.510 574.270 ;
        RECT 1827.730 394.690 1828.910 395.870 ;
        RECT 1829.330 394.690 1830.510 395.870 ;
        RECT 1827.730 393.090 1828.910 394.270 ;
        RECT 1829.330 393.090 1830.510 394.270 ;
        RECT 1827.730 214.690 1828.910 215.870 ;
        RECT 1829.330 214.690 1830.510 215.870 ;
        RECT 1827.730 213.090 1828.910 214.270 ;
        RECT 1829.330 213.090 1830.510 214.270 ;
        RECT 1827.730 34.690 1828.910 35.870 ;
        RECT 1829.330 34.690 1830.510 35.870 ;
        RECT 1827.730 33.090 1828.910 34.270 ;
        RECT 1829.330 33.090 1830.510 34.270 ;
        RECT 1827.730 -12.510 1828.910 -11.330 ;
        RECT 1829.330 -12.510 1830.510 -11.330 ;
        RECT 1827.730 -14.110 1828.910 -12.930 ;
        RECT 1829.330 -14.110 1830.510 -12.930 ;
        RECT 2007.730 3532.610 2008.910 3533.790 ;
        RECT 2009.330 3532.610 2010.510 3533.790 ;
        RECT 2007.730 3531.010 2008.910 3532.190 ;
        RECT 2009.330 3531.010 2010.510 3532.190 ;
        RECT 2007.730 3454.690 2008.910 3455.870 ;
        RECT 2009.330 3454.690 2010.510 3455.870 ;
        RECT 2007.730 3453.090 2008.910 3454.270 ;
        RECT 2009.330 3453.090 2010.510 3454.270 ;
        RECT 2007.730 3274.690 2008.910 3275.870 ;
        RECT 2009.330 3274.690 2010.510 3275.870 ;
        RECT 2007.730 3273.090 2008.910 3274.270 ;
        RECT 2009.330 3273.090 2010.510 3274.270 ;
        RECT 2007.730 3094.690 2008.910 3095.870 ;
        RECT 2009.330 3094.690 2010.510 3095.870 ;
        RECT 2007.730 3093.090 2008.910 3094.270 ;
        RECT 2009.330 3093.090 2010.510 3094.270 ;
        RECT 2007.730 2914.690 2008.910 2915.870 ;
        RECT 2009.330 2914.690 2010.510 2915.870 ;
        RECT 2007.730 2913.090 2008.910 2914.270 ;
        RECT 2009.330 2913.090 2010.510 2914.270 ;
        RECT 2007.730 2734.690 2008.910 2735.870 ;
        RECT 2009.330 2734.690 2010.510 2735.870 ;
        RECT 2007.730 2733.090 2008.910 2734.270 ;
        RECT 2009.330 2733.090 2010.510 2734.270 ;
        RECT 2007.730 2554.690 2008.910 2555.870 ;
        RECT 2009.330 2554.690 2010.510 2555.870 ;
        RECT 2007.730 2553.090 2008.910 2554.270 ;
        RECT 2009.330 2553.090 2010.510 2554.270 ;
        RECT 2007.730 2374.690 2008.910 2375.870 ;
        RECT 2009.330 2374.690 2010.510 2375.870 ;
        RECT 2007.730 2373.090 2008.910 2374.270 ;
        RECT 2009.330 2373.090 2010.510 2374.270 ;
        RECT 2007.730 2194.690 2008.910 2195.870 ;
        RECT 2009.330 2194.690 2010.510 2195.870 ;
        RECT 2007.730 2193.090 2008.910 2194.270 ;
        RECT 2009.330 2193.090 2010.510 2194.270 ;
        RECT 2007.730 2014.690 2008.910 2015.870 ;
        RECT 2009.330 2014.690 2010.510 2015.870 ;
        RECT 2007.730 2013.090 2008.910 2014.270 ;
        RECT 2009.330 2013.090 2010.510 2014.270 ;
        RECT 2007.730 1834.690 2008.910 1835.870 ;
        RECT 2009.330 1834.690 2010.510 1835.870 ;
        RECT 2007.730 1833.090 2008.910 1834.270 ;
        RECT 2009.330 1833.090 2010.510 1834.270 ;
        RECT 2007.730 1654.690 2008.910 1655.870 ;
        RECT 2009.330 1654.690 2010.510 1655.870 ;
        RECT 2007.730 1653.090 2008.910 1654.270 ;
        RECT 2009.330 1653.090 2010.510 1654.270 ;
        RECT 2007.730 1474.690 2008.910 1475.870 ;
        RECT 2009.330 1474.690 2010.510 1475.870 ;
        RECT 2007.730 1473.090 2008.910 1474.270 ;
        RECT 2009.330 1473.090 2010.510 1474.270 ;
        RECT 2007.730 1294.690 2008.910 1295.870 ;
        RECT 2009.330 1294.690 2010.510 1295.870 ;
        RECT 2007.730 1293.090 2008.910 1294.270 ;
        RECT 2009.330 1293.090 2010.510 1294.270 ;
        RECT 2007.730 1114.690 2008.910 1115.870 ;
        RECT 2009.330 1114.690 2010.510 1115.870 ;
        RECT 2007.730 1113.090 2008.910 1114.270 ;
        RECT 2009.330 1113.090 2010.510 1114.270 ;
        RECT 2007.730 934.690 2008.910 935.870 ;
        RECT 2009.330 934.690 2010.510 935.870 ;
        RECT 2007.730 933.090 2008.910 934.270 ;
        RECT 2009.330 933.090 2010.510 934.270 ;
        RECT 2007.730 754.690 2008.910 755.870 ;
        RECT 2009.330 754.690 2010.510 755.870 ;
        RECT 2007.730 753.090 2008.910 754.270 ;
        RECT 2009.330 753.090 2010.510 754.270 ;
        RECT 2007.730 574.690 2008.910 575.870 ;
        RECT 2009.330 574.690 2010.510 575.870 ;
        RECT 2007.730 573.090 2008.910 574.270 ;
        RECT 2009.330 573.090 2010.510 574.270 ;
        RECT 2007.730 394.690 2008.910 395.870 ;
        RECT 2009.330 394.690 2010.510 395.870 ;
        RECT 2007.730 393.090 2008.910 394.270 ;
        RECT 2009.330 393.090 2010.510 394.270 ;
        RECT 2007.730 214.690 2008.910 215.870 ;
        RECT 2009.330 214.690 2010.510 215.870 ;
        RECT 2007.730 213.090 2008.910 214.270 ;
        RECT 2009.330 213.090 2010.510 214.270 ;
        RECT 2007.730 34.690 2008.910 35.870 ;
        RECT 2009.330 34.690 2010.510 35.870 ;
        RECT 2007.730 33.090 2008.910 34.270 ;
        RECT 2009.330 33.090 2010.510 34.270 ;
        RECT 2007.730 -12.510 2008.910 -11.330 ;
        RECT 2009.330 -12.510 2010.510 -11.330 ;
        RECT 2007.730 -14.110 2008.910 -12.930 ;
        RECT 2009.330 -14.110 2010.510 -12.930 ;
        RECT 2187.730 3532.610 2188.910 3533.790 ;
        RECT 2189.330 3532.610 2190.510 3533.790 ;
        RECT 2187.730 3531.010 2188.910 3532.190 ;
        RECT 2189.330 3531.010 2190.510 3532.190 ;
        RECT 2187.730 3454.690 2188.910 3455.870 ;
        RECT 2189.330 3454.690 2190.510 3455.870 ;
        RECT 2187.730 3453.090 2188.910 3454.270 ;
        RECT 2189.330 3453.090 2190.510 3454.270 ;
        RECT 2187.730 3274.690 2188.910 3275.870 ;
        RECT 2189.330 3274.690 2190.510 3275.870 ;
        RECT 2187.730 3273.090 2188.910 3274.270 ;
        RECT 2189.330 3273.090 2190.510 3274.270 ;
        RECT 2187.730 3094.690 2188.910 3095.870 ;
        RECT 2189.330 3094.690 2190.510 3095.870 ;
        RECT 2187.730 3093.090 2188.910 3094.270 ;
        RECT 2189.330 3093.090 2190.510 3094.270 ;
        RECT 2187.730 2914.690 2188.910 2915.870 ;
        RECT 2189.330 2914.690 2190.510 2915.870 ;
        RECT 2187.730 2913.090 2188.910 2914.270 ;
        RECT 2189.330 2913.090 2190.510 2914.270 ;
        RECT 2187.730 2734.690 2188.910 2735.870 ;
        RECT 2189.330 2734.690 2190.510 2735.870 ;
        RECT 2187.730 2733.090 2188.910 2734.270 ;
        RECT 2189.330 2733.090 2190.510 2734.270 ;
        RECT 2187.730 2554.690 2188.910 2555.870 ;
        RECT 2189.330 2554.690 2190.510 2555.870 ;
        RECT 2187.730 2553.090 2188.910 2554.270 ;
        RECT 2189.330 2553.090 2190.510 2554.270 ;
        RECT 2187.730 2374.690 2188.910 2375.870 ;
        RECT 2189.330 2374.690 2190.510 2375.870 ;
        RECT 2187.730 2373.090 2188.910 2374.270 ;
        RECT 2189.330 2373.090 2190.510 2374.270 ;
        RECT 2187.730 2194.690 2188.910 2195.870 ;
        RECT 2189.330 2194.690 2190.510 2195.870 ;
        RECT 2187.730 2193.090 2188.910 2194.270 ;
        RECT 2189.330 2193.090 2190.510 2194.270 ;
        RECT 2187.730 2014.690 2188.910 2015.870 ;
        RECT 2189.330 2014.690 2190.510 2015.870 ;
        RECT 2187.730 2013.090 2188.910 2014.270 ;
        RECT 2189.330 2013.090 2190.510 2014.270 ;
        RECT 2187.730 1834.690 2188.910 1835.870 ;
        RECT 2189.330 1834.690 2190.510 1835.870 ;
        RECT 2187.730 1833.090 2188.910 1834.270 ;
        RECT 2189.330 1833.090 2190.510 1834.270 ;
        RECT 2187.730 1654.690 2188.910 1655.870 ;
        RECT 2189.330 1654.690 2190.510 1655.870 ;
        RECT 2187.730 1653.090 2188.910 1654.270 ;
        RECT 2189.330 1653.090 2190.510 1654.270 ;
        RECT 2187.730 1474.690 2188.910 1475.870 ;
        RECT 2189.330 1474.690 2190.510 1475.870 ;
        RECT 2187.730 1473.090 2188.910 1474.270 ;
        RECT 2189.330 1473.090 2190.510 1474.270 ;
        RECT 2187.730 1294.690 2188.910 1295.870 ;
        RECT 2189.330 1294.690 2190.510 1295.870 ;
        RECT 2187.730 1293.090 2188.910 1294.270 ;
        RECT 2189.330 1293.090 2190.510 1294.270 ;
        RECT 2187.730 1114.690 2188.910 1115.870 ;
        RECT 2189.330 1114.690 2190.510 1115.870 ;
        RECT 2187.730 1113.090 2188.910 1114.270 ;
        RECT 2189.330 1113.090 2190.510 1114.270 ;
        RECT 2187.730 934.690 2188.910 935.870 ;
        RECT 2189.330 934.690 2190.510 935.870 ;
        RECT 2187.730 933.090 2188.910 934.270 ;
        RECT 2189.330 933.090 2190.510 934.270 ;
        RECT 2187.730 754.690 2188.910 755.870 ;
        RECT 2189.330 754.690 2190.510 755.870 ;
        RECT 2187.730 753.090 2188.910 754.270 ;
        RECT 2189.330 753.090 2190.510 754.270 ;
        RECT 2187.730 574.690 2188.910 575.870 ;
        RECT 2189.330 574.690 2190.510 575.870 ;
        RECT 2187.730 573.090 2188.910 574.270 ;
        RECT 2189.330 573.090 2190.510 574.270 ;
        RECT 2187.730 394.690 2188.910 395.870 ;
        RECT 2189.330 394.690 2190.510 395.870 ;
        RECT 2187.730 393.090 2188.910 394.270 ;
        RECT 2189.330 393.090 2190.510 394.270 ;
        RECT 2187.730 214.690 2188.910 215.870 ;
        RECT 2189.330 214.690 2190.510 215.870 ;
        RECT 2187.730 213.090 2188.910 214.270 ;
        RECT 2189.330 213.090 2190.510 214.270 ;
        RECT 2187.730 34.690 2188.910 35.870 ;
        RECT 2189.330 34.690 2190.510 35.870 ;
        RECT 2187.730 33.090 2188.910 34.270 ;
        RECT 2189.330 33.090 2190.510 34.270 ;
        RECT 2187.730 -12.510 2188.910 -11.330 ;
        RECT 2189.330 -12.510 2190.510 -11.330 ;
        RECT 2187.730 -14.110 2188.910 -12.930 ;
        RECT 2189.330 -14.110 2190.510 -12.930 ;
        RECT 2367.730 3532.610 2368.910 3533.790 ;
        RECT 2369.330 3532.610 2370.510 3533.790 ;
        RECT 2367.730 3531.010 2368.910 3532.190 ;
        RECT 2369.330 3531.010 2370.510 3532.190 ;
        RECT 2367.730 3454.690 2368.910 3455.870 ;
        RECT 2369.330 3454.690 2370.510 3455.870 ;
        RECT 2367.730 3453.090 2368.910 3454.270 ;
        RECT 2369.330 3453.090 2370.510 3454.270 ;
        RECT 2367.730 3274.690 2368.910 3275.870 ;
        RECT 2369.330 3274.690 2370.510 3275.870 ;
        RECT 2367.730 3273.090 2368.910 3274.270 ;
        RECT 2369.330 3273.090 2370.510 3274.270 ;
        RECT 2367.730 3094.690 2368.910 3095.870 ;
        RECT 2369.330 3094.690 2370.510 3095.870 ;
        RECT 2367.730 3093.090 2368.910 3094.270 ;
        RECT 2369.330 3093.090 2370.510 3094.270 ;
        RECT 2367.730 2914.690 2368.910 2915.870 ;
        RECT 2369.330 2914.690 2370.510 2915.870 ;
        RECT 2367.730 2913.090 2368.910 2914.270 ;
        RECT 2369.330 2913.090 2370.510 2914.270 ;
        RECT 2367.730 2734.690 2368.910 2735.870 ;
        RECT 2369.330 2734.690 2370.510 2735.870 ;
        RECT 2367.730 2733.090 2368.910 2734.270 ;
        RECT 2369.330 2733.090 2370.510 2734.270 ;
        RECT 2367.730 2554.690 2368.910 2555.870 ;
        RECT 2369.330 2554.690 2370.510 2555.870 ;
        RECT 2367.730 2553.090 2368.910 2554.270 ;
        RECT 2369.330 2553.090 2370.510 2554.270 ;
        RECT 2367.730 2374.690 2368.910 2375.870 ;
        RECT 2369.330 2374.690 2370.510 2375.870 ;
        RECT 2367.730 2373.090 2368.910 2374.270 ;
        RECT 2369.330 2373.090 2370.510 2374.270 ;
        RECT 2367.730 2194.690 2368.910 2195.870 ;
        RECT 2369.330 2194.690 2370.510 2195.870 ;
        RECT 2367.730 2193.090 2368.910 2194.270 ;
        RECT 2369.330 2193.090 2370.510 2194.270 ;
        RECT 2367.730 2014.690 2368.910 2015.870 ;
        RECT 2369.330 2014.690 2370.510 2015.870 ;
        RECT 2367.730 2013.090 2368.910 2014.270 ;
        RECT 2369.330 2013.090 2370.510 2014.270 ;
        RECT 2367.730 1834.690 2368.910 1835.870 ;
        RECT 2369.330 1834.690 2370.510 1835.870 ;
        RECT 2367.730 1833.090 2368.910 1834.270 ;
        RECT 2369.330 1833.090 2370.510 1834.270 ;
        RECT 2367.730 1654.690 2368.910 1655.870 ;
        RECT 2369.330 1654.690 2370.510 1655.870 ;
        RECT 2367.730 1653.090 2368.910 1654.270 ;
        RECT 2369.330 1653.090 2370.510 1654.270 ;
        RECT 2367.730 1474.690 2368.910 1475.870 ;
        RECT 2369.330 1474.690 2370.510 1475.870 ;
        RECT 2367.730 1473.090 2368.910 1474.270 ;
        RECT 2369.330 1473.090 2370.510 1474.270 ;
        RECT 2367.730 1294.690 2368.910 1295.870 ;
        RECT 2369.330 1294.690 2370.510 1295.870 ;
        RECT 2367.730 1293.090 2368.910 1294.270 ;
        RECT 2369.330 1293.090 2370.510 1294.270 ;
        RECT 2367.730 1114.690 2368.910 1115.870 ;
        RECT 2369.330 1114.690 2370.510 1115.870 ;
        RECT 2367.730 1113.090 2368.910 1114.270 ;
        RECT 2369.330 1113.090 2370.510 1114.270 ;
        RECT 2367.730 934.690 2368.910 935.870 ;
        RECT 2369.330 934.690 2370.510 935.870 ;
        RECT 2367.730 933.090 2368.910 934.270 ;
        RECT 2369.330 933.090 2370.510 934.270 ;
        RECT 2367.730 754.690 2368.910 755.870 ;
        RECT 2369.330 754.690 2370.510 755.870 ;
        RECT 2367.730 753.090 2368.910 754.270 ;
        RECT 2369.330 753.090 2370.510 754.270 ;
        RECT 2367.730 574.690 2368.910 575.870 ;
        RECT 2369.330 574.690 2370.510 575.870 ;
        RECT 2367.730 573.090 2368.910 574.270 ;
        RECT 2369.330 573.090 2370.510 574.270 ;
        RECT 2367.730 394.690 2368.910 395.870 ;
        RECT 2369.330 394.690 2370.510 395.870 ;
        RECT 2367.730 393.090 2368.910 394.270 ;
        RECT 2369.330 393.090 2370.510 394.270 ;
        RECT 2367.730 214.690 2368.910 215.870 ;
        RECT 2369.330 214.690 2370.510 215.870 ;
        RECT 2367.730 213.090 2368.910 214.270 ;
        RECT 2369.330 213.090 2370.510 214.270 ;
        RECT 2367.730 34.690 2368.910 35.870 ;
        RECT 2369.330 34.690 2370.510 35.870 ;
        RECT 2367.730 33.090 2368.910 34.270 ;
        RECT 2369.330 33.090 2370.510 34.270 ;
        RECT 2367.730 -12.510 2368.910 -11.330 ;
        RECT 2369.330 -12.510 2370.510 -11.330 ;
        RECT 2367.730 -14.110 2368.910 -12.930 ;
        RECT 2369.330 -14.110 2370.510 -12.930 ;
        RECT 2547.730 3532.610 2548.910 3533.790 ;
        RECT 2549.330 3532.610 2550.510 3533.790 ;
        RECT 2547.730 3531.010 2548.910 3532.190 ;
        RECT 2549.330 3531.010 2550.510 3532.190 ;
        RECT 2547.730 3454.690 2548.910 3455.870 ;
        RECT 2549.330 3454.690 2550.510 3455.870 ;
        RECT 2547.730 3453.090 2548.910 3454.270 ;
        RECT 2549.330 3453.090 2550.510 3454.270 ;
        RECT 2547.730 3274.690 2548.910 3275.870 ;
        RECT 2549.330 3274.690 2550.510 3275.870 ;
        RECT 2547.730 3273.090 2548.910 3274.270 ;
        RECT 2549.330 3273.090 2550.510 3274.270 ;
        RECT 2547.730 3094.690 2548.910 3095.870 ;
        RECT 2549.330 3094.690 2550.510 3095.870 ;
        RECT 2547.730 3093.090 2548.910 3094.270 ;
        RECT 2549.330 3093.090 2550.510 3094.270 ;
        RECT 2547.730 2914.690 2548.910 2915.870 ;
        RECT 2549.330 2914.690 2550.510 2915.870 ;
        RECT 2547.730 2913.090 2548.910 2914.270 ;
        RECT 2549.330 2913.090 2550.510 2914.270 ;
        RECT 2547.730 2734.690 2548.910 2735.870 ;
        RECT 2549.330 2734.690 2550.510 2735.870 ;
        RECT 2547.730 2733.090 2548.910 2734.270 ;
        RECT 2549.330 2733.090 2550.510 2734.270 ;
        RECT 2547.730 2554.690 2548.910 2555.870 ;
        RECT 2549.330 2554.690 2550.510 2555.870 ;
        RECT 2547.730 2553.090 2548.910 2554.270 ;
        RECT 2549.330 2553.090 2550.510 2554.270 ;
        RECT 2547.730 2374.690 2548.910 2375.870 ;
        RECT 2549.330 2374.690 2550.510 2375.870 ;
        RECT 2547.730 2373.090 2548.910 2374.270 ;
        RECT 2549.330 2373.090 2550.510 2374.270 ;
        RECT 2547.730 2194.690 2548.910 2195.870 ;
        RECT 2549.330 2194.690 2550.510 2195.870 ;
        RECT 2547.730 2193.090 2548.910 2194.270 ;
        RECT 2549.330 2193.090 2550.510 2194.270 ;
        RECT 2547.730 2014.690 2548.910 2015.870 ;
        RECT 2549.330 2014.690 2550.510 2015.870 ;
        RECT 2547.730 2013.090 2548.910 2014.270 ;
        RECT 2549.330 2013.090 2550.510 2014.270 ;
        RECT 2547.730 1834.690 2548.910 1835.870 ;
        RECT 2549.330 1834.690 2550.510 1835.870 ;
        RECT 2547.730 1833.090 2548.910 1834.270 ;
        RECT 2549.330 1833.090 2550.510 1834.270 ;
        RECT 2547.730 1654.690 2548.910 1655.870 ;
        RECT 2549.330 1654.690 2550.510 1655.870 ;
        RECT 2547.730 1653.090 2548.910 1654.270 ;
        RECT 2549.330 1653.090 2550.510 1654.270 ;
        RECT 2547.730 1474.690 2548.910 1475.870 ;
        RECT 2549.330 1474.690 2550.510 1475.870 ;
        RECT 2547.730 1473.090 2548.910 1474.270 ;
        RECT 2549.330 1473.090 2550.510 1474.270 ;
        RECT 2547.730 1294.690 2548.910 1295.870 ;
        RECT 2549.330 1294.690 2550.510 1295.870 ;
        RECT 2547.730 1293.090 2548.910 1294.270 ;
        RECT 2549.330 1293.090 2550.510 1294.270 ;
        RECT 2547.730 1114.690 2548.910 1115.870 ;
        RECT 2549.330 1114.690 2550.510 1115.870 ;
        RECT 2547.730 1113.090 2548.910 1114.270 ;
        RECT 2549.330 1113.090 2550.510 1114.270 ;
        RECT 2547.730 934.690 2548.910 935.870 ;
        RECT 2549.330 934.690 2550.510 935.870 ;
        RECT 2547.730 933.090 2548.910 934.270 ;
        RECT 2549.330 933.090 2550.510 934.270 ;
        RECT 2547.730 754.690 2548.910 755.870 ;
        RECT 2549.330 754.690 2550.510 755.870 ;
        RECT 2547.730 753.090 2548.910 754.270 ;
        RECT 2549.330 753.090 2550.510 754.270 ;
        RECT 2547.730 574.690 2548.910 575.870 ;
        RECT 2549.330 574.690 2550.510 575.870 ;
        RECT 2547.730 573.090 2548.910 574.270 ;
        RECT 2549.330 573.090 2550.510 574.270 ;
        RECT 2547.730 394.690 2548.910 395.870 ;
        RECT 2549.330 394.690 2550.510 395.870 ;
        RECT 2547.730 393.090 2548.910 394.270 ;
        RECT 2549.330 393.090 2550.510 394.270 ;
        RECT 2547.730 214.690 2548.910 215.870 ;
        RECT 2549.330 214.690 2550.510 215.870 ;
        RECT 2547.730 213.090 2548.910 214.270 ;
        RECT 2549.330 213.090 2550.510 214.270 ;
        RECT 2547.730 34.690 2548.910 35.870 ;
        RECT 2549.330 34.690 2550.510 35.870 ;
        RECT 2547.730 33.090 2548.910 34.270 ;
        RECT 2549.330 33.090 2550.510 34.270 ;
        RECT 2547.730 -12.510 2548.910 -11.330 ;
        RECT 2549.330 -12.510 2550.510 -11.330 ;
        RECT 2547.730 -14.110 2548.910 -12.930 ;
        RECT 2549.330 -14.110 2550.510 -12.930 ;
        RECT 2727.730 3532.610 2728.910 3533.790 ;
        RECT 2729.330 3532.610 2730.510 3533.790 ;
        RECT 2727.730 3531.010 2728.910 3532.190 ;
        RECT 2729.330 3531.010 2730.510 3532.190 ;
        RECT 2727.730 3454.690 2728.910 3455.870 ;
        RECT 2729.330 3454.690 2730.510 3455.870 ;
        RECT 2727.730 3453.090 2728.910 3454.270 ;
        RECT 2729.330 3453.090 2730.510 3454.270 ;
        RECT 2727.730 3274.690 2728.910 3275.870 ;
        RECT 2729.330 3274.690 2730.510 3275.870 ;
        RECT 2727.730 3273.090 2728.910 3274.270 ;
        RECT 2729.330 3273.090 2730.510 3274.270 ;
        RECT 2727.730 3094.690 2728.910 3095.870 ;
        RECT 2729.330 3094.690 2730.510 3095.870 ;
        RECT 2727.730 3093.090 2728.910 3094.270 ;
        RECT 2729.330 3093.090 2730.510 3094.270 ;
        RECT 2727.730 2914.690 2728.910 2915.870 ;
        RECT 2729.330 2914.690 2730.510 2915.870 ;
        RECT 2727.730 2913.090 2728.910 2914.270 ;
        RECT 2729.330 2913.090 2730.510 2914.270 ;
        RECT 2727.730 2734.690 2728.910 2735.870 ;
        RECT 2729.330 2734.690 2730.510 2735.870 ;
        RECT 2727.730 2733.090 2728.910 2734.270 ;
        RECT 2729.330 2733.090 2730.510 2734.270 ;
        RECT 2727.730 2554.690 2728.910 2555.870 ;
        RECT 2729.330 2554.690 2730.510 2555.870 ;
        RECT 2727.730 2553.090 2728.910 2554.270 ;
        RECT 2729.330 2553.090 2730.510 2554.270 ;
        RECT 2727.730 2374.690 2728.910 2375.870 ;
        RECT 2729.330 2374.690 2730.510 2375.870 ;
        RECT 2727.730 2373.090 2728.910 2374.270 ;
        RECT 2729.330 2373.090 2730.510 2374.270 ;
        RECT 2727.730 2194.690 2728.910 2195.870 ;
        RECT 2729.330 2194.690 2730.510 2195.870 ;
        RECT 2727.730 2193.090 2728.910 2194.270 ;
        RECT 2729.330 2193.090 2730.510 2194.270 ;
        RECT 2727.730 2014.690 2728.910 2015.870 ;
        RECT 2729.330 2014.690 2730.510 2015.870 ;
        RECT 2727.730 2013.090 2728.910 2014.270 ;
        RECT 2729.330 2013.090 2730.510 2014.270 ;
        RECT 2727.730 1834.690 2728.910 1835.870 ;
        RECT 2729.330 1834.690 2730.510 1835.870 ;
        RECT 2727.730 1833.090 2728.910 1834.270 ;
        RECT 2729.330 1833.090 2730.510 1834.270 ;
        RECT 2727.730 1654.690 2728.910 1655.870 ;
        RECT 2729.330 1654.690 2730.510 1655.870 ;
        RECT 2727.730 1653.090 2728.910 1654.270 ;
        RECT 2729.330 1653.090 2730.510 1654.270 ;
        RECT 2727.730 1474.690 2728.910 1475.870 ;
        RECT 2729.330 1474.690 2730.510 1475.870 ;
        RECT 2727.730 1473.090 2728.910 1474.270 ;
        RECT 2729.330 1473.090 2730.510 1474.270 ;
        RECT 2727.730 1294.690 2728.910 1295.870 ;
        RECT 2729.330 1294.690 2730.510 1295.870 ;
        RECT 2727.730 1293.090 2728.910 1294.270 ;
        RECT 2729.330 1293.090 2730.510 1294.270 ;
        RECT 2727.730 1114.690 2728.910 1115.870 ;
        RECT 2729.330 1114.690 2730.510 1115.870 ;
        RECT 2727.730 1113.090 2728.910 1114.270 ;
        RECT 2729.330 1113.090 2730.510 1114.270 ;
        RECT 2727.730 934.690 2728.910 935.870 ;
        RECT 2729.330 934.690 2730.510 935.870 ;
        RECT 2727.730 933.090 2728.910 934.270 ;
        RECT 2729.330 933.090 2730.510 934.270 ;
        RECT 2727.730 754.690 2728.910 755.870 ;
        RECT 2729.330 754.690 2730.510 755.870 ;
        RECT 2727.730 753.090 2728.910 754.270 ;
        RECT 2729.330 753.090 2730.510 754.270 ;
        RECT 2727.730 574.690 2728.910 575.870 ;
        RECT 2729.330 574.690 2730.510 575.870 ;
        RECT 2727.730 573.090 2728.910 574.270 ;
        RECT 2729.330 573.090 2730.510 574.270 ;
        RECT 2727.730 394.690 2728.910 395.870 ;
        RECT 2729.330 394.690 2730.510 395.870 ;
        RECT 2727.730 393.090 2728.910 394.270 ;
        RECT 2729.330 393.090 2730.510 394.270 ;
        RECT 2727.730 214.690 2728.910 215.870 ;
        RECT 2729.330 214.690 2730.510 215.870 ;
        RECT 2727.730 213.090 2728.910 214.270 ;
        RECT 2729.330 213.090 2730.510 214.270 ;
        RECT 2727.730 34.690 2728.910 35.870 ;
        RECT 2729.330 34.690 2730.510 35.870 ;
        RECT 2727.730 33.090 2728.910 34.270 ;
        RECT 2729.330 33.090 2730.510 34.270 ;
        RECT 2727.730 -12.510 2728.910 -11.330 ;
        RECT 2729.330 -12.510 2730.510 -11.330 ;
        RECT 2727.730 -14.110 2728.910 -12.930 ;
        RECT 2729.330 -14.110 2730.510 -12.930 ;
        RECT 2907.730 3532.610 2908.910 3533.790 ;
        RECT 2909.330 3532.610 2910.510 3533.790 ;
        RECT 2907.730 3531.010 2908.910 3532.190 ;
        RECT 2909.330 3531.010 2910.510 3532.190 ;
        RECT 2907.730 3454.690 2908.910 3455.870 ;
        RECT 2909.330 3454.690 2910.510 3455.870 ;
        RECT 2907.730 3453.090 2908.910 3454.270 ;
        RECT 2909.330 3453.090 2910.510 3454.270 ;
        RECT 2907.730 3274.690 2908.910 3275.870 ;
        RECT 2909.330 3274.690 2910.510 3275.870 ;
        RECT 2907.730 3273.090 2908.910 3274.270 ;
        RECT 2909.330 3273.090 2910.510 3274.270 ;
        RECT 2907.730 3094.690 2908.910 3095.870 ;
        RECT 2909.330 3094.690 2910.510 3095.870 ;
        RECT 2907.730 3093.090 2908.910 3094.270 ;
        RECT 2909.330 3093.090 2910.510 3094.270 ;
        RECT 2907.730 2914.690 2908.910 2915.870 ;
        RECT 2909.330 2914.690 2910.510 2915.870 ;
        RECT 2907.730 2913.090 2908.910 2914.270 ;
        RECT 2909.330 2913.090 2910.510 2914.270 ;
        RECT 2907.730 2734.690 2908.910 2735.870 ;
        RECT 2909.330 2734.690 2910.510 2735.870 ;
        RECT 2907.730 2733.090 2908.910 2734.270 ;
        RECT 2909.330 2733.090 2910.510 2734.270 ;
        RECT 2907.730 2554.690 2908.910 2555.870 ;
        RECT 2909.330 2554.690 2910.510 2555.870 ;
        RECT 2907.730 2553.090 2908.910 2554.270 ;
        RECT 2909.330 2553.090 2910.510 2554.270 ;
        RECT 2907.730 2374.690 2908.910 2375.870 ;
        RECT 2909.330 2374.690 2910.510 2375.870 ;
        RECT 2907.730 2373.090 2908.910 2374.270 ;
        RECT 2909.330 2373.090 2910.510 2374.270 ;
        RECT 2907.730 2194.690 2908.910 2195.870 ;
        RECT 2909.330 2194.690 2910.510 2195.870 ;
        RECT 2907.730 2193.090 2908.910 2194.270 ;
        RECT 2909.330 2193.090 2910.510 2194.270 ;
        RECT 2907.730 2014.690 2908.910 2015.870 ;
        RECT 2909.330 2014.690 2910.510 2015.870 ;
        RECT 2907.730 2013.090 2908.910 2014.270 ;
        RECT 2909.330 2013.090 2910.510 2014.270 ;
        RECT 2907.730 1834.690 2908.910 1835.870 ;
        RECT 2909.330 1834.690 2910.510 1835.870 ;
        RECT 2907.730 1833.090 2908.910 1834.270 ;
        RECT 2909.330 1833.090 2910.510 1834.270 ;
        RECT 2907.730 1654.690 2908.910 1655.870 ;
        RECT 2909.330 1654.690 2910.510 1655.870 ;
        RECT 2907.730 1653.090 2908.910 1654.270 ;
        RECT 2909.330 1653.090 2910.510 1654.270 ;
        RECT 2907.730 1474.690 2908.910 1475.870 ;
        RECT 2909.330 1474.690 2910.510 1475.870 ;
        RECT 2907.730 1473.090 2908.910 1474.270 ;
        RECT 2909.330 1473.090 2910.510 1474.270 ;
        RECT 2907.730 1294.690 2908.910 1295.870 ;
        RECT 2909.330 1294.690 2910.510 1295.870 ;
        RECT 2907.730 1293.090 2908.910 1294.270 ;
        RECT 2909.330 1293.090 2910.510 1294.270 ;
        RECT 2907.730 1114.690 2908.910 1115.870 ;
        RECT 2909.330 1114.690 2910.510 1115.870 ;
        RECT 2907.730 1113.090 2908.910 1114.270 ;
        RECT 2909.330 1113.090 2910.510 1114.270 ;
        RECT 2907.730 934.690 2908.910 935.870 ;
        RECT 2909.330 934.690 2910.510 935.870 ;
        RECT 2907.730 933.090 2908.910 934.270 ;
        RECT 2909.330 933.090 2910.510 934.270 ;
        RECT 2907.730 754.690 2908.910 755.870 ;
        RECT 2909.330 754.690 2910.510 755.870 ;
        RECT 2907.730 753.090 2908.910 754.270 ;
        RECT 2909.330 753.090 2910.510 754.270 ;
        RECT 2907.730 574.690 2908.910 575.870 ;
        RECT 2909.330 574.690 2910.510 575.870 ;
        RECT 2907.730 573.090 2908.910 574.270 ;
        RECT 2909.330 573.090 2910.510 574.270 ;
        RECT 2907.730 394.690 2908.910 395.870 ;
        RECT 2909.330 394.690 2910.510 395.870 ;
        RECT 2907.730 393.090 2908.910 394.270 ;
        RECT 2909.330 393.090 2910.510 394.270 ;
        RECT 2907.730 214.690 2908.910 215.870 ;
        RECT 2909.330 214.690 2910.510 215.870 ;
        RECT 2907.730 213.090 2908.910 214.270 ;
        RECT 2909.330 213.090 2910.510 214.270 ;
        RECT 2907.730 34.690 2908.910 35.870 ;
        RECT 2909.330 34.690 2910.510 35.870 ;
        RECT 2907.730 33.090 2908.910 34.270 ;
        RECT 2909.330 33.090 2910.510 34.270 ;
        RECT 2907.730 -12.510 2908.910 -11.330 ;
        RECT 2909.330 -12.510 2910.510 -11.330 ;
        RECT 2907.730 -14.110 2908.910 -12.930 ;
        RECT 2909.330 -14.110 2910.510 -12.930 ;
        RECT 2936.310 3532.610 2937.490 3533.790 ;
        RECT 2937.910 3532.610 2939.090 3533.790 ;
        RECT 2936.310 3531.010 2937.490 3532.190 ;
        RECT 2937.910 3531.010 2939.090 3532.190 ;
        RECT 2936.310 3454.690 2937.490 3455.870 ;
        RECT 2937.910 3454.690 2939.090 3455.870 ;
        RECT 2936.310 3453.090 2937.490 3454.270 ;
        RECT 2937.910 3453.090 2939.090 3454.270 ;
        RECT 2936.310 3274.690 2937.490 3275.870 ;
        RECT 2937.910 3274.690 2939.090 3275.870 ;
        RECT 2936.310 3273.090 2937.490 3274.270 ;
        RECT 2937.910 3273.090 2939.090 3274.270 ;
        RECT 2936.310 3094.690 2937.490 3095.870 ;
        RECT 2937.910 3094.690 2939.090 3095.870 ;
        RECT 2936.310 3093.090 2937.490 3094.270 ;
        RECT 2937.910 3093.090 2939.090 3094.270 ;
        RECT 2936.310 2914.690 2937.490 2915.870 ;
        RECT 2937.910 2914.690 2939.090 2915.870 ;
        RECT 2936.310 2913.090 2937.490 2914.270 ;
        RECT 2937.910 2913.090 2939.090 2914.270 ;
        RECT 2936.310 2734.690 2937.490 2735.870 ;
        RECT 2937.910 2734.690 2939.090 2735.870 ;
        RECT 2936.310 2733.090 2937.490 2734.270 ;
        RECT 2937.910 2733.090 2939.090 2734.270 ;
        RECT 2936.310 2554.690 2937.490 2555.870 ;
        RECT 2937.910 2554.690 2939.090 2555.870 ;
        RECT 2936.310 2553.090 2937.490 2554.270 ;
        RECT 2937.910 2553.090 2939.090 2554.270 ;
        RECT 2936.310 2374.690 2937.490 2375.870 ;
        RECT 2937.910 2374.690 2939.090 2375.870 ;
        RECT 2936.310 2373.090 2937.490 2374.270 ;
        RECT 2937.910 2373.090 2939.090 2374.270 ;
        RECT 2936.310 2194.690 2937.490 2195.870 ;
        RECT 2937.910 2194.690 2939.090 2195.870 ;
        RECT 2936.310 2193.090 2937.490 2194.270 ;
        RECT 2937.910 2193.090 2939.090 2194.270 ;
        RECT 2936.310 2014.690 2937.490 2015.870 ;
        RECT 2937.910 2014.690 2939.090 2015.870 ;
        RECT 2936.310 2013.090 2937.490 2014.270 ;
        RECT 2937.910 2013.090 2939.090 2014.270 ;
        RECT 2936.310 1834.690 2937.490 1835.870 ;
        RECT 2937.910 1834.690 2939.090 1835.870 ;
        RECT 2936.310 1833.090 2937.490 1834.270 ;
        RECT 2937.910 1833.090 2939.090 1834.270 ;
        RECT 2936.310 1654.690 2937.490 1655.870 ;
        RECT 2937.910 1654.690 2939.090 1655.870 ;
        RECT 2936.310 1653.090 2937.490 1654.270 ;
        RECT 2937.910 1653.090 2939.090 1654.270 ;
        RECT 2936.310 1474.690 2937.490 1475.870 ;
        RECT 2937.910 1474.690 2939.090 1475.870 ;
        RECT 2936.310 1473.090 2937.490 1474.270 ;
        RECT 2937.910 1473.090 2939.090 1474.270 ;
        RECT 2936.310 1294.690 2937.490 1295.870 ;
        RECT 2937.910 1294.690 2939.090 1295.870 ;
        RECT 2936.310 1293.090 2937.490 1294.270 ;
        RECT 2937.910 1293.090 2939.090 1294.270 ;
        RECT 2936.310 1114.690 2937.490 1115.870 ;
        RECT 2937.910 1114.690 2939.090 1115.870 ;
        RECT 2936.310 1113.090 2937.490 1114.270 ;
        RECT 2937.910 1113.090 2939.090 1114.270 ;
        RECT 2936.310 934.690 2937.490 935.870 ;
        RECT 2937.910 934.690 2939.090 935.870 ;
        RECT 2936.310 933.090 2937.490 934.270 ;
        RECT 2937.910 933.090 2939.090 934.270 ;
        RECT 2936.310 754.690 2937.490 755.870 ;
        RECT 2937.910 754.690 2939.090 755.870 ;
        RECT 2936.310 753.090 2937.490 754.270 ;
        RECT 2937.910 753.090 2939.090 754.270 ;
        RECT 2936.310 574.690 2937.490 575.870 ;
        RECT 2937.910 574.690 2939.090 575.870 ;
        RECT 2936.310 573.090 2937.490 574.270 ;
        RECT 2937.910 573.090 2939.090 574.270 ;
        RECT 2936.310 394.690 2937.490 395.870 ;
        RECT 2937.910 394.690 2939.090 395.870 ;
        RECT 2936.310 393.090 2937.490 394.270 ;
        RECT 2937.910 393.090 2939.090 394.270 ;
        RECT 2936.310 214.690 2937.490 215.870 ;
        RECT 2937.910 214.690 2939.090 215.870 ;
        RECT 2936.310 213.090 2937.490 214.270 ;
        RECT 2937.910 213.090 2939.090 214.270 ;
        RECT 2936.310 34.690 2937.490 35.870 ;
        RECT 2937.910 34.690 2939.090 35.870 ;
        RECT 2936.310 33.090 2937.490 34.270 ;
        RECT 2937.910 33.090 2939.090 34.270 ;
        RECT 2936.310 -12.510 2937.490 -11.330 ;
        RECT 2937.910 -12.510 2939.090 -11.330 ;
        RECT 2936.310 -14.110 2937.490 -12.930 ;
        RECT 2937.910 -14.110 2939.090 -12.930 ;
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
        RECT -24.430 932.930 2944.050 936.030 ;
        RECT -24.430 752.930 2944.050 756.030 ;
        RECT -24.430 572.930 2944.050 576.030 ;
        RECT -24.430 392.930 2944.050 396.030 ;
        RECT -24.430 212.930 2944.050 216.030 ;
        RECT -24.430 32.930 2944.050 36.030 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
        RECT 226.170 1010.000 229.270 3548.350 ;
        RECT 406.170 1010.000 409.270 3548.350 ;
        RECT 586.170 1010.000 589.270 3548.350 ;
        RECT 766.170 1010.000 769.270 3548.350 ;
        RECT 946.170 1010.000 949.270 3548.350 ;
        RECT 226.170 -28.670 229.270 390.000 ;
        RECT 406.170 -28.670 409.270 390.000 ;
        RECT 586.170 -28.670 589.270 390.000 ;
        RECT 766.170 -28.670 769.270 390.000 ;
        RECT 946.170 -28.670 949.270 390.000 ;
        RECT 1126.170 -28.670 1129.270 3548.350 ;
        RECT 1306.170 -28.670 1309.270 3548.350 ;
        RECT 1486.170 -28.670 1489.270 3548.350 ;
        RECT 1666.170 -28.670 1669.270 3548.350 ;
        RECT 1846.170 -28.670 1849.270 3548.350 ;
        RECT 2026.170 -28.670 2029.270 3548.350 ;
        RECT 2206.170 -28.670 2209.270 3548.350 ;
        RECT 2386.170 -28.670 2389.270 3548.350 ;
        RECT 2566.170 -28.670 2569.270 3548.350 ;
        RECT 2746.170 -28.670 2749.270 3548.350 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
      LAYER via4 ;
        RECT -29.070 3542.210 -27.890 3543.390 ;
        RECT -27.470 3542.210 -26.290 3543.390 ;
        RECT -29.070 3540.610 -27.890 3541.790 ;
        RECT -27.470 3540.610 -26.290 3541.790 ;
        RECT -29.070 3473.290 -27.890 3474.470 ;
        RECT -27.470 3473.290 -26.290 3474.470 ;
        RECT -29.070 3471.690 -27.890 3472.870 ;
        RECT -27.470 3471.690 -26.290 3472.870 ;
        RECT -29.070 3293.290 -27.890 3294.470 ;
        RECT -27.470 3293.290 -26.290 3294.470 ;
        RECT -29.070 3291.690 -27.890 3292.870 ;
        RECT -27.470 3291.690 -26.290 3292.870 ;
        RECT -29.070 3113.290 -27.890 3114.470 ;
        RECT -27.470 3113.290 -26.290 3114.470 ;
        RECT -29.070 3111.690 -27.890 3112.870 ;
        RECT -27.470 3111.690 -26.290 3112.870 ;
        RECT -29.070 2933.290 -27.890 2934.470 ;
        RECT -27.470 2933.290 -26.290 2934.470 ;
        RECT -29.070 2931.690 -27.890 2932.870 ;
        RECT -27.470 2931.690 -26.290 2932.870 ;
        RECT -29.070 2753.290 -27.890 2754.470 ;
        RECT -27.470 2753.290 -26.290 2754.470 ;
        RECT -29.070 2751.690 -27.890 2752.870 ;
        RECT -27.470 2751.690 -26.290 2752.870 ;
        RECT -29.070 2573.290 -27.890 2574.470 ;
        RECT -27.470 2573.290 -26.290 2574.470 ;
        RECT -29.070 2571.690 -27.890 2572.870 ;
        RECT -27.470 2571.690 -26.290 2572.870 ;
        RECT -29.070 2393.290 -27.890 2394.470 ;
        RECT -27.470 2393.290 -26.290 2394.470 ;
        RECT -29.070 2391.690 -27.890 2392.870 ;
        RECT -27.470 2391.690 -26.290 2392.870 ;
        RECT -29.070 2213.290 -27.890 2214.470 ;
        RECT -27.470 2213.290 -26.290 2214.470 ;
        RECT -29.070 2211.690 -27.890 2212.870 ;
        RECT -27.470 2211.690 -26.290 2212.870 ;
        RECT -29.070 2033.290 -27.890 2034.470 ;
        RECT -27.470 2033.290 -26.290 2034.470 ;
        RECT -29.070 2031.690 -27.890 2032.870 ;
        RECT -27.470 2031.690 -26.290 2032.870 ;
        RECT -29.070 1853.290 -27.890 1854.470 ;
        RECT -27.470 1853.290 -26.290 1854.470 ;
        RECT -29.070 1851.690 -27.890 1852.870 ;
        RECT -27.470 1851.690 -26.290 1852.870 ;
        RECT -29.070 1673.290 -27.890 1674.470 ;
        RECT -27.470 1673.290 -26.290 1674.470 ;
        RECT -29.070 1671.690 -27.890 1672.870 ;
        RECT -27.470 1671.690 -26.290 1672.870 ;
        RECT -29.070 1493.290 -27.890 1494.470 ;
        RECT -27.470 1493.290 -26.290 1494.470 ;
        RECT -29.070 1491.690 -27.890 1492.870 ;
        RECT -27.470 1491.690 -26.290 1492.870 ;
        RECT -29.070 1313.290 -27.890 1314.470 ;
        RECT -27.470 1313.290 -26.290 1314.470 ;
        RECT -29.070 1311.690 -27.890 1312.870 ;
        RECT -27.470 1311.690 -26.290 1312.870 ;
        RECT -29.070 1133.290 -27.890 1134.470 ;
        RECT -27.470 1133.290 -26.290 1134.470 ;
        RECT -29.070 1131.690 -27.890 1132.870 ;
        RECT -27.470 1131.690 -26.290 1132.870 ;
        RECT -29.070 953.290 -27.890 954.470 ;
        RECT -27.470 953.290 -26.290 954.470 ;
        RECT -29.070 951.690 -27.890 952.870 ;
        RECT -27.470 951.690 -26.290 952.870 ;
        RECT -29.070 773.290 -27.890 774.470 ;
        RECT -27.470 773.290 -26.290 774.470 ;
        RECT -29.070 771.690 -27.890 772.870 ;
        RECT -27.470 771.690 -26.290 772.870 ;
        RECT -29.070 593.290 -27.890 594.470 ;
        RECT -27.470 593.290 -26.290 594.470 ;
        RECT -29.070 591.690 -27.890 592.870 ;
        RECT -27.470 591.690 -26.290 592.870 ;
        RECT -29.070 413.290 -27.890 414.470 ;
        RECT -27.470 413.290 -26.290 414.470 ;
        RECT -29.070 411.690 -27.890 412.870 ;
        RECT -27.470 411.690 -26.290 412.870 ;
        RECT -29.070 233.290 -27.890 234.470 ;
        RECT -27.470 233.290 -26.290 234.470 ;
        RECT -29.070 231.690 -27.890 232.870 ;
        RECT -27.470 231.690 -26.290 232.870 ;
        RECT -29.070 53.290 -27.890 54.470 ;
        RECT -27.470 53.290 -26.290 54.470 ;
        RECT -29.070 51.690 -27.890 52.870 ;
        RECT -27.470 51.690 -26.290 52.870 ;
        RECT -29.070 -22.110 -27.890 -20.930 ;
        RECT -27.470 -22.110 -26.290 -20.930 ;
        RECT -29.070 -23.710 -27.890 -22.530 ;
        RECT -27.470 -23.710 -26.290 -22.530 ;
        RECT 46.330 3542.210 47.510 3543.390 ;
        RECT 47.930 3542.210 49.110 3543.390 ;
        RECT 46.330 3540.610 47.510 3541.790 ;
        RECT 47.930 3540.610 49.110 3541.790 ;
        RECT 46.330 3473.290 47.510 3474.470 ;
        RECT 47.930 3473.290 49.110 3474.470 ;
        RECT 46.330 3471.690 47.510 3472.870 ;
        RECT 47.930 3471.690 49.110 3472.870 ;
        RECT 46.330 3293.290 47.510 3294.470 ;
        RECT 47.930 3293.290 49.110 3294.470 ;
        RECT 46.330 3291.690 47.510 3292.870 ;
        RECT 47.930 3291.690 49.110 3292.870 ;
        RECT 46.330 3113.290 47.510 3114.470 ;
        RECT 47.930 3113.290 49.110 3114.470 ;
        RECT 46.330 3111.690 47.510 3112.870 ;
        RECT 47.930 3111.690 49.110 3112.870 ;
        RECT 46.330 2933.290 47.510 2934.470 ;
        RECT 47.930 2933.290 49.110 2934.470 ;
        RECT 46.330 2931.690 47.510 2932.870 ;
        RECT 47.930 2931.690 49.110 2932.870 ;
        RECT 46.330 2753.290 47.510 2754.470 ;
        RECT 47.930 2753.290 49.110 2754.470 ;
        RECT 46.330 2751.690 47.510 2752.870 ;
        RECT 47.930 2751.690 49.110 2752.870 ;
        RECT 46.330 2573.290 47.510 2574.470 ;
        RECT 47.930 2573.290 49.110 2574.470 ;
        RECT 46.330 2571.690 47.510 2572.870 ;
        RECT 47.930 2571.690 49.110 2572.870 ;
        RECT 46.330 2393.290 47.510 2394.470 ;
        RECT 47.930 2393.290 49.110 2394.470 ;
        RECT 46.330 2391.690 47.510 2392.870 ;
        RECT 47.930 2391.690 49.110 2392.870 ;
        RECT 46.330 2213.290 47.510 2214.470 ;
        RECT 47.930 2213.290 49.110 2214.470 ;
        RECT 46.330 2211.690 47.510 2212.870 ;
        RECT 47.930 2211.690 49.110 2212.870 ;
        RECT 46.330 2033.290 47.510 2034.470 ;
        RECT 47.930 2033.290 49.110 2034.470 ;
        RECT 46.330 2031.690 47.510 2032.870 ;
        RECT 47.930 2031.690 49.110 2032.870 ;
        RECT 46.330 1853.290 47.510 1854.470 ;
        RECT 47.930 1853.290 49.110 1854.470 ;
        RECT 46.330 1851.690 47.510 1852.870 ;
        RECT 47.930 1851.690 49.110 1852.870 ;
        RECT 46.330 1673.290 47.510 1674.470 ;
        RECT 47.930 1673.290 49.110 1674.470 ;
        RECT 46.330 1671.690 47.510 1672.870 ;
        RECT 47.930 1671.690 49.110 1672.870 ;
        RECT 46.330 1493.290 47.510 1494.470 ;
        RECT 47.930 1493.290 49.110 1494.470 ;
        RECT 46.330 1491.690 47.510 1492.870 ;
        RECT 47.930 1491.690 49.110 1492.870 ;
        RECT 46.330 1313.290 47.510 1314.470 ;
        RECT 47.930 1313.290 49.110 1314.470 ;
        RECT 46.330 1311.690 47.510 1312.870 ;
        RECT 47.930 1311.690 49.110 1312.870 ;
        RECT 46.330 1133.290 47.510 1134.470 ;
        RECT 47.930 1133.290 49.110 1134.470 ;
        RECT 46.330 1131.690 47.510 1132.870 ;
        RECT 47.930 1131.690 49.110 1132.870 ;
        RECT 226.330 3542.210 227.510 3543.390 ;
        RECT 227.930 3542.210 229.110 3543.390 ;
        RECT 226.330 3540.610 227.510 3541.790 ;
        RECT 227.930 3540.610 229.110 3541.790 ;
        RECT 226.330 3473.290 227.510 3474.470 ;
        RECT 227.930 3473.290 229.110 3474.470 ;
        RECT 226.330 3471.690 227.510 3472.870 ;
        RECT 227.930 3471.690 229.110 3472.870 ;
        RECT 226.330 3293.290 227.510 3294.470 ;
        RECT 227.930 3293.290 229.110 3294.470 ;
        RECT 226.330 3291.690 227.510 3292.870 ;
        RECT 227.930 3291.690 229.110 3292.870 ;
        RECT 226.330 3113.290 227.510 3114.470 ;
        RECT 227.930 3113.290 229.110 3114.470 ;
        RECT 226.330 3111.690 227.510 3112.870 ;
        RECT 227.930 3111.690 229.110 3112.870 ;
        RECT 226.330 2933.290 227.510 2934.470 ;
        RECT 227.930 2933.290 229.110 2934.470 ;
        RECT 226.330 2931.690 227.510 2932.870 ;
        RECT 227.930 2931.690 229.110 2932.870 ;
        RECT 226.330 2753.290 227.510 2754.470 ;
        RECT 227.930 2753.290 229.110 2754.470 ;
        RECT 226.330 2751.690 227.510 2752.870 ;
        RECT 227.930 2751.690 229.110 2752.870 ;
        RECT 226.330 2573.290 227.510 2574.470 ;
        RECT 227.930 2573.290 229.110 2574.470 ;
        RECT 226.330 2571.690 227.510 2572.870 ;
        RECT 227.930 2571.690 229.110 2572.870 ;
        RECT 226.330 2393.290 227.510 2394.470 ;
        RECT 227.930 2393.290 229.110 2394.470 ;
        RECT 226.330 2391.690 227.510 2392.870 ;
        RECT 227.930 2391.690 229.110 2392.870 ;
        RECT 226.330 2213.290 227.510 2214.470 ;
        RECT 227.930 2213.290 229.110 2214.470 ;
        RECT 226.330 2211.690 227.510 2212.870 ;
        RECT 227.930 2211.690 229.110 2212.870 ;
        RECT 226.330 2033.290 227.510 2034.470 ;
        RECT 227.930 2033.290 229.110 2034.470 ;
        RECT 226.330 2031.690 227.510 2032.870 ;
        RECT 227.930 2031.690 229.110 2032.870 ;
        RECT 226.330 1853.290 227.510 1854.470 ;
        RECT 227.930 1853.290 229.110 1854.470 ;
        RECT 226.330 1851.690 227.510 1852.870 ;
        RECT 227.930 1851.690 229.110 1852.870 ;
        RECT 226.330 1673.290 227.510 1674.470 ;
        RECT 227.930 1673.290 229.110 1674.470 ;
        RECT 226.330 1671.690 227.510 1672.870 ;
        RECT 227.930 1671.690 229.110 1672.870 ;
        RECT 226.330 1493.290 227.510 1494.470 ;
        RECT 227.930 1493.290 229.110 1494.470 ;
        RECT 226.330 1491.690 227.510 1492.870 ;
        RECT 227.930 1491.690 229.110 1492.870 ;
        RECT 226.330 1313.290 227.510 1314.470 ;
        RECT 227.930 1313.290 229.110 1314.470 ;
        RECT 226.330 1311.690 227.510 1312.870 ;
        RECT 227.930 1311.690 229.110 1312.870 ;
        RECT 226.330 1133.290 227.510 1134.470 ;
        RECT 227.930 1133.290 229.110 1134.470 ;
        RECT 226.330 1131.690 227.510 1132.870 ;
        RECT 227.930 1131.690 229.110 1132.870 ;
        RECT 406.330 3542.210 407.510 3543.390 ;
        RECT 407.930 3542.210 409.110 3543.390 ;
        RECT 406.330 3540.610 407.510 3541.790 ;
        RECT 407.930 3540.610 409.110 3541.790 ;
        RECT 406.330 3473.290 407.510 3474.470 ;
        RECT 407.930 3473.290 409.110 3474.470 ;
        RECT 406.330 3471.690 407.510 3472.870 ;
        RECT 407.930 3471.690 409.110 3472.870 ;
        RECT 406.330 3293.290 407.510 3294.470 ;
        RECT 407.930 3293.290 409.110 3294.470 ;
        RECT 406.330 3291.690 407.510 3292.870 ;
        RECT 407.930 3291.690 409.110 3292.870 ;
        RECT 406.330 3113.290 407.510 3114.470 ;
        RECT 407.930 3113.290 409.110 3114.470 ;
        RECT 406.330 3111.690 407.510 3112.870 ;
        RECT 407.930 3111.690 409.110 3112.870 ;
        RECT 406.330 2933.290 407.510 2934.470 ;
        RECT 407.930 2933.290 409.110 2934.470 ;
        RECT 406.330 2931.690 407.510 2932.870 ;
        RECT 407.930 2931.690 409.110 2932.870 ;
        RECT 406.330 2753.290 407.510 2754.470 ;
        RECT 407.930 2753.290 409.110 2754.470 ;
        RECT 406.330 2751.690 407.510 2752.870 ;
        RECT 407.930 2751.690 409.110 2752.870 ;
        RECT 406.330 2573.290 407.510 2574.470 ;
        RECT 407.930 2573.290 409.110 2574.470 ;
        RECT 406.330 2571.690 407.510 2572.870 ;
        RECT 407.930 2571.690 409.110 2572.870 ;
        RECT 406.330 2393.290 407.510 2394.470 ;
        RECT 407.930 2393.290 409.110 2394.470 ;
        RECT 406.330 2391.690 407.510 2392.870 ;
        RECT 407.930 2391.690 409.110 2392.870 ;
        RECT 406.330 2213.290 407.510 2214.470 ;
        RECT 407.930 2213.290 409.110 2214.470 ;
        RECT 406.330 2211.690 407.510 2212.870 ;
        RECT 407.930 2211.690 409.110 2212.870 ;
        RECT 406.330 2033.290 407.510 2034.470 ;
        RECT 407.930 2033.290 409.110 2034.470 ;
        RECT 406.330 2031.690 407.510 2032.870 ;
        RECT 407.930 2031.690 409.110 2032.870 ;
        RECT 406.330 1853.290 407.510 1854.470 ;
        RECT 407.930 1853.290 409.110 1854.470 ;
        RECT 406.330 1851.690 407.510 1852.870 ;
        RECT 407.930 1851.690 409.110 1852.870 ;
        RECT 406.330 1673.290 407.510 1674.470 ;
        RECT 407.930 1673.290 409.110 1674.470 ;
        RECT 406.330 1671.690 407.510 1672.870 ;
        RECT 407.930 1671.690 409.110 1672.870 ;
        RECT 406.330 1493.290 407.510 1494.470 ;
        RECT 407.930 1493.290 409.110 1494.470 ;
        RECT 406.330 1491.690 407.510 1492.870 ;
        RECT 407.930 1491.690 409.110 1492.870 ;
        RECT 406.330 1313.290 407.510 1314.470 ;
        RECT 407.930 1313.290 409.110 1314.470 ;
        RECT 406.330 1311.690 407.510 1312.870 ;
        RECT 407.930 1311.690 409.110 1312.870 ;
        RECT 406.330 1133.290 407.510 1134.470 ;
        RECT 407.930 1133.290 409.110 1134.470 ;
        RECT 406.330 1131.690 407.510 1132.870 ;
        RECT 407.930 1131.690 409.110 1132.870 ;
        RECT 586.330 3542.210 587.510 3543.390 ;
        RECT 587.930 3542.210 589.110 3543.390 ;
        RECT 586.330 3540.610 587.510 3541.790 ;
        RECT 587.930 3540.610 589.110 3541.790 ;
        RECT 586.330 3473.290 587.510 3474.470 ;
        RECT 587.930 3473.290 589.110 3474.470 ;
        RECT 586.330 3471.690 587.510 3472.870 ;
        RECT 587.930 3471.690 589.110 3472.870 ;
        RECT 586.330 3293.290 587.510 3294.470 ;
        RECT 587.930 3293.290 589.110 3294.470 ;
        RECT 586.330 3291.690 587.510 3292.870 ;
        RECT 587.930 3291.690 589.110 3292.870 ;
        RECT 586.330 3113.290 587.510 3114.470 ;
        RECT 587.930 3113.290 589.110 3114.470 ;
        RECT 586.330 3111.690 587.510 3112.870 ;
        RECT 587.930 3111.690 589.110 3112.870 ;
        RECT 586.330 2933.290 587.510 2934.470 ;
        RECT 587.930 2933.290 589.110 2934.470 ;
        RECT 586.330 2931.690 587.510 2932.870 ;
        RECT 587.930 2931.690 589.110 2932.870 ;
        RECT 586.330 2753.290 587.510 2754.470 ;
        RECT 587.930 2753.290 589.110 2754.470 ;
        RECT 586.330 2751.690 587.510 2752.870 ;
        RECT 587.930 2751.690 589.110 2752.870 ;
        RECT 586.330 2573.290 587.510 2574.470 ;
        RECT 587.930 2573.290 589.110 2574.470 ;
        RECT 586.330 2571.690 587.510 2572.870 ;
        RECT 587.930 2571.690 589.110 2572.870 ;
        RECT 586.330 2393.290 587.510 2394.470 ;
        RECT 587.930 2393.290 589.110 2394.470 ;
        RECT 586.330 2391.690 587.510 2392.870 ;
        RECT 587.930 2391.690 589.110 2392.870 ;
        RECT 586.330 2213.290 587.510 2214.470 ;
        RECT 587.930 2213.290 589.110 2214.470 ;
        RECT 586.330 2211.690 587.510 2212.870 ;
        RECT 587.930 2211.690 589.110 2212.870 ;
        RECT 586.330 2033.290 587.510 2034.470 ;
        RECT 587.930 2033.290 589.110 2034.470 ;
        RECT 586.330 2031.690 587.510 2032.870 ;
        RECT 587.930 2031.690 589.110 2032.870 ;
        RECT 586.330 1853.290 587.510 1854.470 ;
        RECT 587.930 1853.290 589.110 1854.470 ;
        RECT 586.330 1851.690 587.510 1852.870 ;
        RECT 587.930 1851.690 589.110 1852.870 ;
        RECT 586.330 1673.290 587.510 1674.470 ;
        RECT 587.930 1673.290 589.110 1674.470 ;
        RECT 586.330 1671.690 587.510 1672.870 ;
        RECT 587.930 1671.690 589.110 1672.870 ;
        RECT 586.330 1493.290 587.510 1494.470 ;
        RECT 587.930 1493.290 589.110 1494.470 ;
        RECT 586.330 1491.690 587.510 1492.870 ;
        RECT 587.930 1491.690 589.110 1492.870 ;
        RECT 586.330 1313.290 587.510 1314.470 ;
        RECT 587.930 1313.290 589.110 1314.470 ;
        RECT 586.330 1311.690 587.510 1312.870 ;
        RECT 587.930 1311.690 589.110 1312.870 ;
        RECT 586.330 1133.290 587.510 1134.470 ;
        RECT 587.930 1133.290 589.110 1134.470 ;
        RECT 586.330 1131.690 587.510 1132.870 ;
        RECT 587.930 1131.690 589.110 1132.870 ;
        RECT 766.330 3542.210 767.510 3543.390 ;
        RECT 767.930 3542.210 769.110 3543.390 ;
        RECT 766.330 3540.610 767.510 3541.790 ;
        RECT 767.930 3540.610 769.110 3541.790 ;
        RECT 766.330 3473.290 767.510 3474.470 ;
        RECT 767.930 3473.290 769.110 3474.470 ;
        RECT 766.330 3471.690 767.510 3472.870 ;
        RECT 767.930 3471.690 769.110 3472.870 ;
        RECT 766.330 3293.290 767.510 3294.470 ;
        RECT 767.930 3293.290 769.110 3294.470 ;
        RECT 766.330 3291.690 767.510 3292.870 ;
        RECT 767.930 3291.690 769.110 3292.870 ;
        RECT 766.330 3113.290 767.510 3114.470 ;
        RECT 767.930 3113.290 769.110 3114.470 ;
        RECT 766.330 3111.690 767.510 3112.870 ;
        RECT 767.930 3111.690 769.110 3112.870 ;
        RECT 766.330 2933.290 767.510 2934.470 ;
        RECT 767.930 2933.290 769.110 2934.470 ;
        RECT 766.330 2931.690 767.510 2932.870 ;
        RECT 767.930 2931.690 769.110 2932.870 ;
        RECT 766.330 2753.290 767.510 2754.470 ;
        RECT 767.930 2753.290 769.110 2754.470 ;
        RECT 766.330 2751.690 767.510 2752.870 ;
        RECT 767.930 2751.690 769.110 2752.870 ;
        RECT 766.330 2573.290 767.510 2574.470 ;
        RECT 767.930 2573.290 769.110 2574.470 ;
        RECT 766.330 2571.690 767.510 2572.870 ;
        RECT 767.930 2571.690 769.110 2572.870 ;
        RECT 766.330 2393.290 767.510 2394.470 ;
        RECT 767.930 2393.290 769.110 2394.470 ;
        RECT 766.330 2391.690 767.510 2392.870 ;
        RECT 767.930 2391.690 769.110 2392.870 ;
        RECT 766.330 2213.290 767.510 2214.470 ;
        RECT 767.930 2213.290 769.110 2214.470 ;
        RECT 766.330 2211.690 767.510 2212.870 ;
        RECT 767.930 2211.690 769.110 2212.870 ;
        RECT 766.330 2033.290 767.510 2034.470 ;
        RECT 767.930 2033.290 769.110 2034.470 ;
        RECT 766.330 2031.690 767.510 2032.870 ;
        RECT 767.930 2031.690 769.110 2032.870 ;
        RECT 766.330 1853.290 767.510 1854.470 ;
        RECT 767.930 1853.290 769.110 1854.470 ;
        RECT 766.330 1851.690 767.510 1852.870 ;
        RECT 767.930 1851.690 769.110 1852.870 ;
        RECT 766.330 1673.290 767.510 1674.470 ;
        RECT 767.930 1673.290 769.110 1674.470 ;
        RECT 766.330 1671.690 767.510 1672.870 ;
        RECT 767.930 1671.690 769.110 1672.870 ;
        RECT 766.330 1493.290 767.510 1494.470 ;
        RECT 767.930 1493.290 769.110 1494.470 ;
        RECT 766.330 1491.690 767.510 1492.870 ;
        RECT 767.930 1491.690 769.110 1492.870 ;
        RECT 766.330 1313.290 767.510 1314.470 ;
        RECT 767.930 1313.290 769.110 1314.470 ;
        RECT 766.330 1311.690 767.510 1312.870 ;
        RECT 767.930 1311.690 769.110 1312.870 ;
        RECT 766.330 1133.290 767.510 1134.470 ;
        RECT 767.930 1133.290 769.110 1134.470 ;
        RECT 766.330 1131.690 767.510 1132.870 ;
        RECT 767.930 1131.690 769.110 1132.870 ;
        RECT 946.330 3542.210 947.510 3543.390 ;
        RECT 947.930 3542.210 949.110 3543.390 ;
        RECT 946.330 3540.610 947.510 3541.790 ;
        RECT 947.930 3540.610 949.110 3541.790 ;
        RECT 946.330 3473.290 947.510 3474.470 ;
        RECT 947.930 3473.290 949.110 3474.470 ;
        RECT 946.330 3471.690 947.510 3472.870 ;
        RECT 947.930 3471.690 949.110 3472.870 ;
        RECT 946.330 3293.290 947.510 3294.470 ;
        RECT 947.930 3293.290 949.110 3294.470 ;
        RECT 946.330 3291.690 947.510 3292.870 ;
        RECT 947.930 3291.690 949.110 3292.870 ;
        RECT 946.330 3113.290 947.510 3114.470 ;
        RECT 947.930 3113.290 949.110 3114.470 ;
        RECT 946.330 3111.690 947.510 3112.870 ;
        RECT 947.930 3111.690 949.110 3112.870 ;
        RECT 946.330 2933.290 947.510 2934.470 ;
        RECT 947.930 2933.290 949.110 2934.470 ;
        RECT 946.330 2931.690 947.510 2932.870 ;
        RECT 947.930 2931.690 949.110 2932.870 ;
        RECT 946.330 2753.290 947.510 2754.470 ;
        RECT 947.930 2753.290 949.110 2754.470 ;
        RECT 946.330 2751.690 947.510 2752.870 ;
        RECT 947.930 2751.690 949.110 2752.870 ;
        RECT 946.330 2573.290 947.510 2574.470 ;
        RECT 947.930 2573.290 949.110 2574.470 ;
        RECT 946.330 2571.690 947.510 2572.870 ;
        RECT 947.930 2571.690 949.110 2572.870 ;
        RECT 946.330 2393.290 947.510 2394.470 ;
        RECT 947.930 2393.290 949.110 2394.470 ;
        RECT 946.330 2391.690 947.510 2392.870 ;
        RECT 947.930 2391.690 949.110 2392.870 ;
        RECT 946.330 2213.290 947.510 2214.470 ;
        RECT 947.930 2213.290 949.110 2214.470 ;
        RECT 946.330 2211.690 947.510 2212.870 ;
        RECT 947.930 2211.690 949.110 2212.870 ;
        RECT 946.330 2033.290 947.510 2034.470 ;
        RECT 947.930 2033.290 949.110 2034.470 ;
        RECT 946.330 2031.690 947.510 2032.870 ;
        RECT 947.930 2031.690 949.110 2032.870 ;
        RECT 946.330 1853.290 947.510 1854.470 ;
        RECT 947.930 1853.290 949.110 1854.470 ;
        RECT 946.330 1851.690 947.510 1852.870 ;
        RECT 947.930 1851.690 949.110 1852.870 ;
        RECT 946.330 1673.290 947.510 1674.470 ;
        RECT 947.930 1673.290 949.110 1674.470 ;
        RECT 946.330 1671.690 947.510 1672.870 ;
        RECT 947.930 1671.690 949.110 1672.870 ;
        RECT 946.330 1493.290 947.510 1494.470 ;
        RECT 947.930 1493.290 949.110 1494.470 ;
        RECT 946.330 1491.690 947.510 1492.870 ;
        RECT 947.930 1491.690 949.110 1492.870 ;
        RECT 946.330 1313.290 947.510 1314.470 ;
        RECT 947.930 1313.290 949.110 1314.470 ;
        RECT 946.330 1311.690 947.510 1312.870 ;
        RECT 947.930 1311.690 949.110 1312.870 ;
        RECT 946.330 1133.290 947.510 1134.470 ;
        RECT 947.930 1133.290 949.110 1134.470 ;
        RECT 946.330 1131.690 947.510 1132.870 ;
        RECT 947.930 1131.690 949.110 1132.870 ;
        RECT 1126.330 3542.210 1127.510 3543.390 ;
        RECT 1127.930 3542.210 1129.110 3543.390 ;
        RECT 1126.330 3540.610 1127.510 3541.790 ;
        RECT 1127.930 3540.610 1129.110 3541.790 ;
        RECT 1126.330 3473.290 1127.510 3474.470 ;
        RECT 1127.930 3473.290 1129.110 3474.470 ;
        RECT 1126.330 3471.690 1127.510 3472.870 ;
        RECT 1127.930 3471.690 1129.110 3472.870 ;
        RECT 1126.330 3293.290 1127.510 3294.470 ;
        RECT 1127.930 3293.290 1129.110 3294.470 ;
        RECT 1126.330 3291.690 1127.510 3292.870 ;
        RECT 1127.930 3291.690 1129.110 3292.870 ;
        RECT 1126.330 3113.290 1127.510 3114.470 ;
        RECT 1127.930 3113.290 1129.110 3114.470 ;
        RECT 1126.330 3111.690 1127.510 3112.870 ;
        RECT 1127.930 3111.690 1129.110 3112.870 ;
        RECT 1126.330 2933.290 1127.510 2934.470 ;
        RECT 1127.930 2933.290 1129.110 2934.470 ;
        RECT 1126.330 2931.690 1127.510 2932.870 ;
        RECT 1127.930 2931.690 1129.110 2932.870 ;
        RECT 1126.330 2753.290 1127.510 2754.470 ;
        RECT 1127.930 2753.290 1129.110 2754.470 ;
        RECT 1126.330 2751.690 1127.510 2752.870 ;
        RECT 1127.930 2751.690 1129.110 2752.870 ;
        RECT 1126.330 2573.290 1127.510 2574.470 ;
        RECT 1127.930 2573.290 1129.110 2574.470 ;
        RECT 1126.330 2571.690 1127.510 2572.870 ;
        RECT 1127.930 2571.690 1129.110 2572.870 ;
        RECT 1126.330 2393.290 1127.510 2394.470 ;
        RECT 1127.930 2393.290 1129.110 2394.470 ;
        RECT 1126.330 2391.690 1127.510 2392.870 ;
        RECT 1127.930 2391.690 1129.110 2392.870 ;
        RECT 1126.330 2213.290 1127.510 2214.470 ;
        RECT 1127.930 2213.290 1129.110 2214.470 ;
        RECT 1126.330 2211.690 1127.510 2212.870 ;
        RECT 1127.930 2211.690 1129.110 2212.870 ;
        RECT 1126.330 2033.290 1127.510 2034.470 ;
        RECT 1127.930 2033.290 1129.110 2034.470 ;
        RECT 1126.330 2031.690 1127.510 2032.870 ;
        RECT 1127.930 2031.690 1129.110 2032.870 ;
        RECT 1126.330 1853.290 1127.510 1854.470 ;
        RECT 1127.930 1853.290 1129.110 1854.470 ;
        RECT 1126.330 1851.690 1127.510 1852.870 ;
        RECT 1127.930 1851.690 1129.110 1852.870 ;
        RECT 1126.330 1673.290 1127.510 1674.470 ;
        RECT 1127.930 1673.290 1129.110 1674.470 ;
        RECT 1126.330 1671.690 1127.510 1672.870 ;
        RECT 1127.930 1671.690 1129.110 1672.870 ;
        RECT 1126.330 1493.290 1127.510 1494.470 ;
        RECT 1127.930 1493.290 1129.110 1494.470 ;
        RECT 1126.330 1491.690 1127.510 1492.870 ;
        RECT 1127.930 1491.690 1129.110 1492.870 ;
        RECT 1126.330 1313.290 1127.510 1314.470 ;
        RECT 1127.930 1313.290 1129.110 1314.470 ;
        RECT 1126.330 1311.690 1127.510 1312.870 ;
        RECT 1127.930 1311.690 1129.110 1312.870 ;
        RECT 1126.330 1133.290 1127.510 1134.470 ;
        RECT 1127.930 1133.290 1129.110 1134.470 ;
        RECT 1126.330 1131.690 1127.510 1132.870 ;
        RECT 1127.930 1131.690 1129.110 1132.870 ;
        RECT 46.330 953.290 47.510 954.470 ;
        RECT 47.930 953.290 49.110 954.470 ;
        RECT 46.330 951.690 47.510 952.870 ;
        RECT 47.930 951.690 49.110 952.870 ;
        RECT 46.330 773.290 47.510 774.470 ;
        RECT 47.930 773.290 49.110 774.470 ;
        RECT 46.330 771.690 47.510 772.870 ;
        RECT 47.930 771.690 49.110 772.870 ;
        RECT 46.330 593.290 47.510 594.470 ;
        RECT 47.930 593.290 49.110 594.470 ;
        RECT 46.330 591.690 47.510 592.870 ;
        RECT 47.930 591.690 49.110 592.870 ;
        RECT 46.330 413.290 47.510 414.470 ;
        RECT 47.930 413.290 49.110 414.470 ;
        RECT 46.330 411.690 47.510 412.870 ;
        RECT 47.930 411.690 49.110 412.870 ;
        RECT 1126.330 953.290 1127.510 954.470 ;
        RECT 1127.930 953.290 1129.110 954.470 ;
        RECT 1126.330 951.690 1127.510 952.870 ;
        RECT 1127.930 951.690 1129.110 952.870 ;
        RECT 1126.330 773.290 1127.510 774.470 ;
        RECT 1127.930 773.290 1129.110 774.470 ;
        RECT 1126.330 771.690 1127.510 772.870 ;
        RECT 1127.930 771.690 1129.110 772.870 ;
        RECT 1126.330 593.290 1127.510 594.470 ;
        RECT 1127.930 593.290 1129.110 594.470 ;
        RECT 1126.330 591.690 1127.510 592.870 ;
        RECT 1127.930 591.690 1129.110 592.870 ;
        RECT 1126.330 413.290 1127.510 414.470 ;
        RECT 1127.930 413.290 1129.110 414.470 ;
        RECT 1126.330 411.690 1127.510 412.870 ;
        RECT 1127.930 411.690 1129.110 412.870 ;
        RECT 46.330 233.290 47.510 234.470 ;
        RECT 47.930 233.290 49.110 234.470 ;
        RECT 46.330 231.690 47.510 232.870 ;
        RECT 47.930 231.690 49.110 232.870 ;
        RECT 46.330 53.290 47.510 54.470 ;
        RECT 47.930 53.290 49.110 54.470 ;
        RECT 46.330 51.690 47.510 52.870 ;
        RECT 47.930 51.690 49.110 52.870 ;
        RECT 46.330 -22.110 47.510 -20.930 ;
        RECT 47.930 -22.110 49.110 -20.930 ;
        RECT 46.330 -23.710 47.510 -22.530 ;
        RECT 47.930 -23.710 49.110 -22.530 ;
        RECT 226.330 233.290 227.510 234.470 ;
        RECT 227.930 233.290 229.110 234.470 ;
        RECT 226.330 231.690 227.510 232.870 ;
        RECT 227.930 231.690 229.110 232.870 ;
        RECT 226.330 53.290 227.510 54.470 ;
        RECT 227.930 53.290 229.110 54.470 ;
        RECT 226.330 51.690 227.510 52.870 ;
        RECT 227.930 51.690 229.110 52.870 ;
        RECT 226.330 -22.110 227.510 -20.930 ;
        RECT 227.930 -22.110 229.110 -20.930 ;
        RECT 226.330 -23.710 227.510 -22.530 ;
        RECT 227.930 -23.710 229.110 -22.530 ;
        RECT 406.330 233.290 407.510 234.470 ;
        RECT 407.930 233.290 409.110 234.470 ;
        RECT 406.330 231.690 407.510 232.870 ;
        RECT 407.930 231.690 409.110 232.870 ;
        RECT 406.330 53.290 407.510 54.470 ;
        RECT 407.930 53.290 409.110 54.470 ;
        RECT 406.330 51.690 407.510 52.870 ;
        RECT 407.930 51.690 409.110 52.870 ;
        RECT 406.330 -22.110 407.510 -20.930 ;
        RECT 407.930 -22.110 409.110 -20.930 ;
        RECT 406.330 -23.710 407.510 -22.530 ;
        RECT 407.930 -23.710 409.110 -22.530 ;
        RECT 586.330 233.290 587.510 234.470 ;
        RECT 587.930 233.290 589.110 234.470 ;
        RECT 586.330 231.690 587.510 232.870 ;
        RECT 587.930 231.690 589.110 232.870 ;
        RECT 586.330 53.290 587.510 54.470 ;
        RECT 587.930 53.290 589.110 54.470 ;
        RECT 586.330 51.690 587.510 52.870 ;
        RECT 587.930 51.690 589.110 52.870 ;
        RECT 586.330 -22.110 587.510 -20.930 ;
        RECT 587.930 -22.110 589.110 -20.930 ;
        RECT 586.330 -23.710 587.510 -22.530 ;
        RECT 587.930 -23.710 589.110 -22.530 ;
        RECT 766.330 233.290 767.510 234.470 ;
        RECT 767.930 233.290 769.110 234.470 ;
        RECT 766.330 231.690 767.510 232.870 ;
        RECT 767.930 231.690 769.110 232.870 ;
        RECT 766.330 53.290 767.510 54.470 ;
        RECT 767.930 53.290 769.110 54.470 ;
        RECT 766.330 51.690 767.510 52.870 ;
        RECT 767.930 51.690 769.110 52.870 ;
        RECT 766.330 -22.110 767.510 -20.930 ;
        RECT 767.930 -22.110 769.110 -20.930 ;
        RECT 766.330 -23.710 767.510 -22.530 ;
        RECT 767.930 -23.710 769.110 -22.530 ;
        RECT 946.330 233.290 947.510 234.470 ;
        RECT 947.930 233.290 949.110 234.470 ;
        RECT 946.330 231.690 947.510 232.870 ;
        RECT 947.930 231.690 949.110 232.870 ;
        RECT 946.330 53.290 947.510 54.470 ;
        RECT 947.930 53.290 949.110 54.470 ;
        RECT 946.330 51.690 947.510 52.870 ;
        RECT 947.930 51.690 949.110 52.870 ;
        RECT 946.330 -22.110 947.510 -20.930 ;
        RECT 947.930 -22.110 949.110 -20.930 ;
        RECT 946.330 -23.710 947.510 -22.530 ;
        RECT 947.930 -23.710 949.110 -22.530 ;
        RECT 1126.330 233.290 1127.510 234.470 ;
        RECT 1127.930 233.290 1129.110 234.470 ;
        RECT 1126.330 231.690 1127.510 232.870 ;
        RECT 1127.930 231.690 1129.110 232.870 ;
        RECT 1126.330 53.290 1127.510 54.470 ;
        RECT 1127.930 53.290 1129.110 54.470 ;
        RECT 1126.330 51.690 1127.510 52.870 ;
        RECT 1127.930 51.690 1129.110 52.870 ;
        RECT 1126.330 -22.110 1127.510 -20.930 ;
        RECT 1127.930 -22.110 1129.110 -20.930 ;
        RECT 1126.330 -23.710 1127.510 -22.530 ;
        RECT 1127.930 -23.710 1129.110 -22.530 ;
        RECT 1306.330 3542.210 1307.510 3543.390 ;
        RECT 1307.930 3542.210 1309.110 3543.390 ;
        RECT 1306.330 3540.610 1307.510 3541.790 ;
        RECT 1307.930 3540.610 1309.110 3541.790 ;
        RECT 1306.330 3473.290 1307.510 3474.470 ;
        RECT 1307.930 3473.290 1309.110 3474.470 ;
        RECT 1306.330 3471.690 1307.510 3472.870 ;
        RECT 1307.930 3471.690 1309.110 3472.870 ;
        RECT 1306.330 3293.290 1307.510 3294.470 ;
        RECT 1307.930 3293.290 1309.110 3294.470 ;
        RECT 1306.330 3291.690 1307.510 3292.870 ;
        RECT 1307.930 3291.690 1309.110 3292.870 ;
        RECT 1306.330 3113.290 1307.510 3114.470 ;
        RECT 1307.930 3113.290 1309.110 3114.470 ;
        RECT 1306.330 3111.690 1307.510 3112.870 ;
        RECT 1307.930 3111.690 1309.110 3112.870 ;
        RECT 1306.330 2933.290 1307.510 2934.470 ;
        RECT 1307.930 2933.290 1309.110 2934.470 ;
        RECT 1306.330 2931.690 1307.510 2932.870 ;
        RECT 1307.930 2931.690 1309.110 2932.870 ;
        RECT 1306.330 2753.290 1307.510 2754.470 ;
        RECT 1307.930 2753.290 1309.110 2754.470 ;
        RECT 1306.330 2751.690 1307.510 2752.870 ;
        RECT 1307.930 2751.690 1309.110 2752.870 ;
        RECT 1306.330 2573.290 1307.510 2574.470 ;
        RECT 1307.930 2573.290 1309.110 2574.470 ;
        RECT 1306.330 2571.690 1307.510 2572.870 ;
        RECT 1307.930 2571.690 1309.110 2572.870 ;
        RECT 1306.330 2393.290 1307.510 2394.470 ;
        RECT 1307.930 2393.290 1309.110 2394.470 ;
        RECT 1306.330 2391.690 1307.510 2392.870 ;
        RECT 1307.930 2391.690 1309.110 2392.870 ;
        RECT 1306.330 2213.290 1307.510 2214.470 ;
        RECT 1307.930 2213.290 1309.110 2214.470 ;
        RECT 1306.330 2211.690 1307.510 2212.870 ;
        RECT 1307.930 2211.690 1309.110 2212.870 ;
        RECT 1306.330 2033.290 1307.510 2034.470 ;
        RECT 1307.930 2033.290 1309.110 2034.470 ;
        RECT 1306.330 2031.690 1307.510 2032.870 ;
        RECT 1307.930 2031.690 1309.110 2032.870 ;
        RECT 1306.330 1853.290 1307.510 1854.470 ;
        RECT 1307.930 1853.290 1309.110 1854.470 ;
        RECT 1306.330 1851.690 1307.510 1852.870 ;
        RECT 1307.930 1851.690 1309.110 1852.870 ;
        RECT 1306.330 1673.290 1307.510 1674.470 ;
        RECT 1307.930 1673.290 1309.110 1674.470 ;
        RECT 1306.330 1671.690 1307.510 1672.870 ;
        RECT 1307.930 1671.690 1309.110 1672.870 ;
        RECT 1306.330 1493.290 1307.510 1494.470 ;
        RECT 1307.930 1493.290 1309.110 1494.470 ;
        RECT 1306.330 1491.690 1307.510 1492.870 ;
        RECT 1307.930 1491.690 1309.110 1492.870 ;
        RECT 1306.330 1313.290 1307.510 1314.470 ;
        RECT 1307.930 1313.290 1309.110 1314.470 ;
        RECT 1306.330 1311.690 1307.510 1312.870 ;
        RECT 1307.930 1311.690 1309.110 1312.870 ;
        RECT 1306.330 1133.290 1307.510 1134.470 ;
        RECT 1307.930 1133.290 1309.110 1134.470 ;
        RECT 1306.330 1131.690 1307.510 1132.870 ;
        RECT 1307.930 1131.690 1309.110 1132.870 ;
        RECT 1306.330 953.290 1307.510 954.470 ;
        RECT 1307.930 953.290 1309.110 954.470 ;
        RECT 1306.330 951.690 1307.510 952.870 ;
        RECT 1307.930 951.690 1309.110 952.870 ;
        RECT 1306.330 773.290 1307.510 774.470 ;
        RECT 1307.930 773.290 1309.110 774.470 ;
        RECT 1306.330 771.690 1307.510 772.870 ;
        RECT 1307.930 771.690 1309.110 772.870 ;
        RECT 1306.330 593.290 1307.510 594.470 ;
        RECT 1307.930 593.290 1309.110 594.470 ;
        RECT 1306.330 591.690 1307.510 592.870 ;
        RECT 1307.930 591.690 1309.110 592.870 ;
        RECT 1306.330 413.290 1307.510 414.470 ;
        RECT 1307.930 413.290 1309.110 414.470 ;
        RECT 1306.330 411.690 1307.510 412.870 ;
        RECT 1307.930 411.690 1309.110 412.870 ;
        RECT 1306.330 233.290 1307.510 234.470 ;
        RECT 1307.930 233.290 1309.110 234.470 ;
        RECT 1306.330 231.690 1307.510 232.870 ;
        RECT 1307.930 231.690 1309.110 232.870 ;
        RECT 1306.330 53.290 1307.510 54.470 ;
        RECT 1307.930 53.290 1309.110 54.470 ;
        RECT 1306.330 51.690 1307.510 52.870 ;
        RECT 1307.930 51.690 1309.110 52.870 ;
        RECT 1306.330 -22.110 1307.510 -20.930 ;
        RECT 1307.930 -22.110 1309.110 -20.930 ;
        RECT 1306.330 -23.710 1307.510 -22.530 ;
        RECT 1307.930 -23.710 1309.110 -22.530 ;
        RECT 1486.330 3542.210 1487.510 3543.390 ;
        RECT 1487.930 3542.210 1489.110 3543.390 ;
        RECT 1486.330 3540.610 1487.510 3541.790 ;
        RECT 1487.930 3540.610 1489.110 3541.790 ;
        RECT 1486.330 3473.290 1487.510 3474.470 ;
        RECT 1487.930 3473.290 1489.110 3474.470 ;
        RECT 1486.330 3471.690 1487.510 3472.870 ;
        RECT 1487.930 3471.690 1489.110 3472.870 ;
        RECT 1486.330 3293.290 1487.510 3294.470 ;
        RECT 1487.930 3293.290 1489.110 3294.470 ;
        RECT 1486.330 3291.690 1487.510 3292.870 ;
        RECT 1487.930 3291.690 1489.110 3292.870 ;
        RECT 1486.330 3113.290 1487.510 3114.470 ;
        RECT 1487.930 3113.290 1489.110 3114.470 ;
        RECT 1486.330 3111.690 1487.510 3112.870 ;
        RECT 1487.930 3111.690 1489.110 3112.870 ;
        RECT 1486.330 2933.290 1487.510 2934.470 ;
        RECT 1487.930 2933.290 1489.110 2934.470 ;
        RECT 1486.330 2931.690 1487.510 2932.870 ;
        RECT 1487.930 2931.690 1489.110 2932.870 ;
        RECT 1486.330 2753.290 1487.510 2754.470 ;
        RECT 1487.930 2753.290 1489.110 2754.470 ;
        RECT 1486.330 2751.690 1487.510 2752.870 ;
        RECT 1487.930 2751.690 1489.110 2752.870 ;
        RECT 1486.330 2573.290 1487.510 2574.470 ;
        RECT 1487.930 2573.290 1489.110 2574.470 ;
        RECT 1486.330 2571.690 1487.510 2572.870 ;
        RECT 1487.930 2571.690 1489.110 2572.870 ;
        RECT 1486.330 2393.290 1487.510 2394.470 ;
        RECT 1487.930 2393.290 1489.110 2394.470 ;
        RECT 1486.330 2391.690 1487.510 2392.870 ;
        RECT 1487.930 2391.690 1489.110 2392.870 ;
        RECT 1486.330 2213.290 1487.510 2214.470 ;
        RECT 1487.930 2213.290 1489.110 2214.470 ;
        RECT 1486.330 2211.690 1487.510 2212.870 ;
        RECT 1487.930 2211.690 1489.110 2212.870 ;
        RECT 1486.330 2033.290 1487.510 2034.470 ;
        RECT 1487.930 2033.290 1489.110 2034.470 ;
        RECT 1486.330 2031.690 1487.510 2032.870 ;
        RECT 1487.930 2031.690 1489.110 2032.870 ;
        RECT 1486.330 1853.290 1487.510 1854.470 ;
        RECT 1487.930 1853.290 1489.110 1854.470 ;
        RECT 1486.330 1851.690 1487.510 1852.870 ;
        RECT 1487.930 1851.690 1489.110 1852.870 ;
        RECT 1486.330 1673.290 1487.510 1674.470 ;
        RECT 1487.930 1673.290 1489.110 1674.470 ;
        RECT 1486.330 1671.690 1487.510 1672.870 ;
        RECT 1487.930 1671.690 1489.110 1672.870 ;
        RECT 1486.330 1493.290 1487.510 1494.470 ;
        RECT 1487.930 1493.290 1489.110 1494.470 ;
        RECT 1486.330 1491.690 1487.510 1492.870 ;
        RECT 1487.930 1491.690 1489.110 1492.870 ;
        RECT 1486.330 1313.290 1487.510 1314.470 ;
        RECT 1487.930 1313.290 1489.110 1314.470 ;
        RECT 1486.330 1311.690 1487.510 1312.870 ;
        RECT 1487.930 1311.690 1489.110 1312.870 ;
        RECT 1486.330 1133.290 1487.510 1134.470 ;
        RECT 1487.930 1133.290 1489.110 1134.470 ;
        RECT 1486.330 1131.690 1487.510 1132.870 ;
        RECT 1487.930 1131.690 1489.110 1132.870 ;
        RECT 1486.330 953.290 1487.510 954.470 ;
        RECT 1487.930 953.290 1489.110 954.470 ;
        RECT 1486.330 951.690 1487.510 952.870 ;
        RECT 1487.930 951.690 1489.110 952.870 ;
        RECT 1486.330 773.290 1487.510 774.470 ;
        RECT 1487.930 773.290 1489.110 774.470 ;
        RECT 1486.330 771.690 1487.510 772.870 ;
        RECT 1487.930 771.690 1489.110 772.870 ;
        RECT 1486.330 593.290 1487.510 594.470 ;
        RECT 1487.930 593.290 1489.110 594.470 ;
        RECT 1486.330 591.690 1487.510 592.870 ;
        RECT 1487.930 591.690 1489.110 592.870 ;
        RECT 1486.330 413.290 1487.510 414.470 ;
        RECT 1487.930 413.290 1489.110 414.470 ;
        RECT 1486.330 411.690 1487.510 412.870 ;
        RECT 1487.930 411.690 1489.110 412.870 ;
        RECT 1486.330 233.290 1487.510 234.470 ;
        RECT 1487.930 233.290 1489.110 234.470 ;
        RECT 1486.330 231.690 1487.510 232.870 ;
        RECT 1487.930 231.690 1489.110 232.870 ;
        RECT 1486.330 53.290 1487.510 54.470 ;
        RECT 1487.930 53.290 1489.110 54.470 ;
        RECT 1486.330 51.690 1487.510 52.870 ;
        RECT 1487.930 51.690 1489.110 52.870 ;
        RECT 1486.330 -22.110 1487.510 -20.930 ;
        RECT 1487.930 -22.110 1489.110 -20.930 ;
        RECT 1486.330 -23.710 1487.510 -22.530 ;
        RECT 1487.930 -23.710 1489.110 -22.530 ;
        RECT 1666.330 3542.210 1667.510 3543.390 ;
        RECT 1667.930 3542.210 1669.110 3543.390 ;
        RECT 1666.330 3540.610 1667.510 3541.790 ;
        RECT 1667.930 3540.610 1669.110 3541.790 ;
        RECT 1666.330 3473.290 1667.510 3474.470 ;
        RECT 1667.930 3473.290 1669.110 3474.470 ;
        RECT 1666.330 3471.690 1667.510 3472.870 ;
        RECT 1667.930 3471.690 1669.110 3472.870 ;
        RECT 1666.330 3293.290 1667.510 3294.470 ;
        RECT 1667.930 3293.290 1669.110 3294.470 ;
        RECT 1666.330 3291.690 1667.510 3292.870 ;
        RECT 1667.930 3291.690 1669.110 3292.870 ;
        RECT 1666.330 3113.290 1667.510 3114.470 ;
        RECT 1667.930 3113.290 1669.110 3114.470 ;
        RECT 1666.330 3111.690 1667.510 3112.870 ;
        RECT 1667.930 3111.690 1669.110 3112.870 ;
        RECT 1666.330 2933.290 1667.510 2934.470 ;
        RECT 1667.930 2933.290 1669.110 2934.470 ;
        RECT 1666.330 2931.690 1667.510 2932.870 ;
        RECT 1667.930 2931.690 1669.110 2932.870 ;
        RECT 1666.330 2753.290 1667.510 2754.470 ;
        RECT 1667.930 2753.290 1669.110 2754.470 ;
        RECT 1666.330 2751.690 1667.510 2752.870 ;
        RECT 1667.930 2751.690 1669.110 2752.870 ;
        RECT 1666.330 2573.290 1667.510 2574.470 ;
        RECT 1667.930 2573.290 1669.110 2574.470 ;
        RECT 1666.330 2571.690 1667.510 2572.870 ;
        RECT 1667.930 2571.690 1669.110 2572.870 ;
        RECT 1666.330 2393.290 1667.510 2394.470 ;
        RECT 1667.930 2393.290 1669.110 2394.470 ;
        RECT 1666.330 2391.690 1667.510 2392.870 ;
        RECT 1667.930 2391.690 1669.110 2392.870 ;
        RECT 1666.330 2213.290 1667.510 2214.470 ;
        RECT 1667.930 2213.290 1669.110 2214.470 ;
        RECT 1666.330 2211.690 1667.510 2212.870 ;
        RECT 1667.930 2211.690 1669.110 2212.870 ;
        RECT 1666.330 2033.290 1667.510 2034.470 ;
        RECT 1667.930 2033.290 1669.110 2034.470 ;
        RECT 1666.330 2031.690 1667.510 2032.870 ;
        RECT 1667.930 2031.690 1669.110 2032.870 ;
        RECT 1666.330 1853.290 1667.510 1854.470 ;
        RECT 1667.930 1853.290 1669.110 1854.470 ;
        RECT 1666.330 1851.690 1667.510 1852.870 ;
        RECT 1667.930 1851.690 1669.110 1852.870 ;
        RECT 1666.330 1673.290 1667.510 1674.470 ;
        RECT 1667.930 1673.290 1669.110 1674.470 ;
        RECT 1666.330 1671.690 1667.510 1672.870 ;
        RECT 1667.930 1671.690 1669.110 1672.870 ;
        RECT 1666.330 1493.290 1667.510 1494.470 ;
        RECT 1667.930 1493.290 1669.110 1494.470 ;
        RECT 1666.330 1491.690 1667.510 1492.870 ;
        RECT 1667.930 1491.690 1669.110 1492.870 ;
        RECT 1666.330 1313.290 1667.510 1314.470 ;
        RECT 1667.930 1313.290 1669.110 1314.470 ;
        RECT 1666.330 1311.690 1667.510 1312.870 ;
        RECT 1667.930 1311.690 1669.110 1312.870 ;
        RECT 1666.330 1133.290 1667.510 1134.470 ;
        RECT 1667.930 1133.290 1669.110 1134.470 ;
        RECT 1666.330 1131.690 1667.510 1132.870 ;
        RECT 1667.930 1131.690 1669.110 1132.870 ;
        RECT 1666.330 953.290 1667.510 954.470 ;
        RECT 1667.930 953.290 1669.110 954.470 ;
        RECT 1666.330 951.690 1667.510 952.870 ;
        RECT 1667.930 951.690 1669.110 952.870 ;
        RECT 1666.330 773.290 1667.510 774.470 ;
        RECT 1667.930 773.290 1669.110 774.470 ;
        RECT 1666.330 771.690 1667.510 772.870 ;
        RECT 1667.930 771.690 1669.110 772.870 ;
        RECT 1666.330 593.290 1667.510 594.470 ;
        RECT 1667.930 593.290 1669.110 594.470 ;
        RECT 1666.330 591.690 1667.510 592.870 ;
        RECT 1667.930 591.690 1669.110 592.870 ;
        RECT 1666.330 413.290 1667.510 414.470 ;
        RECT 1667.930 413.290 1669.110 414.470 ;
        RECT 1666.330 411.690 1667.510 412.870 ;
        RECT 1667.930 411.690 1669.110 412.870 ;
        RECT 1666.330 233.290 1667.510 234.470 ;
        RECT 1667.930 233.290 1669.110 234.470 ;
        RECT 1666.330 231.690 1667.510 232.870 ;
        RECT 1667.930 231.690 1669.110 232.870 ;
        RECT 1666.330 53.290 1667.510 54.470 ;
        RECT 1667.930 53.290 1669.110 54.470 ;
        RECT 1666.330 51.690 1667.510 52.870 ;
        RECT 1667.930 51.690 1669.110 52.870 ;
        RECT 1666.330 -22.110 1667.510 -20.930 ;
        RECT 1667.930 -22.110 1669.110 -20.930 ;
        RECT 1666.330 -23.710 1667.510 -22.530 ;
        RECT 1667.930 -23.710 1669.110 -22.530 ;
        RECT 1846.330 3542.210 1847.510 3543.390 ;
        RECT 1847.930 3542.210 1849.110 3543.390 ;
        RECT 1846.330 3540.610 1847.510 3541.790 ;
        RECT 1847.930 3540.610 1849.110 3541.790 ;
        RECT 1846.330 3473.290 1847.510 3474.470 ;
        RECT 1847.930 3473.290 1849.110 3474.470 ;
        RECT 1846.330 3471.690 1847.510 3472.870 ;
        RECT 1847.930 3471.690 1849.110 3472.870 ;
        RECT 1846.330 3293.290 1847.510 3294.470 ;
        RECT 1847.930 3293.290 1849.110 3294.470 ;
        RECT 1846.330 3291.690 1847.510 3292.870 ;
        RECT 1847.930 3291.690 1849.110 3292.870 ;
        RECT 1846.330 3113.290 1847.510 3114.470 ;
        RECT 1847.930 3113.290 1849.110 3114.470 ;
        RECT 1846.330 3111.690 1847.510 3112.870 ;
        RECT 1847.930 3111.690 1849.110 3112.870 ;
        RECT 1846.330 2933.290 1847.510 2934.470 ;
        RECT 1847.930 2933.290 1849.110 2934.470 ;
        RECT 1846.330 2931.690 1847.510 2932.870 ;
        RECT 1847.930 2931.690 1849.110 2932.870 ;
        RECT 1846.330 2753.290 1847.510 2754.470 ;
        RECT 1847.930 2753.290 1849.110 2754.470 ;
        RECT 1846.330 2751.690 1847.510 2752.870 ;
        RECT 1847.930 2751.690 1849.110 2752.870 ;
        RECT 1846.330 2573.290 1847.510 2574.470 ;
        RECT 1847.930 2573.290 1849.110 2574.470 ;
        RECT 1846.330 2571.690 1847.510 2572.870 ;
        RECT 1847.930 2571.690 1849.110 2572.870 ;
        RECT 1846.330 2393.290 1847.510 2394.470 ;
        RECT 1847.930 2393.290 1849.110 2394.470 ;
        RECT 1846.330 2391.690 1847.510 2392.870 ;
        RECT 1847.930 2391.690 1849.110 2392.870 ;
        RECT 1846.330 2213.290 1847.510 2214.470 ;
        RECT 1847.930 2213.290 1849.110 2214.470 ;
        RECT 1846.330 2211.690 1847.510 2212.870 ;
        RECT 1847.930 2211.690 1849.110 2212.870 ;
        RECT 1846.330 2033.290 1847.510 2034.470 ;
        RECT 1847.930 2033.290 1849.110 2034.470 ;
        RECT 1846.330 2031.690 1847.510 2032.870 ;
        RECT 1847.930 2031.690 1849.110 2032.870 ;
        RECT 1846.330 1853.290 1847.510 1854.470 ;
        RECT 1847.930 1853.290 1849.110 1854.470 ;
        RECT 1846.330 1851.690 1847.510 1852.870 ;
        RECT 1847.930 1851.690 1849.110 1852.870 ;
        RECT 1846.330 1673.290 1847.510 1674.470 ;
        RECT 1847.930 1673.290 1849.110 1674.470 ;
        RECT 1846.330 1671.690 1847.510 1672.870 ;
        RECT 1847.930 1671.690 1849.110 1672.870 ;
        RECT 1846.330 1493.290 1847.510 1494.470 ;
        RECT 1847.930 1493.290 1849.110 1494.470 ;
        RECT 1846.330 1491.690 1847.510 1492.870 ;
        RECT 1847.930 1491.690 1849.110 1492.870 ;
        RECT 1846.330 1313.290 1847.510 1314.470 ;
        RECT 1847.930 1313.290 1849.110 1314.470 ;
        RECT 1846.330 1311.690 1847.510 1312.870 ;
        RECT 1847.930 1311.690 1849.110 1312.870 ;
        RECT 1846.330 1133.290 1847.510 1134.470 ;
        RECT 1847.930 1133.290 1849.110 1134.470 ;
        RECT 1846.330 1131.690 1847.510 1132.870 ;
        RECT 1847.930 1131.690 1849.110 1132.870 ;
        RECT 1846.330 953.290 1847.510 954.470 ;
        RECT 1847.930 953.290 1849.110 954.470 ;
        RECT 1846.330 951.690 1847.510 952.870 ;
        RECT 1847.930 951.690 1849.110 952.870 ;
        RECT 1846.330 773.290 1847.510 774.470 ;
        RECT 1847.930 773.290 1849.110 774.470 ;
        RECT 1846.330 771.690 1847.510 772.870 ;
        RECT 1847.930 771.690 1849.110 772.870 ;
        RECT 1846.330 593.290 1847.510 594.470 ;
        RECT 1847.930 593.290 1849.110 594.470 ;
        RECT 1846.330 591.690 1847.510 592.870 ;
        RECT 1847.930 591.690 1849.110 592.870 ;
        RECT 1846.330 413.290 1847.510 414.470 ;
        RECT 1847.930 413.290 1849.110 414.470 ;
        RECT 1846.330 411.690 1847.510 412.870 ;
        RECT 1847.930 411.690 1849.110 412.870 ;
        RECT 1846.330 233.290 1847.510 234.470 ;
        RECT 1847.930 233.290 1849.110 234.470 ;
        RECT 1846.330 231.690 1847.510 232.870 ;
        RECT 1847.930 231.690 1849.110 232.870 ;
        RECT 1846.330 53.290 1847.510 54.470 ;
        RECT 1847.930 53.290 1849.110 54.470 ;
        RECT 1846.330 51.690 1847.510 52.870 ;
        RECT 1847.930 51.690 1849.110 52.870 ;
        RECT 1846.330 -22.110 1847.510 -20.930 ;
        RECT 1847.930 -22.110 1849.110 -20.930 ;
        RECT 1846.330 -23.710 1847.510 -22.530 ;
        RECT 1847.930 -23.710 1849.110 -22.530 ;
        RECT 2026.330 3542.210 2027.510 3543.390 ;
        RECT 2027.930 3542.210 2029.110 3543.390 ;
        RECT 2026.330 3540.610 2027.510 3541.790 ;
        RECT 2027.930 3540.610 2029.110 3541.790 ;
        RECT 2026.330 3473.290 2027.510 3474.470 ;
        RECT 2027.930 3473.290 2029.110 3474.470 ;
        RECT 2026.330 3471.690 2027.510 3472.870 ;
        RECT 2027.930 3471.690 2029.110 3472.870 ;
        RECT 2026.330 3293.290 2027.510 3294.470 ;
        RECT 2027.930 3293.290 2029.110 3294.470 ;
        RECT 2026.330 3291.690 2027.510 3292.870 ;
        RECT 2027.930 3291.690 2029.110 3292.870 ;
        RECT 2026.330 3113.290 2027.510 3114.470 ;
        RECT 2027.930 3113.290 2029.110 3114.470 ;
        RECT 2026.330 3111.690 2027.510 3112.870 ;
        RECT 2027.930 3111.690 2029.110 3112.870 ;
        RECT 2026.330 2933.290 2027.510 2934.470 ;
        RECT 2027.930 2933.290 2029.110 2934.470 ;
        RECT 2026.330 2931.690 2027.510 2932.870 ;
        RECT 2027.930 2931.690 2029.110 2932.870 ;
        RECT 2026.330 2753.290 2027.510 2754.470 ;
        RECT 2027.930 2753.290 2029.110 2754.470 ;
        RECT 2026.330 2751.690 2027.510 2752.870 ;
        RECT 2027.930 2751.690 2029.110 2752.870 ;
        RECT 2026.330 2573.290 2027.510 2574.470 ;
        RECT 2027.930 2573.290 2029.110 2574.470 ;
        RECT 2026.330 2571.690 2027.510 2572.870 ;
        RECT 2027.930 2571.690 2029.110 2572.870 ;
        RECT 2026.330 2393.290 2027.510 2394.470 ;
        RECT 2027.930 2393.290 2029.110 2394.470 ;
        RECT 2026.330 2391.690 2027.510 2392.870 ;
        RECT 2027.930 2391.690 2029.110 2392.870 ;
        RECT 2026.330 2213.290 2027.510 2214.470 ;
        RECT 2027.930 2213.290 2029.110 2214.470 ;
        RECT 2026.330 2211.690 2027.510 2212.870 ;
        RECT 2027.930 2211.690 2029.110 2212.870 ;
        RECT 2026.330 2033.290 2027.510 2034.470 ;
        RECT 2027.930 2033.290 2029.110 2034.470 ;
        RECT 2026.330 2031.690 2027.510 2032.870 ;
        RECT 2027.930 2031.690 2029.110 2032.870 ;
        RECT 2026.330 1853.290 2027.510 1854.470 ;
        RECT 2027.930 1853.290 2029.110 1854.470 ;
        RECT 2026.330 1851.690 2027.510 1852.870 ;
        RECT 2027.930 1851.690 2029.110 1852.870 ;
        RECT 2026.330 1673.290 2027.510 1674.470 ;
        RECT 2027.930 1673.290 2029.110 1674.470 ;
        RECT 2026.330 1671.690 2027.510 1672.870 ;
        RECT 2027.930 1671.690 2029.110 1672.870 ;
        RECT 2026.330 1493.290 2027.510 1494.470 ;
        RECT 2027.930 1493.290 2029.110 1494.470 ;
        RECT 2026.330 1491.690 2027.510 1492.870 ;
        RECT 2027.930 1491.690 2029.110 1492.870 ;
        RECT 2026.330 1313.290 2027.510 1314.470 ;
        RECT 2027.930 1313.290 2029.110 1314.470 ;
        RECT 2026.330 1311.690 2027.510 1312.870 ;
        RECT 2027.930 1311.690 2029.110 1312.870 ;
        RECT 2026.330 1133.290 2027.510 1134.470 ;
        RECT 2027.930 1133.290 2029.110 1134.470 ;
        RECT 2026.330 1131.690 2027.510 1132.870 ;
        RECT 2027.930 1131.690 2029.110 1132.870 ;
        RECT 2026.330 953.290 2027.510 954.470 ;
        RECT 2027.930 953.290 2029.110 954.470 ;
        RECT 2026.330 951.690 2027.510 952.870 ;
        RECT 2027.930 951.690 2029.110 952.870 ;
        RECT 2026.330 773.290 2027.510 774.470 ;
        RECT 2027.930 773.290 2029.110 774.470 ;
        RECT 2026.330 771.690 2027.510 772.870 ;
        RECT 2027.930 771.690 2029.110 772.870 ;
        RECT 2026.330 593.290 2027.510 594.470 ;
        RECT 2027.930 593.290 2029.110 594.470 ;
        RECT 2026.330 591.690 2027.510 592.870 ;
        RECT 2027.930 591.690 2029.110 592.870 ;
        RECT 2026.330 413.290 2027.510 414.470 ;
        RECT 2027.930 413.290 2029.110 414.470 ;
        RECT 2026.330 411.690 2027.510 412.870 ;
        RECT 2027.930 411.690 2029.110 412.870 ;
        RECT 2026.330 233.290 2027.510 234.470 ;
        RECT 2027.930 233.290 2029.110 234.470 ;
        RECT 2026.330 231.690 2027.510 232.870 ;
        RECT 2027.930 231.690 2029.110 232.870 ;
        RECT 2026.330 53.290 2027.510 54.470 ;
        RECT 2027.930 53.290 2029.110 54.470 ;
        RECT 2026.330 51.690 2027.510 52.870 ;
        RECT 2027.930 51.690 2029.110 52.870 ;
        RECT 2026.330 -22.110 2027.510 -20.930 ;
        RECT 2027.930 -22.110 2029.110 -20.930 ;
        RECT 2026.330 -23.710 2027.510 -22.530 ;
        RECT 2027.930 -23.710 2029.110 -22.530 ;
        RECT 2206.330 3542.210 2207.510 3543.390 ;
        RECT 2207.930 3542.210 2209.110 3543.390 ;
        RECT 2206.330 3540.610 2207.510 3541.790 ;
        RECT 2207.930 3540.610 2209.110 3541.790 ;
        RECT 2206.330 3473.290 2207.510 3474.470 ;
        RECT 2207.930 3473.290 2209.110 3474.470 ;
        RECT 2206.330 3471.690 2207.510 3472.870 ;
        RECT 2207.930 3471.690 2209.110 3472.870 ;
        RECT 2206.330 3293.290 2207.510 3294.470 ;
        RECT 2207.930 3293.290 2209.110 3294.470 ;
        RECT 2206.330 3291.690 2207.510 3292.870 ;
        RECT 2207.930 3291.690 2209.110 3292.870 ;
        RECT 2206.330 3113.290 2207.510 3114.470 ;
        RECT 2207.930 3113.290 2209.110 3114.470 ;
        RECT 2206.330 3111.690 2207.510 3112.870 ;
        RECT 2207.930 3111.690 2209.110 3112.870 ;
        RECT 2206.330 2933.290 2207.510 2934.470 ;
        RECT 2207.930 2933.290 2209.110 2934.470 ;
        RECT 2206.330 2931.690 2207.510 2932.870 ;
        RECT 2207.930 2931.690 2209.110 2932.870 ;
        RECT 2206.330 2753.290 2207.510 2754.470 ;
        RECT 2207.930 2753.290 2209.110 2754.470 ;
        RECT 2206.330 2751.690 2207.510 2752.870 ;
        RECT 2207.930 2751.690 2209.110 2752.870 ;
        RECT 2206.330 2573.290 2207.510 2574.470 ;
        RECT 2207.930 2573.290 2209.110 2574.470 ;
        RECT 2206.330 2571.690 2207.510 2572.870 ;
        RECT 2207.930 2571.690 2209.110 2572.870 ;
        RECT 2206.330 2393.290 2207.510 2394.470 ;
        RECT 2207.930 2393.290 2209.110 2394.470 ;
        RECT 2206.330 2391.690 2207.510 2392.870 ;
        RECT 2207.930 2391.690 2209.110 2392.870 ;
        RECT 2206.330 2213.290 2207.510 2214.470 ;
        RECT 2207.930 2213.290 2209.110 2214.470 ;
        RECT 2206.330 2211.690 2207.510 2212.870 ;
        RECT 2207.930 2211.690 2209.110 2212.870 ;
        RECT 2206.330 2033.290 2207.510 2034.470 ;
        RECT 2207.930 2033.290 2209.110 2034.470 ;
        RECT 2206.330 2031.690 2207.510 2032.870 ;
        RECT 2207.930 2031.690 2209.110 2032.870 ;
        RECT 2206.330 1853.290 2207.510 1854.470 ;
        RECT 2207.930 1853.290 2209.110 1854.470 ;
        RECT 2206.330 1851.690 2207.510 1852.870 ;
        RECT 2207.930 1851.690 2209.110 1852.870 ;
        RECT 2206.330 1673.290 2207.510 1674.470 ;
        RECT 2207.930 1673.290 2209.110 1674.470 ;
        RECT 2206.330 1671.690 2207.510 1672.870 ;
        RECT 2207.930 1671.690 2209.110 1672.870 ;
        RECT 2206.330 1493.290 2207.510 1494.470 ;
        RECT 2207.930 1493.290 2209.110 1494.470 ;
        RECT 2206.330 1491.690 2207.510 1492.870 ;
        RECT 2207.930 1491.690 2209.110 1492.870 ;
        RECT 2206.330 1313.290 2207.510 1314.470 ;
        RECT 2207.930 1313.290 2209.110 1314.470 ;
        RECT 2206.330 1311.690 2207.510 1312.870 ;
        RECT 2207.930 1311.690 2209.110 1312.870 ;
        RECT 2206.330 1133.290 2207.510 1134.470 ;
        RECT 2207.930 1133.290 2209.110 1134.470 ;
        RECT 2206.330 1131.690 2207.510 1132.870 ;
        RECT 2207.930 1131.690 2209.110 1132.870 ;
        RECT 2206.330 953.290 2207.510 954.470 ;
        RECT 2207.930 953.290 2209.110 954.470 ;
        RECT 2206.330 951.690 2207.510 952.870 ;
        RECT 2207.930 951.690 2209.110 952.870 ;
        RECT 2206.330 773.290 2207.510 774.470 ;
        RECT 2207.930 773.290 2209.110 774.470 ;
        RECT 2206.330 771.690 2207.510 772.870 ;
        RECT 2207.930 771.690 2209.110 772.870 ;
        RECT 2206.330 593.290 2207.510 594.470 ;
        RECT 2207.930 593.290 2209.110 594.470 ;
        RECT 2206.330 591.690 2207.510 592.870 ;
        RECT 2207.930 591.690 2209.110 592.870 ;
        RECT 2206.330 413.290 2207.510 414.470 ;
        RECT 2207.930 413.290 2209.110 414.470 ;
        RECT 2206.330 411.690 2207.510 412.870 ;
        RECT 2207.930 411.690 2209.110 412.870 ;
        RECT 2206.330 233.290 2207.510 234.470 ;
        RECT 2207.930 233.290 2209.110 234.470 ;
        RECT 2206.330 231.690 2207.510 232.870 ;
        RECT 2207.930 231.690 2209.110 232.870 ;
        RECT 2206.330 53.290 2207.510 54.470 ;
        RECT 2207.930 53.290 2209.110 54.470 ;
        RECT 2206.330 51.690 2207.510 52.870 ;
        RECT 2207.930 51.690 2209.110 52.870 ;
        RECT 2206.330 -22.110 2207.510 -20.930 ;
        RECT 2207.930 -22.110 2209.110 -20.930 ;
        RECT 2206.330 -23.710 2207.510 -22.530 ;
        RECT 2207.930 -23.710 2209.110 -22.530 ;
        RECT 2386.330 3542.210 2387.510 3543.390 ;
        RECT 2387.930 3542.210 2389.110 3543.390 ;
        RECT 2386.330 3540.610 2387.510 3541.790 ;
        RECT 2387.930 3540.610 2389.110 3541.790 ;
        RECT 2386.330 3473.290 2387.510 3474.470 ;
        RECT 2387.930 3473.290 2389.110 3474.470 ;
        RECT 2386.330 3471.690 2387.510 3472.870 ;
        RECT 2387.930 3471.690 2389.110 3472.870 ;
        RECT 2386.330 3293.290 2387.510 3294.470 ;
        RECT 2387.930 3293.290 2389.110 3294.470 ;
        RECT 2386.330 3291.690 2387.510 3292.870 ;
        RECT 2387.930 3291.690 2389.110 3292.870 ;
        RECT 2386.330 3113.290 2387.510 3114.470 ;
        RECT 2387.930 3113.290 2389.110 3114.470 ;
        RECT 2386.330 3111.690 2387.510 3112.870 ;
        RECT 2387.930 3111.690 2389.110 3112.870 ;
        RECT 2386.330 2933.290 2387.510 2934.470 ;
        RECT 2387.930 2933.290 2389.110 2934.470 ;
        RECT 2386.330 2931.690 2387.510 2932.870 ;
        RECT 2387.930 2931.690 2389.110 2932.870 ;
        RECT 2386.330 2753.290 2387.510 2754.470 ;
        RECT 2387.930 2753.290 2389.110 2754.470 ;
        RECT 2386.330 2751.690 2387.510 2752.870 ;
        RECT 2387.930 2751.690 2389.110 2752.870 ;
        RECT 2386.330 2573.290 2387.510 2574.470 ;
        RECT 2387.930 2573.290 2389.110 2574.470 ;
        RECT 2386.330 2571.690 2387.510 2572.870 ;
        RECT 2387.930 2571.690 2389.110 2572.870 ;
        RECT 2386.330 2393.290 2387.510 2394.470 ;
        RECT 2387.930 2393.290 2389.110 2394.470 ;
        RECT 2386.330 2391.690 2387.510 2392.870 ;
        RECT 2387.930 2391.690 2389.110 2392.870 ;
        RECT 2386.330 2213.290 2387.510 2214.470 ;
        RECT 2387.930 2213.290 2389.110 2214.470 ;
        RECT 2386.330 2211.690 2387.510 2212.870 ;
        RECT 2387.930 2211.690 2389.110 2212.870 ;
        RECT 2386.330 2033.290 2387.510 2034.470 ;
        RECT 2387.930 2033.290 2389.110 2034.470 ;
        RECT 2386.330 2031.690 2387.510 2032.870 ;
        RECT 2387.930 2031.690 2389.110 2032.870 ;
        RECT 2386.330 1853.290 2387.510 1854.470 ;
        RECT 2387.930 1853.290 2389.110 1854.470 ;
        RECT 2386.330 1851.690 2387.510 1852.870 ;
        RECT 2387.930 1851.690 2389.110 1852.870 ;
        RECT 2386.330 1673.290 2387.510 1674.470 ;
        RECT 2387.930 1673.290 2389.110 1674.470 ;
        RECT 2386.330 1671.690 2387.510 1672.870 ;
        RECT 2387.930 1671.690 2389.110 1672.870 ;
        RECT 2386.330 1493.290 2387.510 1494.470 ;
        RECT 2387.930 1493.290 2389.110 1494.470 ;
        RECT 2386.330 1491.690 2387.510 1492.870 ;
        RECT 2387.930 1491.690 2389.110 1492.870 ;
        RECT 2386.330 1313.290 2387.510 1314.470 ;
        RECT 2387.930 1313.290 2389.110 1314.470 ;
        RECT 2386.330 1311.690 2387.510 1312.870 ;
        RECT 2387.930 1311.690 2389.110 1312.870 ;
        RECT 2386.330 1133.290 2387.510 1134.470 ;
        RECT 2387.930 1133.290 2389.110 1134.470 ;
        RECT 2386.330 1131.690 2387.510 1132.870 ;
        RECT 2387.930 1131.690 2389.110 1132.870 ;
        RECT 2386.330 953.290 2387.510 954.470 ;
        RECT 2387.930 953.290 2389.110 954.470 ;
        RECT 2386.330 951.690 2387.510 952.870 ;
        RECT 2387.930 951.690 2389.110 952.870 ;
        RECT 2386.330 773.290 2387.510 774.470 ;
        RECT 2387.930 773.290 2389.110 774.470 ;
        RECT 2386.330 771.690 2387.510 772.870 ;
        RECT 2387.930 771.690 2389.110 772.870 ;
        RECT 2386.330 593.290 2387.510 594.470 ;
        RECT 2387.930 593.290 2389.110 594.470 ;
        RECT 2386.330 591.690 2387.510 592.870 ;
        RECT 2387.930 591.690 2389.110 592.870 ;
        RECT 2386.330 413.290 2387.510 414.470 ;
        RECT 2387.930 413.290 2389.110 414.470 ;
        RECT 2386.330 411.690 2387.510 412.870 ;
        RECT 2387.930 411.690 2389.110 412.870 ;
        RECT 2386.330 233.290 2387.510 234.470 ;
        RECT 2387.930 233.290 2389.110 234.470 ;
        RECT 2386.330 231.690 2387.510 232.870 ;
        RECT 2387.930 231.690 2389.110 232.870 ;
        RECT 2386.330 53.290 2387.510 54.470 ;
        RECT 2387.930 53.290 2389.110 54.470 ;
        RECT 2386.330 51.690 2387.510 52.870 ;
        RECT 2387.930 51.690 2389.110 52.870 ;
        RECT 2386.330 -22.110 2387.510 -20.930 ;
        RECT 2387.930 -22.110 2389.110 -20.930 ;
        RECT 2386.330 -23.710 2387.510 -22.530 ;
        RECT 2387.930 -23.710 2389.110 -22.530 ;
        RECT 2566.330 3542.210 2567.510 3543.390 ;
        RECT 2567.930 3542.210 2569.110 3543.390 ;
        RECT 2566.330 3540.610 2567.510 3541.790 ;
        RECT 2567.930 3540.610 2569.110 3541.790 ;
        RECT 2566.330 3473.290 2567.510 3474.470 ;
        RECT 2567.930 3473.290 2569.110 3474.470 ;
        RECT 2566.330 3471.690 2567.510 3472.870 ;
        RECT 2567.930 3471.690 2569.110 3472.870 ;
        RECT 2566.330 3293.290 2567.510 3294.470 ;
        RECT 2567.930 3293.290 2569.110 3294.470 ;
        RECT 2566.330 3291.690 2567.510 3292.870 ;
        RECT 2567.930 3291.690 2569.110 3292.870 ;
        RECT 2566.330 3113.290 2567.510 3114.470 ;
        RECT 2567.930 3113.290 2569.110 3114.470 ;
        RECT 2566.330 3111.690 2567.510 3112.870 ;
        RECT 2567.930 3111.690 2569.110 3112.870 ;
        RECT 2566.330 2933.290 2567.510 2934.470 ;
        RECT 2567.930 2933.290 2569.110 2934.470 ;
        RECT 2566.330 2931.690 2567.510 2932.870 ;
        RECT 2567.930 2931.690 2569.110 2932.870 ;
        RECT 2566.330 2753.290 2567.510 2754.470 ;
        RECT 2567.930 2753.290 2569.110 2754.470 ;
        RECT 2566.330 2751.690 2567.510 2752.870 ;
        RECT 2567.930 2751.690 2569.110 2752.870 ;
        RECT 2566.330 2573.290 2567.510 2574.470 ;
        RECT 2567.930 2573.290 2569.110 2574.470 ;
        RECT 2566.330 2571.690 2567.510 2572.870 ;
        RECT 2567.930 2571.690 2569.110 2572.870 ;
        RECT 2566.330 2393.290 2567.510 2394.470 ;
        RECT 2567.930 2393.290 2569.110 2394.470 ;
        RECT 2566.330 2391.690 2567.510 2392.870 ;
        RECT 2567.930 2391.690 2569.110 2392.870 ;
        RECT 2566.330 2213.290 2567.510 2214.470 ;
        RECT 2567.930 2213.290 2569.110 2214.470 ;
        RECT 2566.330 2211.690 2567.510 2212.870 ;
        RECT 2567.930 2211.690 2569.110 2212.870 ;
        RECT 2566.330 2033.290 2567.510 2034.470 ;
        RECT 2567.930 2033.290 2569.110 2034.470 ;
        RECT 2566.330 2031.690 2567.510 2032.870 ;
        RECT 2567.930 2031.690 2569.110 2032.870 ;
        RECT 2566.330 1853.290 2567.510 1854.470 ;
        RECT 2567.930 1853.290 2569.110 1854.470 ;
        RECT 2566.330 1851.690 2567.510 1852.870 ;
        RECT 2567.930 1851.690 2569.110 1852.870 ;
        RECT 2566.330 1673.290 2567.510 1674.470 ;
        RECT 2567.930 1673.290 2569.110 1674.470 ;
        RECT 2566.330 1671.690 2567.510 1672.870 ;
        RECT 2567.930 1671.690 2569.110 1672.870 ;
        RECT 2566.330 1493.290 2567.510 1494.470 ;
        RECT 2567.930 1493.290 2569.110 1494.470 ;
        RECT 2566.330 1491.690 2567.510 1492.870 ;
        RECT 2567.930 1491.690 2569.110 1492.870 ;
        RECT 2566.330 1313.290 2567.510 1314.470 ;
        RECT 2567.930 1313.290 2569.110 1314.470 ;
        RECT 2566.330 1311.690 2567.510 1312.870 ;
        RECT 2567.930 1311.690 2569.110 1312.870 ;
        RECT 2566.330 1133.290 2567.510 1134.470 ;
        RECT 2567.930 1133.290 2569.110 1134.470 ;
        RECT 2566.330 1131.690 2567.510 1132.870 ;
        RECT 2567.930 1131.690 2569.110 1132.870 ;
        RECT 2566.330 953.290 2567.510 954.470 ;
        RECT 2567.930 953.290 2569.110 954.470 ;
        RECT 2566.330 951.690 2567.510 952.870 ;
        RECT 2567.930 951.690 2569.110 952.870 ;
        RECT 2566.330 773.290 2567.510 774.470 ;
        RECT 2567.930 773.290 2569.110 774.470 ;
        RECT 2566.330 771.690 2567.510 772.870 ;
        RECT 2567.930 771.690 2569.110 772.870 ;
        RECT 2566.330 593.290 2567.510 594.470 ;
        RECT 2567.930 593.290 2569.110 594.470 ;
        RECT 2566.330 591.690 2567.510 592.870 ;
        RECT 2567.930 591.690 2569.110 592.870 ;
        RECT 2566.330 413.290 2567.510 414.470 ;
        RECT 2567.930 413.290 2569.110 414.470 ;
        RECT 2566.330 411.690 2567.510 412.870 ;
        RECT 2567.930 411.690 2569.110 412.870 ;
        RECT 2566.330 233.290 2567.510 234.470 ;
        RECT 2567.930 233.290 2569.110 234.470 ;
        RECT 2566.330 231.690 2567.510 232.870 ;
        RECT 2567.930 231.690 2569.110 232.870 ;
        RECT 2566.330 53.290 2567.510 54.470 ;
        RECT 2567.930 53.290 2569.110 54.470 ;
        RECT 2566.330 51.690 2567.510 52.870 ;
        RECT 2567.930 51.690 2569.110 52.870 ;
        RECT 2566.330 -22.110 2567.510 -20.930 ;
        RECT 2567.930 -22.110 2569.110 -20.930 ;
        RECT 2566.330 -23.710 2567.510 -22.530 ;
        RECT 2567.930 -23.710 2569.110 -22.530 ;
        RECT 2746.330 3542.210 2747.510 3543.390 ;
        RECT 2747.930 3542.210 2749.110 3543.390 ;
        RECT 2746.330 3540.610 2747.510 3541.790 ;
        RECT 2747.930 3540.610 2749.110 3541.790 ;
        RECT 2746.330 3473.290 2747.510 3474.470 ;
        RECT 2747.930 3473.290 2749.110 3474.470 ;
        RECT 2746.330 3471.690 2747.510 3472.870 ;
        RECT 2747.930 3471.690 2749.110 3472.870 ;
        RECT 2746.330 3293.290 2747.510 3294.470 ;
        RECT 2747.930 3293.290 2749.110 3294.470 ;
        RECT 2746.330 3291.690 2747.510 3292.870 ;
        RECT 2747.930 3291.690 2749.110 3292.870 ;
        RECT 2746.330 3113.290 2747.510 3114.470 ;
        RECT 2747.930 3113.290 2749.110 3114.470 ;
        RECT 2746.330 3111.690 2747.510 3112.870 ;
        RECT 2747.930 3111.690 2749.110 3112.870 ;
        RECT 2746.330 2933.290 2747.510 2934.470 ;
        RECT 2747.930 2933.290 2749.110 2934.470 ;
        RECT 2746.330 2931.690 2747.510 2932.870 ;
        RECT 2747.930 2931.690 2749.110 2932.870 ;
        RECT 2746.330 2753.290 2747.510 2754.470 ;
        RECT 2747.930 2753.290 2749.110 2754.470 ;
        RECT 2746.330 2751.690 2747.510 2752.870 ;
        RECT 2747.930 2751.690 2749.110 2752.870 ;
        RECT 2746.330 2573.290 2747.510 2574.470 ;
        RECT 2747.930 2573.290 2749.110 2574.470 ;
        RECT 2746.330 2571.690 2747.510 2572.870 ;
        RECT 2747.930 2571.690 2749.110 2572.870 ;
        RECT 2746.330 2393.290 2747.510 2394.470 ;
        RECT 2747.930 2393.290 2749.110 2394.470 ;
        RECT 2746.330 2391.690 2747.510 2392.870 ;
        RECT 2747.930 2391.690 2749.110 2392.870 ;
        RECT 2746.330 2213.290 2747.510 2214.470 ;
        RECT 2747.930 2213.290 2749.110 2214.470 ;
        RECT 2746.330 2211.690 2747.510 2212.870 ;
        RECT 2747.930 2211.690 2749.110 2212.870 ;
        RECT 2746.330 2033.290 2747.510 2034.470 ;
        RECT 2747.930 2033.290 2749.110 2034.470 ;
        RECT 2746.330 2031.690 2747.510 2032.870 ;
        RECT 2747.930 2031.690 2749.110 2032.870 ;
        RECT 2746.330 1853.290 2747.510 1854.470 ;
        RECT 2747.930 1853.290 2749.110 1854.470 ;
        RECT 2746.330 1851.690 2747.510 1852.870 ;
        RECT 2747.930 1851.690 2749.110 1852.870 ;
        RECT 2746.330 1673.290 2747.510 1674.470 ;
        RECT 2747.930 1673.290 2749.110 1674.470 ;
        RECT 2746.330 1671.690 2747.510 1672.870 ;
        RECT 2747.930 1671.690 2749.110 1672.870 ;
        RECT 2746.330 1493.290 2747.510 1494.470 ;
        RECT 2747.930 1493.290 2749.110 1494.470 ;
        RECT 2746.330 1491.690 2747.510 1492.870 ;
        RECT 2747.930 1491.690 2749.110 1492.870 ;
        RECT 2746.330 1313.290 2747.510 1314.470 ;
        RECT 2747.930 1313.290 2749.110 1314.470 ;
        RECT 2746.330 1311.690 2747.510 1312.870 ;
        RECT 2747.930 1311.690 2749.110 1312.870 ;
        RECT 2746.330 1133.290 2747.510 1134.470 ;
        RECT 2747.930 1133.290 2749.110 1134.470 ;
        RECT 2746.330 1131.690 2747.510 1132.870 ;
        RECT 2747.930 1131.690 2749.110 1132.870 ;
        RECT 2746.330 953.290 2747.510 954.470 ;
        RECT 2747.930 953.290 2749.110 954.470 ;
        RECT 2746.330 951.690 2747.510 952.870 ;
        RECT 2747.930 951.690 2749.110 952.870 ;
        RECT 2746.330 773.290 2747.510 774.470 ;
        RECT 2747.930 773.290 2749.110 774.470 ;
        RECT 2746.330 771.690 2747.510 772.870 ;
        RECT 2747.930 771.690 2749.110 772.870 ;
        RECT 2746.330 593.290 2747.510 594.470 ;
        RECT 2747.930 593.290 2749.110 594.470 ;
        RECT 2746.330 591.690 2747.510 592.870 ;
        RECT 2747.930 591.690 2749.110 592.870 ;
        RECT 2746.330 413.290 2747.510 414.470 ;
        RECT 2747.930 413.290 2749.110 414.470 ;
        RECT 2746.330 411.690 2747.510 412.870 ;
        RECT 2747.930 411.690 2749.110 412.870 ;
        RECT 2746.330 233.290 2747.510 234.470 ;
        RECT 2747.930 233.290 2749.110 234.470 ;
        RECT 2746.330 231.690 2747.510 232.870 ;
        RECT 2747.930 231.690 2749.110 232.870 ;
        RECT 2746.330 53.290 2747.510 54.470 ;
        RECT 2747.930 53.290 2749.110 54.470 ;
        RECT 2746.330 51.690 2747.510 52.870 ;
        RECT 2747.930 51.690 2749.110 52.870 ;
        RECT 2746.330 -22.110 2747.510 -20.930 ;
        RECT 2747.930 -22.110 2749.110 -20.930 ;
        RECT 2746.330 -23.710 2747.510 -22.530 ;
        RECT 2747.930 -23.710 2749.110 -22.530 ;
        RECT 2945.910 3542.210 2947.090 3543.390 ;
        RECT 2947.510 3542.210 2948.690 3543.390 ;
        RECT 2945.910 3540.610 2947.090 3541.790 ;
        RECT 2947.510 3540.610 2948.690 3541.790 ;
        RECT 2945.910 3473.290 2947.090 3474.470 ;
        RECT 2947.510 3473.290 2948.690 3474.470 ;
        RECT 2945.910 3471.690 2947.090 3472.870 ;
        RECT 2947.510 3471.690 2948.690 3472.870 ;
        RECT 2945.910 3293.290 2947.090 3294.470 ;
        RECT 2947.510 3293.290 2948.690 3294.470 ;
        RECT 2945.910 3291.690 2947.090 3292.870 ;
        RECT 2947.510 3291.690 2948.690 3292.870 ;
        RECT 2945.910 3113.290 2947.090 3114.470 ;
        RECT 2947.510 3113.290 2948.690 3114.470 ;
        RECT 2945.910 3111.690 2947.090 3112.870 ;
        RECT 2947.510 3111.690 2948.690 3112.870 ;
        RECT 2945.910 2933.290 2947.090 2934.470 ;
        RECT 2947.510 2933.290 2948.690 2934.470 ;
        RECT 2945.910 2931.690 2947.090 2932.870 ;
        RECT 2947.510 2931.690 2948.690 2932.870 ;
        RECT 2945.910 2753.290 2947.090 2754.470 ;
        RECT 2947.510 2753.290 2948.690 2754.470 ;
        RECT 2945.910 2751.690 2947.090 2752.870 ;
        RECT 2947.510 2751.690 2948.690 2752.870 ;
        RECT 2945.910 2573.290 2947.090 2574.470 ;
        RECT 2947.510 2573.290 2948.690 2574.470 ;
        RECT 2945.910 2571.690 2947.090 2572.870 ;
        RECT 2947.510 2571.690 2948.690 2572.870 ;
        RECT 2945.910 2393.290 2947.090 2394.470 ;
        RECT 2947.510 2393.290 2948.690 2394.470 ;
        RECT 2945.910 2391.690 2947.090 2392.870 ;
        RECT 2947.510 2391.690 2948.690 2392.870 ;
        RECT 2945.910 2213.290 2947.090 2214.470 ;
        RECT 2947.510 2213.290 2948.690 2214.470 ;
        RECT 2945.910 2211.690 2947.090 2212.870 ;
        RECT 2947.510 2211.690 2948.690 2212.870 ;
        RECT 2945.910 2033.290 2947.090 2034.470 ;
        RECT 2947.510 2033.290 2948.690 2034.470 ;
        RECT 2945.910 2031.690 2947.090 2032.870 ;
        RECT 2947.510 2031.690 2948.690 2032.870 ;
        RECT 2945.910 1853.290 2947.090 1854.470 ;
        RECT 2947.510 1853.290 2948.690 1854.470 ;
        RECT 2945.910 1851.690 2947.090 1852.870 ;
        RECT 2947.510 1851.690 2948.690 1852.870 ;
        RECT 2945.910 1673.290 2947.090 1674.470 ;
        RECT 2947.510 1673.290 2948.690 1674.470 ;
        RECT 2945.910 1671.690 2947.090 1672.870 ;
        RECT 2947.510 1671.690 2948.690 1672.870 ;
        RECT 2945.910 1493.290 2947.090 1494.470 ;
        RECT 2947.510 1493.290 2948.690 1494.470 ;
        RECT 2945.910 1491.690 2947.090 1492.870 ;
        RECT 2947.510 1491.690 2948.690 1492.870 ;
        RECT 2945.910 1313.290 2947.090 1314.470 ;
        RECT 2947.510 1313.290 2948.690 1314.470 ;
        RECT 2945.910 1311.690 2947.090 1312.870 ;
        RECT 2947.510 1311.690 2948.690 1312.870 ;
        RECT 2945.910 1133.290 2947.090 1134.470 ;
        RECT 2947.510 1133.290 2948.690 1134.470 ;
        RECT 2945.910 1131.690 2947.090 1132.870 ;
        RECT 2947.510 1131.690 2948.690 1132.870 ;
        RECT 2945.910 953.290 2947.090 954.470 ;
        RECT 2947.510 953.290 2948.690 954.470 ;
        RECT 2945.910 951.690 2947.090 952.870 ;
        RECT 2947.510 951.690 2948.690 952.870 ;
        RECT 2945.910 773.290 2947.090 774.470 ;
        RECT 2947.510 773.290 2948.690 774.470 ;
        RECT 2945.910 771.690 2947.090 772.870 ;
        RECT 2947.510 771.690 2948.690 772.870 ;
        RECT 2945.910 593.290 2947.090 594.470 ;
        RECT 2947.510 593.290 2948.690 594.470 ;
        RECT 2945.910 591.690 2947.090 592.870 ;
        RECT 2947.510 591.690 2948.690 592.870 ;
        RECT 2945.910 413.290 2947.090 414.470 ;
        RECT 2947.510 413.290 2948.690 414.470 ;
        RECT 2945.910 411.690 2947.090 412.870 ;
        RECT 2947.510 411.690 2948.690 412.870 ;
        RECT 2945.910 233.290 2947.090 234.470 ;
        RECT 2947.510 233.290 2948.690 234.470 ;
        RECT 2945.910 231.690 2947.090 232.870 ;
        RECT 2947.510 231.690 2948.690 232.870 ;
        RECT 2945.910 53.290 2947.090 54.470 ;
        RECT 2947.510 53.290 2948.690 54.470 ;
        RECT 2945.910 51.690 2947.090 52.870 ;
        RECT 2947.510 51.690 2948.690 52.870 ;
        RECT 2945.910 -22.110 2947.090 -20.930 ;
        RECT 2947.510 -22.110 2948.690 -20.930 ;
        RECT 2945.910 -23.710 2947.090 -22.530 ;
        RECT 2947.510 -23.710 2948.690 -22.530 ;
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
        RECT -34.030 951.530 2953.650 954.630 ;
        RECT -34.030 771.530 2953.650 774.630 ;
        RECT -34.030 591.530 2953.650 594.630 ;
        RECT -34.030 411.530 2953.650 414.630 ;
        RECT -34.030 231.530 2953.650 234.630 ;
        RECT -34.030 51.530 2953.650 54.630 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
        RECT 244.770 1010.000 247.870 3557.950 ;
        RECT 424.770 1010.000 427.870 3557.950 ;
        RECT 604.770 1010.000 607.870 3557.950 ;
        RECT 784.770 1010.000 787.870 3557.950 ;
        RECT 964.770 1010.000 967.870 3557.950 ;
        RECT 244.770 -38.270 247.870 390.000 ;
        RECT 424.770 -38.270 427.870 390.000 ;
        RECT 604.770 -38.270 607.870 390.000 ;
        RECT 784.770 -38.270 787.870 390.000 ;
        RECT 964.770 -38.270 967.870 390.000 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
        RECT 1684.770 -38.270 1687.870 3557.950 ;
        RECT 1864.770 -38.270 1867.870 3557.950 ;
        RECT 2044.770 -38.270 2047.870 3557.950 ;
        RECT 2224.770 -38.270 2227.870 3557.950 ;
        RECT 2404.770 -38.270 2407.870 3557.950 ;
        RECT 2584.770 -38.270 2587.870 3557.950 ;
        RECT 2764.770 -38.270 2767.870 3557.950 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
      LAYER via4 ;
        RECT -38.670 3551.810 -37.490 3552.990 ;
        RECT -37.070 3551.810 -35.890 3552.990 ;
        RECT -38.670 3550.210 -37.490 3551.390 ;
        RECT -37.070 3550.210 -35.890 3551.390 ;
        RECT -38.670 3491.890 -37.490 3493.070 ;
        RECT -37.070 3491.890 -35.890 3493.070 ;
        RECT -38.670 3490.290 -37.490 3491.470 ;
        RECT -37.070 3490.290 -35.890 3491.470 ;
        RECT -38.670 3311.890 -37.490 3313.070 ;
        RECT -37.070 3311.890 -35.890 3313.070 ;
        RECT -38.670 3310.290 -37.490 3311.470 ;
        RECT -37.070 3310.290 -35.890 3311.470 ;
        RECT -38.670 3131.890 -37.490 3133.070 ;
        RECT -37.070 3131.890 -35.890 3133.070 ;
        RECT -38.670 3130.290 -37.490 3131.470 ;
        RECT -37.070 3130.290 -35.890 3131.470 ;
        RECT -38.670 2951.890 -37.490 2953.070 ;
        RECT -37.070 2951.890 -35.890 2953.070 ;
        RECT -38.670 2950.290 -37.490 2951.470 ;
        RECT -37.070 2950.290 -35.890 2951.470 ;
        RECT -38.670 2771.890 -37.490 2773.070 ;
        RECT -37.070 2771.890 -35.890 2773.070 ;
        RECT -38.670 2770.290 -37.490 2771.470 ;
        RECT -37.070 2770.290 -35.890 2771.470 ;
        RECT -38.670 2591.890 -37.490 2593.070 ;
        RECT -37.070 2591.890 -35.890 2593.070 ;
        RECT -38.670 2590.290 -37.490 2591.470 ;
        RECT -37.070 2590.290 -35.890 2591.470 ;
        RECT -38.670 2411.890 -37.490 2413.070 ;
        RECT -37.070 2411.890 -35.890 2413.070 ;
        RECT -38.670 2410.290 -37.490 2411.470 ;
        RECT -37.070 2410.290 -35.890 2411.470 ;
        RECT -38.670 2231.890 -37.490 2233.070 ;
        RECT -37.070 2231.890 -35.890 2233.070 ;
        RECT -38.670 2230.290 -37.490 2231.470 ;
        RECT -37.070 2230.290 -35.890 2231.470 ;
        RECT -38.670 2051.890 -37.490 2053.070 ;
        RECT -37.070 2051.890 -35.890 2053.070 ;
        RECT -38.670 2050.290 -37.490 2051.470 ;
        RECT -37.070 2050.290 -35.890 2051.470 ;
        RECT -38.670 1871.890 -37.490 1873.070 ;
        RECT -37.070 1871.890 -35.890 1873.070 ;
        RECT -38.670 1870.290 -37.490 1871.470 ;
        RECT -37.070 1870.290 -35.890 1871.470 ;
        RECT -38.670 1691.890 -37.490 1693.070 ;
        RECT -37.070 1691.890 -35.890 1693.070 ;
        RECT -38.670 1690.290 -37.490 1691.470 ;
        RECT -37.070 1690.290 -35.890 1691.470 ;
        RECT -38.670 1511.890 -37.490 1513.070 ;
        RECT -37.070 1511.890 -35.890 1513.070 ;
        RECT -38.670 1510.290 -37.490 1511.470 ;
        RECT -37.070 1510.290 -35.890 1511.470 ;
        RECT -38.670 1331.890 -37.490 1333.070 ;
        RECT -37.070 1331.890 -35.890 1333.070 ;
        RECT -38.670 1330.290 -37.490 1331.470 ;
        RECT -37.070 1330.290 -35.890 1331.470 ;
        RECT -38.670 1151.890 -37.490 1153.070 ;
        RECT -37.070 1151.890 -35.890 1153.070 ;
        RECT -38.670 1150.290 -37.490 1151.470 ;
        RECT -37.070 1150.290 -35.890 1151.470 ;
        RECT -38.670 971.890 -37.490 973.070 ;
        RECT -37.070 971.890 -35.890 973.070 ;
        RECT -38.670 970.290 -37.490 971.470 ;
        RECT -37.070 970.290 -35.890 971.470 ;
        RECT -38.670 791.890 -37.490 793.070 ;
        RECT -37.070 791.890 -35.890 793.070 ;
        RECT -38.670 790.290 -37.490 791.470 ;
        RECT -37.070 790.290 -35.890 791.470 ;
        RECT -38.670 611.890 -37.490 613.070 ;
        RECT -37.070 611.890 -35.890 613.070 ;
        RECT -38.670 610.290 -37.490 611.470 ;
        RECT -37.070 610.290 -35.890 611.470 ;
        RECT -38.670 431.890 -37.490 433.070 ;
        RECT -37.070 431.890 -35.890 433.070 ;
        RECT -38.670 430.290 -37.490 431.470 ;
        RECT -37.070 430.290 -35.890 431.470 ;
        RECT -38.670 251.890 -37.490 253.070 ;
        RECT -37.070 251.890 -35.890 253.070 ;
        RECT -38.670 250.290 -37.490 251.470 ;
        RECT -37.070 250.290 -35.890 251.470 ;
        RECT -38.670 71.890 -37.490 73.070 ;
        RECT -37.070 71.890 -35.890 73.070 ;
        RECT -38.670 70.290 -37.490 71.470 ;
        RECT -37.070 70.290 -35.890 71.470 ;
        RECT -38.670 -31.710 -37.490 -30.530 ;
        RECT -37.070 -31.710 -35.890 -30.530 ;
        RECT -38.670 -33.310 -37.490 -32.130 ;
        RECT -37.070 -33.310 -35.890 -32.130 ;
        RECT 64.930 3551.810 66.110 3552.990 ;
        RECT 66.530 3551.810 67.710 3552.990 ;
        RECT 64.930 3550.210 66.110 3551.390 ;
        RECT 66.530 3550.210 67.710 3551.390 ;
        RECT 64.930 3491.890 66.110 3493.070 ;
        RECT 66.530 3491.890 67.710 3493.070 ;
        RECT 64.930 3490.290 66.110 3491.470 ;
        RECT 66.530 3490.290 67.710 3491.470 ;
        RECT 64.930 3311.890 66.110 3313.070 ;
        RECT 66.530 3311.890 67.710 3313.070 ;
        RECT 64.930 3310.290 66.110 3311.470 ;
        RECT 66.530 3310.290 67.710 3311.470 ;
        RECT 64.930 3131.890 66.110 3133.070 ;
        RECT 66.530 3131.890 67.710 3133.070 ;
        RECT 64.930 3130.290 66.110 3131.470 ;
        RECT 66.530 3130.290 67.710 3131.470 ;
        RECT 64.930 2951.890 66.110 2953.070 ;
        RECT 66.530 2951.890 67.710 2953.070 ;
        RECT 64.930 2950.290 66.110 2951.470 ;
        RECT 66.530 2950.290 67.710 2951.470 ;
        RECT 64.930 2771.890 66.110 2773.070 ;
        RECT 66.530 2771.890 67.710 2773.070 ;
        RECT 64.930 2770.290 66.110 2771.470 ;
        RECT 66.530 2770.290 67.710 2771.470 ;
        RECT 64.930 2591.890 66.110 2593.070 ;
        RECT 66.530 2591.890 67.710 2593.070 ;
        RECT 64.930 2590.290 66.110 2591.470 ;
        RECT 66.530 2590.290 67.710 2591.470 ;
        RECT 64.930 2411.890 66.110 2413.070 ;
        RECT 66.530 2411.890 67.710 2413.070 ;
        RECT 64.930 2410.290 66.110 2411.470 ;
        RECT 66.530 2410.290 67.710 2411.470 ;
        RECT 64.930 2231.890 66.110 2233.070 ;
        RECT 66.530 2231.890 67.710 2233.070 ;
        RECT 64.930 2230.290 66.110 2231.470 ;
        RECT 66.530 2230.290 67.710 2231.470 ;
        RECT 64.930 2051.890 66.110 2053.070 ;
        RECT 66.530 2051.890 67.710 2053.070 ;
        RECT 64.930 2050.290 66.110 2051.470 ;
        RECT 66.530 2050.290 67.710 2051.470 ;
        RECT 64.930 1871.890 66.110 1873.070 ;
        RECT 66.530 1871.890 67.710 1873.070 ;
        RECT 64.930 1870.290 66.110 1871.470 ;
        RECT 66.530 1870.290 67.710 1871.470 ;
        RECT 64.930 1691.890 66.110 1693.070 ;
        RECT 66.530 1691.890 67.710 1693.070 ;
        RECT 64.930 1690.290 66.110 1691.470 ;
        RECT 66.530 1690.290 67.710 1691.470 ;
        RECT 64.930 1511.890 66.110 1513.070 ;
        RECT 66.530 1511.890 67.710 1513.070 ;
        RECT 64.930 1510.290 66.110 1511.470 ;
        RECT 66.530 1510.290 67.710 1511.470 ;
        RECT 64.930 1331.890 66.110 1333.070 ;
        RECT 66.530 1331.890 67.710 1333.070 ;
        RECT 64.930 1330.290 66.110 1331.470 ;
        RECT 66.530 1330.290 67.710 1331.470 ;
        RECT 64.930 1151.890 66.110 1153.070 ;
        RECT 66.530 1151.890 67.710 1153.070 ;
        RECT 64.930 1150.290 66.110 1151.470 ;
        RECT 66.530 1150.290 67.710 1151.470 ;
        RECT 244.930 3551.810 246.110 3552.990 ;
        RECT 246.530 3551.810 247.710 3552.990 ;
        RECT 244.930 3550.210 246.110 3551.390 ;
        RECT 246.530 3550.210 247.710 3551.390 ;
        RECT 244.930 3491.890 246.110 3493.070 ;
        RECT 246.530 3491.890 247.710 3493.070 ;
        RECT 244.930 3490.290 246.110 3491.470 ;
        RECT 246.530 3490.290 247.710 3491.470 ;
        RECT 244.930 3311.890 246.110 3313.070 ;
        RECT 246.530 3311.890 247.710 3313.070 ;
        RECT 244.930 3310.290 246.110 3311.470 ;
        RECT 246.530 3310.290 247.710 3311.470 ;
        RECT 244.930 3131.890 246.110 3133.070 ;
        RECT 246.530 3131.890 247.710 3133.070 ;
        RECT 244.930 3130.290 246.110 3131.470 ;
        RECT 246.530 3130.290 247.710 3131.470 ;
        RECT 244.930 2951.890 246.110 2953.070 ;
        RECT 246.530 2951.890 247.710 2953.070 ;
        RECT 244.930 2950.290 246.110 2951.470 ;
        RECT 246.530 2950.290 247.710 2951.470 ;
        RECT 244.930 2771.890 246.110 2773.070 ;
        RECT 246.530 2771.890 247.710 2773.070 ;
        RECT 244.930 2770.290 246.110 2771.470 ;
        RECT 246.530 2770.290 247.710 2771.470 ;
        RECT 244.930 2591.890 246.110 2593.070 ;
        RECT 246.530 2591.890 247.710 2593.070 ;
        RECT 244.930 2590.290 246.110 2591.470 ;
        RECT 246.530 2590.290 247.710 2591.470 ;
        RECT 244.930 2411.890 246.110 2413.070 ;
        RECT 246.530 2411.890 247.710 2413.070 ;
        RECT 244.930 2410.290 246.110 2411.470 ;
        RECT 246.530 2410.290 247.710 2411.470 ;
        RECT 244.930 2231.890 246.110 2233.070 ;
        RECT 246.530 2231.890 247.710 2233.070 ;
        RECT 244.930 2230.290 246.110 2231.470 ;
        RECT 246.530 2230.290 247.710 2231.470 ;
        RECT 244.930 2051.890 246.110 2053.070 ;
        RECT 246.530 2051.890 247.710 2053.070 ;
        RECT 244.930 2050.290 246.110 2051.470 ;
        RECT 246.530 2050.290 247.710 2051.470 ;
        RECT 244.930 1871.890 246.110 1873.070 ;
        RECT 246.530 1871.890 247.710 1873.070 ;
        RECT 244.930 1870.290 246.110 1871.470 ;
        RECT 246.530 1870.290 247.710 1871.470 ;
        RECT 244.930 1691.890 246.110 1693.070 ;
        RECT 246.530 1691.890 247.710 1693.070 ;
        RECT 244.930 1690.290 246.110 1691.470 ;
        RECT 246.530 1690.290 247.710 1691.470 ;
        RECT 244.930 1511.890 246.110 1513.070 ;
        RECT 246.530 1511.890 247.710 1513.070 ;
        RECT 244.930 1510.290 246.110 1511.470 ;
        RECT 246.530 1510.290 247.710 1511.470 ;
        RECT 244.930 1331.890 246.110 1333.070 ;
        RECT 246.530 1331.890 247.710 1333.070 ;
        RECT 244.930 1330.290 246.110 1331.470 ;
        RECT 246.530 1330.290 247.710 1331.470 ;
        RECT 244.930 1151.890 246.110 1153.070 ;
        RECT 246.530 1151.890 247.710 1153.070 ;
        RECT 244.930 1150.290 246.110 1151.470 ;
        RECT 246.530 1150.290 247.710 1151.470 ;
        RECT 424.930 3551.810 426.110 3552.990 ;
        RECT 426.530 3551.810 427.710 3552.990 ;
        RECT 424.930 3550.210 426.110 3551.390 ;
        RECT 426.530 3550.210 427.710 3551.390 ;
        RECT 424.930 3491.890 426.110 3493.070 ;
        RECT 426.530 3491.890 427.710 3493.070 ;
        RECT 424.930 3490.290 426.110 3491.470 ;
        RECT 426.530 3490.290 427.710 3491.470 ;
        RECT 424.930 3311.890 426.110 3313.070 ;
        RECT 426.530 3311.890 427.710 3313.070 ;
        RECT 424.930 3310.290 426.110 3311.470 ;
        RECT 426.530 3310.290 427.710 3311.470 ;
        RECT 424.930 3131.890 426.110 3133.070 ;
        RECT 426.530 3131.890 427.710 3133.070 ;
        RECT 424.930 3130.290 426.110 3131.470 ;
        RECT 426.530 3130.290 427.710 3131.470 ;
        RECT 424.930 2951.890 426.110 2953.070 ;
        RECT 426.530 2951.890 427.710 2953.070 ;
        RECT 424.930 2950.290 426.110 2951.470 ;
        RECT 426.530 2950.290 427.710 2951.470 ;
        RECT 424.930 2771.890 426.110 2773.070 ;
        RECT 426.530 2771.890 427.710 2773.070 ;
        RECT 424.930 2770.290 426.110 2771.470 ;
        RECT 426.530 2770.290 427.710 2771.470 ;
        RECT 424.930 2591.890 426.110 2593.070 ;
        RECT 426.530 2591.890 427.710 2593.070 ;
        RECT 424.930 2590.290 426.110 2591.470 ;
        RECT 426.530 2590.290 427.710 2591.470 ;
        RECT 424.930 2411.890 426.110 2413.070 ;
        RECT 426.530 2411.890 427.710 2413.070 ;
        RECT 424.930 2410.290 426.110 2411.470 ;
        RECT 426.530 2410.290 427.710 2411.470 ;
        RECT 424.930 2231.890 426.110 2233.070 ;
        RECT 426.530 2231.890 427.710 2233.070 ;
        RECT 424.930 2230.290 426.110 2231.470 ;
        RECT 426.530 2230.290 427.710 2231.470 ;
        RECT 424.930 2051.890 426.110 2053.070 ;
        RECT 426.530 2051.890 427.710 2053.070 ;
        RECT 424.930 2050.290 426.110 2051.470 ;
        RECT 426.530 2050.290 427.710 2051.470 ;
        RECT 424.930 1871.890 426.110 1873.070 ;
        RECT 426.530 1871.890 427.710 1873.070 ;
        RECT 424.930 1870.290 426.110 1871.470 ;
        RECT 426.530 1870.290 427.710 1871.470 ;
        RECT 424.930 1691.890 426.110 1693.070 ;
        RECT 426.530 1691.890 427.710 1693.070 ;
        RECT 424.930 1690.290 426.110 1691.470 ;
        RECT 426.530 1690.290 427.710 1691.470 ;
        RECT 424.930 1511.890 426.110 1513.070 ;
        RECT 426.530 1511.890 427.710 1513.070 ;
        RECT 424.930 1510.290 426.110 1511.470 ;
        RECT 426.530 1510.290 427.710 1511.470 ;
        RECT 424.930 1331.890 426.110 1333.070 ;
        RECT 426.530 1331.890 427.710 1333.070 ;
        RECT 424.930 1330.290 426.110 1331.470 ;
        RECT 426.530 1330.290 427.710 1331.470 ;
        RECT 424.930 1151.890 426.110 1153.070 ;
        RECT 426.530 1151.890 427.710 1153.070 ;
        RECT 424.930 1150.290 426.110 1151.470 ;
        RECT 426.530 1150.290 427.710 1151.470 ;
        RECT 604.930 3551.810 606.110 3552.990 ;
        RECT 606.530 3551.810 607.710 3552.990 ;
        RECT 604.930 3550.210 606.110 3551.390 ;
        RECT 606.530 3550.210 607.710 3551.390 ;
        RECT 604.930 3491.890 606.110 3493.070 ;
        RECT 606.530 3491.890 607.710 3493.070 ;
        RECT 604.930 3490.290 606.110 3491.470 ;
        RECT 606.530 3490.290 607.710 3491.470 ;
        RECT 604.930 3311.890 606.110 3313.070 ;
        RECT 606.530 3311.890 607.710 3313.070 ;
        RECT 604.930 3310.290 606.110 3311.470 ;
        RECT 606.530 3310.290 607.710 3311.470 ;
        RECT 604.930 3131.890 606.110 3133.070 ;
        RECT 606.530 3131.890 607.710 3133.070 ;
        RECT 604.930 3130.290 606.110 3131.470 ;
        RECT 606.530 3130.290 607.710 3131.470 ;
        RECT 604.930 2951.890 606.110 2953.070 ;
        RECT 606.530 2951.890 607.710 2953.070 ;
        RECT 604.930 2950.290 606.110 2951.470 ;
        RECT 606.530 2950.290 607.710 2951.470 ;
        RECT 604.930 2771.890 606.110 2773.070 ;
        RECT 606.530 2771.890 607.710 2773.070 ;
        RECT 604.930 2770.290 606.110 2771.470 ;
        RECT 606.530 2770.290 607.710 2771.470 ;
        RECT 604.930 2591.890 606.110 2593.070 ;
        RECT 606.530 2591.890 607.710 2593.070 ;
        RECT 604.930 2590.290 606.110 2591.470 ;
        RECT 606.530 2590.290 607.710 2591.470 ;
        RECT 604.930 2411.890 606.110 2413.070 ;
        RECT 606.530 2411.890 607.710 2413.070 ;
        RECT 604.930 2410.290 606.110 2411.470 ;
        RECT 606.530 2410.290 607.710 2411.470 ;
        RECT 604.930 2231.890 606.110 2233.070 ;
        RECT 606.530 2231.890 607.710 2233.070 ;
        RECT 604.930 2230.290 606.110 2231.470 ;
        RECT 606.530 2230.290 607.710 2231.470 ;
        RECT 604.930 2051.890 606.110 2053.070 ;
        RECT 606.530 2051.890 607.710 2053.070 ;
        RECT 604.930 2050.290 606.110 2051.470 ;
        RECT 606.530 2050.290 607.710 2051.470 ;
        RECT 604.930 1871.890 606.110 1873.070 ;
        RECT 606.530 1871.890 607.710 1873.070 ;
        RECT 604.930 1870.290 606.110 1871.470 ;
        RECT 606.530 1870.290 607.710 1871.470 ;
        RECT 604.930 1691.890 606.110 1693.070 ;
        RECT 606.530 1691.890 607.710 1693.070 ;
        RECT 604.930 1690.290 606.110 1691.470 ;
        RECT 606.530 1690.290 607.710 1691.470 ;
        RECT 604.930 1511.890 606.110 1513.070 ;
        RECT 606.530 1511.890 607.710 1513.070 ;
        RECT 604.930 1510.290 606.110 1511.470 ;
        RECT 606.530 1510.290 607.710 1511.470 ;
        RECT 604.930 1331.890 606.110 1333.070 ;
        RECT 606.530 1331.890 607.710 1333.070 ;
        RECT 604.930 1330.290 606.110 1331.470 ;
        RECT 606.530 1330.290 607.710 1331.470 ;
        RECT 604.930 1151.890 606.110 1153.070 ;
        RECT 606.530 1151.890 607.710 1153.070 ;
        RECT 604.930 1150.290 606.110 1151.470 ;
        RECT 606.530 1150.290 607.710 1151.470 ;
        RECT 784.930 3551.810 786.110 3552.990 ;
        RECT 786.530 3551.810 787.710 3552.990 ;
        RECT 784.930 3550.210 786.110 3551.390 ;
        RECT 786.530 3550.210 787.710 3551.390 ;
        RECT 784.930 3491.890 786.110 3493.070 ;
        RECT 786.530 3491.890 787.710 3493.070 ;
        RECT 784.930 3490.290 786.110 3491.470 ;
        RECT 786.530 3490.290 787.710 3491.470 ;
        RECT 784.930 3311.890 786.110 3313.070 ;
        RECT 786.530 3311.890 787.710 3313.070 ;
        RECT 784.930 3310.290 786.110 3311.470 ;
        RECT 786.530 3310.290 787.710 3311.470 ;
        RECT 784.930 3131.890 786.110 3133.070 ;
        RECT 786.530 3131.890 787.710 3133.070 ;
        RECT 784.930 3130.290 786.110 3131.470 ;
        RECT 786.530 3130.290 787.710 3131.470 ;
        RECT 784.930 2951.890 786.110 2953.070 ;
        RECT 786.530 2951.890 787.710 2953.070 ;
        RECT 784.930 2950.290 786.110 2951.470 ;
        RECT 786.530 2950.290 787.710 2951.470 ;
        RECT 784.930 2771.890 786.110 2773.070 ;
        RECT 786.530 2771.890 787.710 2773.070 ;
        RECT 784.930 2770.290 786.110 2771.470 ;
        RECT 786.530 2770.290 787.710 2771.470 ;
        RECT 784.930 2591.890 786.110 2593.070 ;
        RECT 786.530 2591.890 787.710 2593.070 ;
        RECT 784.930 2590.290 786.110 2591.470 ;
        RECT 786.530 2590.290 787.710 2591.470 ;
        RECT 784.930 2411.890 786.110 2413.070 ;
        RECT 786.530 2411.890 787.710 2413.070 ;
        RECT 784.930 2410.290 786.110 2411.470 ;
        RECT 786.530 2410.290 787.710 2411.470 ;
        RECT 784.930 2231.890 786.110 2233.070 ;
        RECT 786.530 2231.890 787.710 2233.070 ;
        RECT 784.930 2230.290 786.110 2231.470 ;
        RECT 786.530 2230.290 787.710 2231.470 ;
        RECT 784.930 2051.890 786.110 2053.070 ;
        RECT 786.530 2051.890 787.710 2053.070 ;
        RECT 784.930 2050.290 786.110 2051.470 ;
        RECT 786.530 2050.290 787.710 2051.470 ;
        RECT 784.930 1871.890 786.110 1873.070 ;
        RECT 786.530 1871.890 787.710 1873.070 ;
        RECT 784.930 1870.290 786.110 1871.470 ;
        RECT 786.530 1870.290 787.710 1871.470 ;
        RECT 784.930 1691.890 786.110 1693.070 ;
        RECT 786.530 1691.890 787.710 1693.070 ;
        RECT 784.930 1690.290 786.110 1691.470 ;
        RECT 786.530 1690.290 787.710 1691.470 ;
        RECT 784.930 1511.890 786.110 1513.070 ;
        RECT 786.530 1511.890 787.710 1513.070 ;
        RECT 784.930 1510.290 786.110 1511.470 ;
        RECT 786.530 1510.290 787.710 1511.470 ;
        RECT 784.930 1331.890 786.110 1333.070 ;
        RECT 786.530 1331.890 787.710 1333.070 ;
        RECT 784.930 1330.290 786.110 1331.470 ;
        RECT 786.530 1330.290 787.710 1331.470 ;
        RECT 784.930 1151.890 786.110 1153.070 ;
        RECT 786.530 1151.890 787.710 1153.070 ;
        RECT 784.930 1150.290 786.110 1151.470 ;
        RECT 786.530 1150.290 787.710 1151.470 ;
        RECT 964.930 3551.810 966.110 3552.990 ;
        RECT 966.530 3551.810 967.710 3552.990 ;
        RECT 964.930 3550.210 966.110 3551.390 ;
        RECT 966.530 3550.210 967.710 3551.390 ;
        RECT 964.930 3491.890 966.110 3493.070 ;
        RECT 966.530 3491.890 967.710 3493.070 ;
        RECT 964.930 3490.290 966.110 3491.470 ;
        RECT 966.530 3490.290 967.710 3491.470 ;
        RECT 964.930 3311.890 966.110 3313.070 ;
        RECT 966.530 3311.890 967.710 3313.070 ;
        RECT 964.930 3310.290 966.110 3311.470 ;
        RECT 966.530 3310.290 967.710 3311.470 ;
        RECT 964.930 3131.890 966.110 3133.070 ;
        RECT 966.530 3131.890 967.710 3133.070 ;
        RECT 964.930 3130.290 966.110 3131.470 ;
        RECT 966.530 3130.290 967.710 3131.470 ;
        RECT 964.930 2951.890 966.110 2953.070 ;
        RECT 966.530 2951.890 967.710 2953.070 ;
        RECT 964.930 2950.290 966.110 2951.470 ;
        RECT 966.530 2950.290 967.710 2951.470 ;
        RECT 964.930 2771.890 966.110 2773.070 ;
        RECT 966.530 2771.890 967.710 2773.070 ;
        RECT 964.930 2770.290 966.110 2771.470 ;
        RECT 966.530 2770.290 967.710 2771.470 ;
        RECT 964.930 2591.890 966.110 2593.070 ;
        RECT 966.530 2591.890 967.710 2593.070 ;
        RECT 964.930 2590.290 966.110 2591.470 ;
        RECT 966.530 2590.290 967.710 2591.470 ;
        RECT 964.930 2411.890 966.110 2413.070 ;
        RECT 966.530 2411.890 967.710 2413.070 ;
        RECT 964.930 2410.290 966.110 2411.470 ;
        RECT 966.530 2410.290 967.710 2411.470 ;
        RECT 964.930 2231.890 966.110 2233.070 ;
        RECT 966.530 2231.890 967.710 2233.070 ;
        RECT 964.930 2230.290 966.110 2231.470 ;
        RECT 966.530 2230.290 967.710 2231.470 ;
        RECT 964.930 2051.890 966.110 2053.070 ;
        RECT 966.530 2051.890 967.710 2053.070 ;
        RECT 964.930 2050.290 966.110 2051.470 ;
        RECT 966.530 2050.290 967.710 2051.470 ;
        RECT 964.930 1871.890 966.110 1873.070 ;
        RECT 966.530 1871.890 967.710 1873.070 ;
        RECT 964.930 1870.290 966.110 1871.470 ;
        RECT 966.530 1870.290 967.710 1871.470 ;
        RECT 964.930 1691.890 966.110 1693.070 ;
        RECT 966.530 1691.890 967.710 1693.070 ;
        RECT 964.930 1690.290 966.110 1691.470 ;
        RECT 966.530 1690.290 967.710 1691.470 ;
        RECT 964.930 1511.890 966.110 1513.070 ;
        RECT 966.530 1511.890 967.710 1513.070 ;
        RECT 964.930 1510.290 966.110 1511.470 ;
        RECT 966.530 1510.290 967.710 1511.470 ;
        RECT 964.930 1331.890 966.110 1333.070 ;
        RECT 966.530 1331.890 967.710 1333.070 ;
        RECT 964.930 1330.290 966.110 1331.470 ;
        RECT 966.530 1330.290 967.710 1331.470 ;
        RECT 964.930 1151.890 966.110 1153.070 ;
        RECT 966.530 1151.890 967.710 1153.070 ;
        RECT 964.930 1150.290 966.110 1151.470 ;
        RECT 966.530 1150.290 967.710 1151.470 ;
        RECT 1144.930 3551.810 1146.110 3552.990 ;
        RECT 1146.530 3551.810 1147.710 3552.990 ;
        RECT 1144.930 3550.210 1146.110 3551.390 ;
        RECT 1146.530 3550.210 1147.710 3551.390 ;
        RECT 1144.930 3491.890 1146.110 3493.070 ;
        RECT 1146.530 3491.890 1147.710 3493.070 ;
        RECT 1144.930 3490.290 1146.110 3491.470 ;
        RECT 1146.530 3490.290 1147.710 3491.470 ;
        RECT 1144.930 3311.890 1146.110 3313.070 ;
        RECT 1146.530 3311.890 1147.710 3313.070 ;
        RECT 1144.930 3310.290 1146.110 3311.470 ;
        RECT 1146.530 3310.290 1147.710 3311.470 ;
        RECT 1144.930 3131.890 1146.110 3133.070 ;
        RECT 1146.530 3131.890 1147.710 3133.070 ;
        RECT 1144.930 3130.290 1146.110 3131.470 ;
        RECT 1146.530 3130.290 1147.710 3131.470 ;
        RECT 1144.930 2951.890 1146.110 2953.070 ;
        RECT 1146.530 2951.890 1147.710 2953.070 ;
        RECT 1144.930 2950.290 1146.110 2951.470 ;
        RECT 1146.530 2950.290 1147.710 2951.470 ;
        RECT 1144.930 2771.890 1146.110 2773.070 ;
        RECT 1146.530 2771.890 1147.710 2773.070 ;
        RECT 1144.930 2770.290 1146.110 2771.470 ;
        RECT 1146.530 2770.290 1147.710 2771.470 ;
        RECT 1144.930 2591.890 1146.110 2593.070 ;
        RECT 1146.530 2591.890 1147.710 2593.070 ;
        RECT 1144.930 2590.290 1146.110 2591.470 ;
        RECT 1146.530 2590.290 1147.710 2591.470 ;
        RECT 1144.930 2411.890 1146.110 2413.070 ;
        RECT 1146.530 2411.890 1147.710 2413.070 ;
        RECT 1144.930 2410.290 1146.110 2411.470 ;
        RECT 1146.530 2410.290 1147.710 2411.470 ;
        RECT 1144.930 2231.890 1146.110 2233.070 ;
        RECT 1146.530 2231.890 1147.710 2233.070 ;
        RECT 1144.930 2230.290 1146.110 2231.470 ;
        RECT 1146.530 2230.290 1147.710 2231.470 ;
        RECT 1144.930 2051.890 1146.110 2053.070 ;
        RECT 1146.530 2051.890 1147.710 2053.070 ;
        RECT 1144.930 2050.290 1146.110 2051.470 ;
        RECT 1146.530 2050.290 1147.710 2051.470 ;
        RECT 1144.930 1871.890 1146.110 1873.070 ;
        RECT 1146.530 1871.890 1147.710 1873.070 ;
        RECT 1144.930 1870.290 1146.110 1871.470 ;
        RECT 1146.530 1870.290 1147.710 1871.470 ;
        RECT 1144.930 1691.890 1146.110 1693.070 ;
        RECT 1146.530 1691.890 1147.710 1693.070 ;
        RECT 1144.930 1690.290 1146.110 1691.470 ;
        RECT 1146.530 1690.290 1147.710 1691.470 ;
        RECT 1144.930 1511.890 1146.110 1513.070 ;
        RECT 1146.530 1511.890 1147.710 1513.070 ;
        RECT 1144.930 1510.290 1146.110 1511.470 ;
        RECT 1146.530 1510.290 1147.710 1511.470 ;
        RECT 1144.930 1331.890 1146.110 1333.070 ;
        RECT 1146.530 1331.890 1147.710 1333.070 ;
        RECT 1144.930 1330.290 1146.110 1331.470 ;
        RECT 1146.530 1330.290 1147.710 1331.470 ;
        RECT 1144.930 1151.890 1146.110 1153.070 ;
        RECT 1146.530 1151.890 1147.710 1153.070 ;
        RECT 1144.930 1150.290 1146.110 1151.470 ;
        RECT 1146.530 1150.290 1147.710 1151.470 ;
        RECT 64.930 971.890 66.110 973.070 ;
        RECT 66.530 971.890 67.710 973.070 ;
        RECT 64.930 970.290 66.110 971.470 ;
        RECT 66.530 970.290 67.710 971.470 ;
        RECT 64.930 791.890 66.110 793.070 ;
        RECT 66.530 791.890 67.710 793.070 ;
        RECT 64.930 790.290 66.110 791.470 ;
        RECT 66.530 790.290 67.710 791.470 ;
        RECT 64.930 611.890 66.110 613.070 ;
        RECT 66.530 611.890 67.710 613.070 ;
        RECT 64.930 610.290 66.110 611.470 ;
        RECT 66.530 610.290 67.710 611.470 ;
        RECT 64.930 431.890 66.110 433.070 ;
        RECT 66.530 431.890 67.710 433.070 ;
        RECT 64.930 430.290 66.110 431.470 ;
        RECT 66.530 430.290 67.710 431.470 ;
        RECT 1144.930 971.890 1146.110 973.070 ;
        RECT 1146.530 971.890 1147.710 973.070 ;
        RECT 1144.930 970.290 1146.110 971.470 ;
        RECT 1146.530 970.290 1147.710 971.470 ;
        RECT 1144.930 791.890 1146.110 793.070 ;
        RECT 1146.530 791.890 1147.710 793.070 ;
        RECT 1144.930 790.290 1146.110 791.470 ;
        RECT 1146.530 790.290 1147.710 791.470 ;
        RECT 1144.930 611.890 1146.110 613.070 ;
        RECT 1146.530 611.890 1147.710 613.070 ;
        RECT 1144.930 610.290 1146.110 611.470 ;
        RECT 1146.530 610.290 1147.710 611.470 ;
        RECT 1144.930 431.890 1146.110 433.070 ;
        RECT 1146.530 431.890 1147.710 433.070 ;
        RECT 1144.930 430.290 1146.110 431.470 ;
        RECT 1146.530 430.290 1147.710 431.470 ;
        RECT 64.930 251.890 66.110 253.070 ;
        RECT 66.530 251.890 67.710 253.070 ;
        RECT 64.930 250.290 66.110 251.470 ;
        RECT 66.530 250.290 67.710 251.470 ;
        RECT 64.930 71.890 66.110 73.070 ;
        RECT 66.530 71.890 67.710 73.070 ;
        RECT 64.930 70.290 66.110 71.470 ;
        RECT 66.530 70.290 67.710 71.470 ;
        RECT 64.930 -31.710 66.110 -30.530 ;
        RECT 66.530 -31.710 67.710 -30.530 ;
        RECT 64.930 -33.310 66.110 -32.130 ;
        RECT 66.530 -33.310 67.710 -32.130 ;
        RECT 244.930 251.890 246.110 253.070 ;
        RECT 246.530 251.890 247.710 253.070 ;
        RECT 244.930 250.290 246.110 251.470 ;
        RECT 246.530 250.290 247.710 251.470 ;
        RECT 244.930 71.890 246.110 73.070 ;
        RECT 246.530 71.890 247.710 73.070 ;
        RECT 244.930 70.290 246.110 71.470 ;
        RECT 246.530 70.290 247.710 71.470 ;
        RECT 244.930 -31.710 246.110 -30.530 ;
        RECT 246.530 -31.710 247.710 -30.530 ;
        RECT 244.930 -33.310 246.110 -32.130 ;
        RECT 246.530 -33.310 247.710 -32.130 ;
        RECT 424.930 251.890 426.110 253.070 ;
        RECT 426.530 251.890 427.710 253.070 ;
        RECT 424.930 250.290 426.110 251.470 ;
        RECT 426.530 250.290 427.710 251.470 ;
        RECT 424.930 71.890 426.110 73.070 ;
        RECT 426.530 71.890 427.710 73.070 ;
        RECT 424.930 70.290 426.110 71.470 ;
        RECT 426.530 70.290 427.710 71.470 ;
        RECT 424.930 -31.710 426.110 -30.530 ;
        RECT 426.530 -31.710 427.710 -30.530 ;
        RECT 424.930 -33.310 426.110 -32.130 ;
        RECT 426.530 -33.310 427.710 -32.130 ;
        RECT 604.930 251.890 606.110 253.070 ;
        RECT 606.530 251.890 607.710 253.070 ;
        RECT 604.930 250.290 606.110 251.470 ;
        RECT 606.530 250.290 607.710 251.470 ;
        RECT 604.930 71.890 606.110 73.070 ;
        RECT 606.530 71.890 607.710 73.070 ;
        RECT 604.930 70.290 606.110 71.470 ;
        RECT 606.530 70.290 607.710 71.470 ;
        RECT 604.930 -31.710 606.110 -30.530 ;
        RECT 606.530 -31.710 607.710 -30.530 ;
        RECT 604.930 -33.310 606.110 -32.130 ;
        RECT 606.530 -33.310 607.710 -32.130 ;
        RECT 784.930 251.890 786.110 253.070 ;
        RECT 786.530 251.890 787.710 253.070 ;
        RECT 784.930 250.290 786.110 251.470 ;
        RECT 786.530 250.290 787.710 251.470 ;
        RECT 784.930 71.890 786.110 73.070 ;
        RECT 786.530 71.890 787.710 73.070 ;
        RECT 784.930 70.290 786.110 71.470 ;
        RECT 786.530 70.290 787.710 71.470 ;
        RECT 784.930 -31.710 786.110 -30.530 ;
        RECT 786.530 -31.710 787.710 -30.530 ;
        RECT 784.930 -33.310 786.110 -32.130 ;
        RECT 786.530 -33.310 787.710 -32.130 ;
        RECT 964.930 251.890 966.110 253.070 ;
        RECT 966.530 251.890 967.710 253.070 ;
        RECT 964.930 250.290 966.110 251.470 ;
        RECT 966.530 250.290 967.710 251.470 ;
        RECT 964.930 71.890 966.110 73.070 ;
        RECT 966.530 71.890 967.710 73.070 ;
        RECT 964.930 70.290 966.110 71.470 ;
        RECT 966.530 70.290 967.710 71.470 ;
        RECT 964.930 -31.710 966.110 -30.530 ;
        RECT 966.530 -31.710 967.710 -30.530 ;
        RECT 964.930 -33.310 966.110 -32.130 ;
        RECT 966.530 -33.310 967.710 -32.130 ;
        RECT 1144.930 251.890 1146.110 253.070 ;
        RECT 1146.530 251.890 1147.710 253.070 ;
        RECT 1144.930 250.290 1146.110 251.470 ;
        RECT 1146.530 250.290 1147.710 251.470 ;
        RECT 1144.930 71.890 1146.110 73.070 ;
        RECT 1146.530 71.890 1147.710 73.070 ;
        RECT 1144.930 70.290 1146.110 71.470 ;
        RECT 1146.530 70.290 1147.710 71.470 ;
        RECT 1144.930 -31.710 1146.110 -30.530 ;
        RECT 1146.530 -31.710 1147.710 -30.530 ;
        RECT 1144.930 -33.310 1146.110 -32.130 ;
        RECT 1146.530 -33.310 1147.710 -32.130 ;
        RECT 1324.930 3551.810 1326.110 3552.990 ;
        RECT 1326.530 3551.810 1327.710 3552.990 ;
        RECT 1324.930 3550.210 1326.110 3551.390 ;
        RECT 1326.530 3550.210 1327.710 3551.390 ;
        RECT 1324.930 3491.890 1326.110 3493.070 ;
        RECT 1326.530 3491.890 1327.710 3493.070 ;
        RECT 1324.930 3490.290 1326.110 3491.470 ;
        RECT 1326.530 3490.290 1327.710 3491.470 ;
        RECT 1324.930 3311.890 1326.110 3313.070 ;
        RECT 1326.530 3311.890 1327.710 3313.070 ;
        RECT 1324.930 3310.290 1326.110 3311.470 ;
        RECT 1326.530 3310.290 1327.710 3311.470 ;
        RECT 1324.930 3131.890 1326.110 3133.070 ;
        RECT 1326.530 3131.890 1327.710 3133.070 ;
        RECT 1324.930 3130.290 1326.110 3131.470 ;
        RECT 1326.530 3130.290 1327.710 3131.470 ;
        RECT 1324.930 2951.890 1326.110 2953.070 ;
        RECT 1326.530 2951.890 1327.710 2953.070 ;
        RECT 1324.930 2950.290 1326.110 2951.470 ;
        RECT 1326.530 2950.290 1327.710 2951.470 ;
        RECT 1324.930 2771.890 1326.110 2773.070 ;
        RECT 1326.530 2771.890 1327.710 2773.070 ;
        RECT 1324.930 2770.290 1326.110 2771.470 ;
        RECT 1326.530 2770.290 1327.710 2771.470 ;
        RECT 1324.930 2591.890 1326.110 2593.070 ;
        RECT 1326.530 2591.890 1327.710 2593.070 ;
        RECT 1324.930 2590.290 1326.110 2591.470 ;
        RECT 1326.530 2590.290 1327.710 2591.470 ;
        RECT 1324.930 2411.890 1326.110 2413.070 ;
        RECT 1326.530 2411.890 1327.710 2413.070 ;
        RECT 1324.930 2410.290 1326.110 2411.470 ;
        RECT 1326.530 2410.290 1327.710 2411.470 ;
        RECT 1324.930 2231.890 1326.110 2233.070 ;
        RECT 1326.530 2231.890 1327.710 2233.070 ;
        RECT 1324.930 2230.290 1326.110 2231.470 ;
        RECT 1326.530 2230.290 1327.710 2231.470 ;
        RECT 1324.930 2051.890 1326.110 2053.070 ;
        RECT 1326.530 2051.890 1327.710 2053.070 ;
        RECT 1324.930 2050.290 1326.110 2051.470 ;
        RECT 1326.530 2050.290 1327.710 2051.470 ;
        RECT 1324.930 1871.890 1326.110 1873.070 ;
        RECT 1326.530 1871.890 1327.710 1873.070 ;
        RECT 1324.930 1870.290 1326.110 1871.470 ;
        RECT 1326.530 1870.290 1327.710 1871.470 ;
        RECT 1324.930 1691.890 1326.110 1693.070 ;
        RECT 1326.530 1691.890 1327.710 1693.070 ;
        RECT 1324.930 1690.290 1326.110 1691.470 ;
        RECT 1326.530 1690.290 1327.710 1691.470 ;
        RECT 1324.930 1511.890 1326.110 1513.070 ;
        RECT 1326.530 1511.890 1327.710 1513.070 ;
        RECT 1324.930 1510.290 1326.110 1511.470 ;
        RECT 1326.530 1510.290 1327.710 1511.470 ;
        RECT 1324.930 1331.890 1326.110 1333.070 ;
        RECT 1326.530 1331.890 1327.710 1333.070 ;
        RECT 1324.930 1330.290 1326.110 1331.470 ;
        RECT 1326.530 1330.290 1327.710 1331.470 ;
        RECT 1324.930 1151.890 1326.110 1153.070 ;
        RECT 1326.530 1151.890 1327.710 1153.070 ;
        RECT 1324.930 1150.290 1326.110 1151.470 ;
        RECT 1326.530 1150.290 1327.710 1151.470 ;
        RECT 1324.930 971.890 1326.110 973.070 ;
        RECT 1326.530 971.890 1327.710 973.070 ;
        RECT 1324.930 970.290 1326.110 971.470 ;
        RECT 1326.530 970.290 1327.710 971.470 ;
        RECT 1324.930 791.890 1326.110 793.070 ;
        RECT 1326.530 791.890 1327.710 793.070 ;
        RECT 1324.930 790.290 1326.110 791.470 ;
        RECT 1326.530 790.290 1327.710 791.470 ;
        RECT 1324.930 611.890 1326.110 613.070 ;
        RECT 1326.530 611.890 1327.710 613.070 ;
        RECT 1324.930 610.290 1326.110 611.470 ;
        RECT 1326.530 610.290 1327.710 611.470 ;
        RECT 1324.930 431.890 1326.110 433.070 ;
        RECT 1326.530 431.890 1327.710 433.070 ;
        RECT 1324.930 430.290 1326.110 431.470 ;
        RECT 1326.530 430.290 1327.710 431.470 ;
        RECT 1324.930 251.890 1326.110 253.070 ;
        RECT 1326.530 251.890 1327.710 253.070 ;
        RECT 1324.930 250.290 1326.110 251.470 ;
        RECT 1326.530 250.290 1327.710 251.470 ;
        RECT 1324.930 71.890 1326.110 73.070 ;
        RECT 1326.530 71.890 1327.710 73.070 ;
        RECT 1324.930 70.290 1326.110 71.470 ;
        RECT 1326.530 70.290 1327.710 71.470 ;
        RECT 1324.930 -31.710 1326.110 -30.530 ;
        RECT 1326.530 -31.710 1327.710 -30.530 ;
        RECT 1324.930 -33.310 1326.110 -32.130 ;
        RECT 1326.530 -33.310 1327.710 -32.130 ;
        RECT 1504.930 3551.810 1506.110 3552.990 ;
        RECT 1506.530 3551.810 1507.710 3552.990 ;
        RECT 1504.930 3550.210 1506.110 3551.390 ;
        RECT 1506.530 3550.210 1507.710 3551.390 ;
        RECT 1504.930 3491.890 1506.110 3493.070 ;
        RECT 1506.530 3491.890 1507.710 3493.070 ;
        RECT 1504.930 3490.290 1506.110 3491.470 ;
        RECT 1506.530 3490.290 1507.710 3491.470 ;
        RECT 1504.930 3311.890 1506.110 3313.070 ;
        RECT 1506.530 3311.890 1507.710 3313.070 ;
        RECT 1504.930 3310.290 1506.110 3311.470 ;
        RECT 1506.530 3310.290 1507.710 3311.470 ;
        RECT 1504.930 3131.890 1506.110 3133.070 ;
        RECT 1506.530 3131.890 1507.710 3133.070 ;
        RECT 1504.930 3130.290 1506.110 3131.470 ;
        RECT 1506.530 3130.290 1507.710 3131.470 ;
        RECT 1504.930 2951.890 1506.110 2953.070 ;
        RECT 1506.530 2951.890 1507.710 2953.070 ;
        RECT 1504.930 2950.290 1506.110 2951.470 ;
        RECT 1506.530 2950.290 1507.710 2951.470 ;
        RECT 1504.930 2771.890 1506.110 2773.070 ;
        RECT 1506.530 2771.890 1507.710 2773.070 ;
        RECT 1504.930 2770.290 1506.110 2771.470 ;
        RECT 1506.530 2770.290 1507.710 2771.470 ;
        RECT 1504.930 2591.890 1506.110 2593.070 ;
        RECT 1506.530 2591.890 1507.710 2593.070 ;
        RECT 1504.930 2590.290 1506.110 2591.470 ;
        RECT 1506.530 2590.290 1507.710 2591.470 ;
        RECT 1504.930 2411.890 1506.110 2413.070 ;
        RECT 1506.530 2411.890 1507.710 2413.070 ;
        RECT 1504.930 2410.290 1506.110 2411.470 ;
        RECT 1506.530 2410.290 1507.710 2411.470 ;
        RECT 1504.930 2231.890 1506.110 2233.070 ;
        RECT 1506.530 2231.890 1507.710 2233.070 ;
        RECT 1504.930 2230.290 1506.110 2231.470 ;
        RECT 1506.530 2230.290 1507.710 2231.470 ;
        RECT 1504.930 2051.890 1506.110 2053.070 ;
        RECT 1506.530 2051.890 1507.710 2053.070 ;
        RECT 1504.930 2050.290 1506.110 2051.470 ;
        RECT 1506.530 2050.290 1507.710 2051.470 ;
        RECT 1504.930 1871.890 1506.110 1873.070 ;
        RECT 1506.530 1871.890 1507.710 1873.070 ;
        RECT 1504.930 1870.290 1506.110 1871.470 ;
        RECT 1506.530 1870.290 1507.710 1871.470 ;
        RECT 1504.930 1691.890 1506.110 1693.070 ;
        RECT 1506.530 1691.890 1507.710 1693.070 ;
        RECT 1504.930 1690.290 1506.110 1691.470 ;
        RECT 1506.530 1690.290 1507.710 1691.470 ;
        RECT 1504.930 1511.890 1506.110 1513.070 ;
        RECT 1506.530 1511.890 1507.710 1513.070 ;
        RECT 1504.930 1510.290 1506.110 1511.470 ;
        RECT 1506.530 1510.290 1507.710 1511.470 ;
        RECT 1504.930 1331.890 1506.110 1333.070 ;
        RECT 1506.530 1331.890 1507.710 1333.070 ;
        RECT 1504.930 1330.290 1506.110 1331.470 ;
        RECT 1506.530 1330.290 1507.710 1331.470 ;
        RECT 1504.930 1151.890 1506.110 1153.070 ;
        RECT 1506.530 1151.890 1507.710 1153.070 ;
        RECT 1504.930 1150.290 1506.110 1151.470 ;
        RECT 1506.530 1150.290 1507.710 1151.470 ;
        RECT 1504.930 971.890 1506.110 973.070 ;
        RECT 1506.530 971.890 1507.710 973.070 ;
        RECT 1504.930 970.290 1506.110 971.470 ;
        RECT 1506.530 970.290 1507.710 971.470 ;
        RECT 1504.930 791.890 1506.110 793.070 ;
        RECT 1506.530 791.890 1507.710 793.070 ;
        RECT 1504.930 790.290 1506.110 791.470 ;
        RECT 1506.530 790.290 1507.710 791.470 ;
        RECT 1504.930 611.890 1506.110 613.070 ;
        RECT 1506.530 611.890 1507.710 613.070 ;
        RECT 1504.930 610.290 1506.110 611.470 ;
        RECT 1506.530 610.290 1507.710 611.470 ;
        RECT 1504.930 431.890 1506.110 433.070 ;
        RECT 1506.530 431.890 1507.710 433.070 ;
        RECT 1504.930 430.290 1506.110 431.470 ;
        RECT 1506.530 430.290 1507.710 431.470 ;
        RECT 1504.930 251.890 1506.110 253.070 ;
        RECT 1506.530 251.890 1507.710 253.070 ;
        RECT 1504.930 250.290 1506.110 251.470 ;
        RECT 1506.530 250.290 1507.710 251.470 ;
        RECT 1504.930 71.890 1506.110 73.070 ;
        RECT 1506.530 71.890 1507.710 73.070 ;
        RECT 1504.930 70.290 1506.110 71.470 ;
        RECT 1506.530 70.290 1507.710 71.470 ;
        RECT 1504.930 -31.710 1506.110 -30.530 ;
        RECT 1506.530 -31.710 1507.710 -30.530 ;
        RECT 1504.930 -33.310 1506.110 -32.130 ;
        RECT 1506.530 -33.310 1507.710 -32.130 ;
        RECT 1684.930 3551.810 1686.110 3552.990 ;
        RECT 1686.530 3551.810 1687.710 3552.990 ;
        RECT 1684.930 3550.210 1686.110 3551.390 ;
        RECT 1686.530 3550.210 1687.710 3551.390 ;
        RECT 1684.930 3491.890 1686.110 3493.070 ;
        RECT 1686.530 3491.890 1687.710 3493.070 ;
        RECT 1684.930 3490.290 1686.110 3491.470 ;
        RECT 1686.530 3490.290 1687.710 3491.470 ;
        RECT 1684.930 3311.890 1686.110 3313.070 ;
        RECT 1686.530 3311.890 1687.710 3313.070 ;
        RECT 1684.930 3310.290 1686.110 3311.470 ;
        RECT 1686.530 3310.290 1687.710 3311.470 ;
        RECT 1684.930 3131.890 1686.110 3133.070 ;
        RECT 1686.530 3131.890 1687.710 3133.070 ;
        RECT 1684.930 3130.290 1686.110 3131.470 ;
        RECT 1686.530 3130.290 1687.710 3131.470 ;
        RECT 1684.930 2951.890 1686.110 2953.070 ;
        RECT 1686.530 2951.890 1687.710 2953.070 ;
        RECT 1684.930 2950.290 1686.110 2951.470 ;
        RECT 1686.530 2950.290 1687.710 2951.470 ;
        RECT 1684.930 2771.890 1686.110 2773.070 ;
        RECT 1686.530 2771.890 1687.710 2773.070 ;
        RECT 1684.930 2770.290 1686.110 2771.470 ;
        RECT 1686.530 2770.290 1687.710 2771.470 ;
        RECT 1684.930 2591.890 1686.110 2593.070 ;
        RECT 1686.530 2591.890 1687.710 2593.070 ;
        RECT 1684.930 2590.290 1686.110 2591.470 ;
        RECT 1686.530 2590.290 1687.710 2591.470 ;
        RECT 1684.930 2411.890 1686.110 2413.070 ;
        RECT 1686.530 2411.890 1687.710 2413.070 ;
        RECT 1684.930 2410.290 1686.110 2411.470 ;
        RECT 1686.530 2410.290 1687.710 2411.470 ;
        RECT 1684.930 2231.890 1686.110 2233.070 ;
        RECT 1686.530 2231.890 1687.710 2233.070 ;
        RECT 1684.930 2230.290 1686.110 2231.470 ;
        RECT 1686.530 2230.290 1687.710 2231.470 ;
        RECT 1684.930 2051.890 1686.110 2053.070 ;
        RECT 1686.530 2051.890 1687.710 2053.070 ;
        RECT 1684.930 2050.290 1686.110 2051.470 ;
        RECT 1686.530 2050.290 1687.710 2051.470 ;
        RECT 1684.930 1871.890 1686.110 1873.070 ;
        RECT 1686.530 1871.890 1687.710 1873.070 ;
        RECT 1684.930 1870.290 1686.110 1871.470 ;
        RECT 1686.530 1870.290 1687.710 1871.470 ;
        RECT 1684.930 1691.890 1686.110 1693.070 ;
        RECT 1686.530 1691.890 1687.710 1693.070 ;
        RECT 1684.930 1690.290 1686.110 1691.470 ;
        RECT 1686.530 1690.290 1687.710 1691.470 ;
        RECT 1684.930 1511.890 1686.110 1513.070 ;
        RECT 1686.530 1511.890 1687.710 1513.070 ;
        RECT 1684.930 1510.290 1686.110 1511.470 ;
        RECT 1686.530 1510.290 1687.710 1511.470 ;
        RECT 1684.930 1331.890 1686.110 1333.070 ;
        RECT 1686.530 1331.890 1687.710 1333.070 ;
        RECT 1684.930 1330.290 1686.110 1331.470 ;
        RECT 1686.530 1330.290 1687.710 1331.470 ;
        RECT 1684.930 1151.890 1686.110 1153.070 ;
        RECT 1686.530 1151.890 1687.710 1153.070 ;
        RECT 1684.930 1150.290 1686.110 1151.470 ;
        RECT 1686.530 1150.290 1687.710 1151.470 ;
        RECT 1684.930 971.890 1686.110 973.070 ;
        RECT 1686.530 971.890 1687.710 973.070 ;
        RECT 1684.930 970.290 1686.110 971.470 ;
        RECT 1686.530 970.290 1687.710 971.470 ;
        RECT 1684.930 791.890 1686.110 793.070 ;
        RECT 1686.530 791.890 1687.710 793.070 ;
        RECT 1684.930 790.290 1686.110 791.470 ;
        RECT 1686.530 790.290 1687.710 791.470 ;
        RECT 1684.930 611.890 1686.110 613.070 ;
        RECT 1686.530 611.890 1687.710 613.070 ;
        RECT 1684.930 610.290 1686.110 611.470 ;
        RECT 1686.530 610.290 1687.710 611.470 ;
        RECT 1684.930 431.890 1686.110 433.070 ;
        RECT 1686.530 431.890 1687.710 433.070 ;
        RECT 1684.930 430.290 1686.110 431.470 ;
        RECT 1686.530 430.290 1687.710 431.470 ;
        RECT 1684.930 251.890 1686.110 253.070 ;
        RECT 1686.530 251.890 1687.710 253.070 ;
        RECT 1684.930 250.290 1686.110 251.470 ;
        RECT 1686.530 250.290 1687.710 251.470 ;
        RECT 1684.930 71.890 1686.110 73.070 ;
        RECT 1686.530 71.890 1687.710 73.070 ;
        RECT 1684.930 70.290 1686.110 71.470 ;
        RECT 1686.530 70.290 1687.710 71.470 ;
        RECT 1684.930 -31.710 1686.110 -30.530 ;
        RECT 1686.530 -31.710 1687.710 -30.530 ;
        RECT 1684.930 -33.310 1686.110 -32.130 ;
        RECT 1686.530 -33.310 1687.710 -32.130 ;
        RECT 1864.930 3551.810 1866.110 3552.990 ;
        RECT 1866.530 3551.810 1867.710 3552.990 ;
        RECT 1864.930 3550.210 1866.110 3551.390 ;
        RECT 1866.530 3550.210 1867.710 3551.390 ;
        RECT 1864.930 3491.890 1866.110 3493.070 ;
        RECT 1866.530 3491.890 1867.710 3493.070 ;
        RECT 1864.930 3490.290 1866.110 3491.470 ;
        RECT 1866.530 3490.290 1867.710 3491.470 ;
        RECT 1864.930 3311.890 1866.110 3313.070 ;
        RECT 1866.530 3311.890 1867.710 3313.070 ;
        RECT 1864.930 3310.290 1866.110 3311.470 ;
        RECT 1866.530 3310.290 1867.710 3311.470 ;
        RECT 1864.930 3131.890 1866.110 3133.070 ;
        RECT 1866.530 3131.890 1867.710 3133.070 ;
        RECT 1864.930 3130.290 1866.110 3131.470 ;
        RECT 1866.530 3130.290 1867.710 3131.470 ;
        RECT 1864.930 2951.890 1866.110 2953.070 ;
        RECT 1866.530 2951.890 1867.710 2953.070 ;
        RECT 1864.930 2950.290 1866.110 2951.470 ;
        RECT 1866.530 2950.290 1867.710 2951.470 ;
        RECT 1864.930 2771.890 1866.110 2773.070 ;
        RECT 1866.530 2771.890 1867.710 2773.070 ;
        RECT 1864.930 2770.290 1866.110 2771.470 ;
        RECT 1866.530 2770.290 1867.710 2771.470 ;
        RECT 1864.930 2591.890 1866.110 2593.070 ;
        RECT 1866.530 2591.890 1867.710 2593.070 ;
        RECT 1864.930 2590.290 1866.110 2591.470 ;
        RECT 1866.530 2590.290 1867.710 2591.470 ;
        RECT 1864.930 2411.890 1866.110 2413.070 ;
        RECT 1866.530 2411.890 1867.710 2413.070 ;
        RECT 1864.930 2410.290 1866.110 2411.470 ;
        RECT 1866.530 2410.290 1867.710 2411.470 ;
        RECT 1864.930 2231.890 1866.110 2233.070 ;
        RECT 1866.530 2231.890 1867.710 2233.070 ;
        RECT 1864.930 2230.290 1866.110 2231.470 ;
        RECT 1866.530 2230.290 1867.710 2231.470 ;
        RECT 1864.930 2051.890 1866.110 2053.070 ;
        RECT 1866.530 2051.890 1867.710 2053.070 ;
        RECT 1864.930 2050.290 1866.110 2051.470 ;
        RECT 1866.530 2050.290 1867.710 2051.470 ;
        RECT 1864.930 1871.890 1866.110 1873.070 ;
        RECT 1866.530 1871.890 1867.710 1873.070 ;
        RECT 1864.930 1870.290 1866.110 1871.470 ;
        RECT 1866.530 1870.290 1867.710 1871.470 ;
        RECT 1864.930 1691.890 1866.110 1693.070 ;
        RECT 1866.530 1691.890 1867.710 1693.070 ;
        RECT 1864.930 1690.290 1866.110 1691.470 ;
        RECT 1866.530 1690.290 1867.710 1691.470 ;
        RECT 1864.930 1511.890 1866.110 1513.070 ;
        RECT 1866.530 1511.890 1867.710 1513.070 ;
        RECT 1864.930 1510.290 1866.110 1511.470 ;
        RECT 1866.530 1510.290 1867.710 1511.470 ;
        RECT 1864.930 1331.890 1866.110 1333.070 ;
        RECT 1866.530 1331.890 1867.710 1333.070 ;
        RECT 1864.930 1330.290 1866.110 1331.470 ;
        RECT 1866.530 1330.290 1867.710 1331.470 ;
        RECT 1864.930 1151.890 1866.110 1153.070 ;
        RECT 1866.530 1151.890 1867.710 1153.070 ;
        RECT 1864.930 1150.290 1866.110 1151.470 ;
        RECT 1866.530 1150.290 1867.710 1151.470 ;
        RECT 1864.930 971.890 1866.110 973.070 ;
        RECT 1866.530 971.890 1867.710 973.070 ;
        RECT 1864.930 970.290 1866.110 971.470 ;
        RECT 1866.530 970.290 1867.710 971.470 ;
        RECT 1864.930 791.890 1866.110 793.070 ;
        RECT 1866.530 791.890 1867.710 793.070 ;
        RECT 1864.930 790.290 1866.110 791.470 ;
        RECT 1866.530 790.290 1867.710 791.470 ;
        RECT 1864.930 611.890 1866.110 613.070 ;
        RECT 1866.530 611.890 1867.710 613.070 ;
        RECT 1864.930 610.290 1866.110 611.470 ;
        RECT 1866.530 610.290 1867.710 611.470 ;
        RECT 1864.930 431.890 1866.110 433.070 ;
        RECT 1866.530 431.890 1867.710 433.070 ;
        RECT 1864.930 430.290 1866.110 431.470 ;
        RECT 1866.530 430.290 1867.710 431.470 ;
        RECT 1864.930 251.890 1866.110 253.070 ;
        RECT 1866.530 251.890 1867.710 253.070 ;
        RECT 1864.930 250.290 1866.110 251.470 ;
        RECT 1866.530 250.290 1867.710 251.470 ;
        RECT 1864.930 71.890 1866.110 73.070 ;
        RECT 1866.530 71.890 1867.710 73.070 ;
        RECT 1864.930 70.290 1866.110 71.470 ;
        RECT 1866.530 70.290 1867.710 71.470 ;
        RECT 1864.930 -31.710 1866.110 -30.530 ;
        RECT 1866.530 -31.710 1867.710 -30.530 ;
        RECT 1864.930 -33.310 1866.110 -32.130 ;
        RECT 1866.530 -33.310 1867.710 -32.130 ;
        RECT 2044.930 3551.810 2046.110 3552.990 ;
        RECT 2046.530 3551.810 2047.710 3552.990 ;
        RECT 2044.930 3550.210 2046.110 3551.390 ;
        RECT 2046.530 3550.210 2047.710 3551.390 ;
        RECT 2044.930 3491.890 2046.110 3493.070 ;
        RECT 2046.530 3491.890 2047.710 3493.070 ;
        RECT 2044.930 3490.290 2046.110 3491.470 ;
        RECT 2046.530 3490.290 2047.710 3491.470 ;
        RECT 2044.930 3311.890 2046.110 3313.070 ;
        RECT 2046.530 3311.890 2047.710 3313.070 ;
        RECT 2044.930 3310.290 2046.110 3311.470 ;
        RECT 2046.530 3310.290 2047.710 3311.470 ;
        RECT 2044.930 3131.890 2046.110 3133.070 ;
        RECT 2046.530 3131.890 2047.710 3133.070 ;
        RECT 2044.930 3130.290 2046.110 3131.470 ;
        RECT 2046.530 3130.290 2047.710 3131.470 ;
        RECT 2044.930 2951.890 2046.110 2953.070 ;
        RECT 2046.530 2951.890 2047.710 2953.070 ;
        RECT 2044.930 2950.290 2046.110 2951.470 ;
        RECT 2046.530 2950.290 2047.710 2951.470 ;
        RECT 2044.930 2771.890 2046.110 2773.070 ;
        RECT 2046.530 2771.890 2047.710 2773.070 ;
        RECT 2044.930 2770.290 2046.110 2771.470 ;
        RECT 2046.530 2770.290 2047.710 2771.470 ;
        RECT 2044.930 2591.890 2046.110 2593.070 ;
        RECT 2046.530 2591.890 2047.710 2593.070 ;
        RECT 2044.930 2590.290 2046.110 2591.470 ;
        RECT 2046.530 2590.290 2047.710 2591.470 ;
        RECT 2044.930 2411.890 2046.110 2413.070 ;
        RECT 2046.530 2411.890 2047.710 2413.070 ;
        RECT 2044.930 2410.290 2046.110 2411.470 ;
        RECT 2046.530 2410.290 2047.710 2411.470 ;
        RECT 2044.930 2231.890 2046.110 2233.070 ;
        RECT 2046.530 2231.890 2047.710 2233.070 ;
        RECT 2044.930 2230.290 2046.110 2231.470 ;
        RECT 2046.530 2230.290 2047.710 2231.470 ;
        RECT 2044.930 2051.890 2046.110 2053.070 ;
        RECT 2046.530 2051.890 2047.710 2053.070 ;
        RECT 2044.930 2050.290 2046.110 2051.470 ;
        RECT 2046.530 2050.290 2047.710 2051.470 ;
        RECT 2044.930 1871.890 2046.110 1873.070 ;
        RECT 2046.530 1871.890 2047.710 1873.070 ;
        RECT 2044.930 1870.290 2046.110 1871.470 ;
        RECT 2046.530 1870.290 2047.710 1871.470 ;
        RECT 2044.930 1691.890 2046.110 1693.070 ;
        RECT 2046.530 1691.890 2047.710 1693.070 ;
        RECT 2044.930 1690.290 2046.110 1691.470 ;
        RECT 2046.530 1690.290 2047.710 1691.470 ;
        RECT 2044.930 1511.890 2046.110 1513.070 ;
        RECT 2046.530 1511.890 2047.710 1513.070 ;
        RECT 2044.930 1510.290 2046.110 1511.470 ;
        RECT 2046.530 1510.290 2047.710 1511.470 ;
        RECT 2044.930 1331.890 2046.110 1333.070 ;
        RECT 2046.530 1331.890 2047.710 1333.070 ;
        RECT 2044.930 1330.290 2046.110 1331.470 ;
        RECT 2046.530 1330.290 2047.710 1331.470 ;
        RECT 2044.930 1151.890 2046.110 1153.070 ;
        RECT 2046.530 1151.890 2047.710 1153.070 ;
        RECT 2044.930 1150.290 2046.110 1151.470 ;
        RECT 2046.530 1150.290 2047.710 1151.470 ;
        RECT 2044.930 971.890 2046.110 973.070 ;
        RECT 2046.530 971.890 2047.710 973.070 ;
        RECT 2044.930 970.290 2046.110 971.470 ;
        RECT 2046.530 970.290 2047.710 971.470 ;
        RECT 2044.930 791.890 2046.110 793.070 ;
        RECT 2046.530 791.890 2047.710 793.070 ;
        RECT 2044.930 790.290 2046.110 791.470 ;
        RECT 2046.530 790.290 2047.710 791.470 ;
        RECT 2044.930 611.890 2046.110 613.070 ;
        RECT 2046.530 611.890 2047.710 613.070 ;
        RECT 2044.930 610.290 2046.110 611.470 ;
        RECT 2046.530 610.290 2047.710 611.470 ;
        RECT 2044.930 431.890 2046.110 433.070 ;
        RECT 2046.530 431.890 2047.710 433.070 ;
        RECT 2044.930 430.290 2046.110 431.470 ;
        RECT 2046.530 430.290 2047.710 431.470 ;
        RECT 2044.930 251.890 2046.110 253.070 ;
        RECT 2046.530 251.890 2047.710 253.070 ;
        RECT 2044.930 250.290 2046.110 251.470 ;
        RECT 2046.530 250.290 2047.710 251.470 ;
        RECT 2044.930 71.890 2046.110 73.070 ;
        RECT 2046.530 71.890 2047.710 73.070 ;
        RECT 2044.930 70.290 2046.110 71.470 ;
        RECT 2046.530 70.290 2047.710 71.470 ;
        RECT 2044.930 -31.710 2046.110 -30.530 ;
        RECT 2046.530 -31.710 2047.710 -30.530 ;
        RECT 2044.930 -33.310 2046.110 -32.130 ;
        RECT 2046.530 -33.310 2047.710 -32.130 ;
        RECT 2224.930 3551.810 2226.110 3552.990 ;
        RECT 2226.530 3551.810 2227.710 3552.990 ;
        RECT 2224.930 3550.210 2226.110 3551.390 ;
        RECT 2226.530 3550.210 2227.710 3551.390 ;
        RECT 2224.930 3491.890 2226.110 3493.070 ;
        RECT 2226.530 3491.890 2227.710 3493.070 ;
        RECT 2224.930 3490.290 2226.110 3491.470 ;
        RECT 2226.530 3490.290 2227.710 3491.470 ;
        RECT 2224.930 3311.890 2226.110 3313.070 ;
        RECT 2226.530 3311.890 2227.710 3313.070 ;
        RECT 2224.930 3310.290 2226.110 3311.470 ;
        RECT 2226.530 3310.290 2227.710 3311.470 ;
        RECT 2224.930 3131.890 2226.110 3133.070 ;
        RECT 2226.530 3131.890 2227.710 3133.070 ;
        RECT 2224.930 3130.290 2226.110 3131.470 ;
        RECT 2226.530 3130.290 2227.710 3131.470 ;
        RECT 2224.930 2951.890 2226.110 2953.070 ;
        RECT 2226.530 2951.890 2227.710 2953.070 ;
        RECT 2224.930 2950.290 2226.110 2951.470 ;
        RECT 2226.530 2950.290 2227.710 2951.470 ;
        RECT 2224.930 2771.890 2226.110 2773.070 ;
        RECT 2226.530 2771.890 2227.710 2773.070 ;
        RECT 2224.930 2770.290 2226.110 2771.470 ;
        RECT 2226.530 2770.290 2227.710 2771.470 ;
        RECT 2224.930 2591.890 2226.110 2593.070 ;
        RECT 2226.530 2591.890 2227.710 2593.070 ;
        RECT 2224.930 2590.290 2226.110 2591.470 ;
        RECT 2226.530 2590.290 2227.710 2591.470 ;
        RECT 2224.930 2411.890 2226.110 2413.070 ;
        RECT 2226.530 2411.890 2227.710 2413.070 ;
        RECT 2224.930 2410.290 2226.110 2411.470 ;
        RECT 2226.530 2410.290 2227.710 2411.470 ;
        RECT 2224.930 2231.890 2226.110 2233.070 ;
        RECT 2226.530 2231.890 2227.710 2233.070 ;
        RECT 2224.930 2230.290 2226.110 2231.470 ;
        RECT 2226.530 2230.290 2227.710 2231.470 ;
        RECT 2224.930 2051.890 2226.110 2053.070 ;
        RECT 2226.530 2051.890 2227.710 2053.070 ;
        RECT 2224.930 2050.290 2226.110 2051.470 ;
        RECT 2226.530 2050.290 2227.710 2051.470 ;
        RECT 2224.930 1871.890 2226.110 1873.070 ;
        RECT 2226.530 1871.890 2227.710 1873.070 ;
        RECT 2224.930 1870.290 2226.110 1871.470 ;
        RECT 2226.530 1870.290 2227.710 1871.470 ;
        RECT 2224.930 1691.890 2226.110 1693.070 ;
        RECT 2226.530 1691.890 2227.710 1693.070 ;
        RECT 2224.930 1690.290 2226.110 1691.470 ;
        RECT 2226.530 1690.290 2227.710 1691.470 ;
        RECT 2224.930 1511.890 2226.110 1513.070 ;
        RECT 2226.530 1511.890 2227.710 1513.070 ;
        RECT 2224.930 1510.290 2226.110 1511.470 ;
        RECT 2226.530 1510.290 2227.710 1511.470 ;
        RECT 2224.930 1331.890 2226.110 1333.070 ;
        RECT 2226.530 1331.890 2227.710 1333.070 ;
        RECT 2224.930 1330.290 2226.110 1331.470 ;
        RECT 2226.530 1330.290 2227.710 1331.470 ;
        RECT 2224.930 1151.890 2226.110 1153.070 ;
        RECT 2226.530 1151.890 2227.710 1153.070 ;
        RECT 2224.930 1150.290 2226.110 1151.470 ;
        RECT 2226.530 1150.290 2227.710 1151.470 ;
        RECT 2224.930 971.890 2226.110 973.070 ;
        RECT 2226.530 971.890 2227.710 973.070 ;
        RECT 2224.930 970.290 2226.110 971.470 ;
        RECT 2226.530 970.290 2227.710 971.470 ;
        RECT 2224.930 791.890 2226.110 793.070 ;
        RECT 2226.530 791.890 2227.710 793.070 ;
        RECT 2224.930 790.290 2226.110 791.470 ;
        RECT 2226.530 790.290 2227.710 791.470 ;
        RECT 2224.930 611.890 2226.110 613.070 ;
        RECT 2226.530 611.890 2227.710 613.070 ;
        RECT 2224.930 610.290 2226.110 611.470 ;
        RECT 2226.530 610.290 2227.710 611.470 ;
        RECT 2224.930 431.890 2226.110 433.070 ;
        RECT 2226.530 431.890 2227.710 433.070 ;
        RECT 2224.930 430.290 2226.110 431.470 ;
        RECT 2226.530 430.290 2227.710 431.470 ;
        RECT 2224.930 251.890 2226.110 253.070 ;
        RECT 2226.530 251.890 2227.710 253.070 ;
        RECT 2224.930 250.290 2226.110 251.470 ;
        RECT 2226.530 250.290 2227.710 251.470 ;
        RECT 2224.930 71.890 2226.110 73.070 ;
        RECT 2226.530 71.890 2227.710 73.070 ;
        RECT 2224.930 70.290 2226.110 71.470 ;
        RECT 2226.530 70.290 2227.710 71.470 ;
        RECT 2224.930 -31.710 2226.110 -30.530 ;
        RECT 2226.530 -31.710 2227.710 -30.530 ;
        RECT 2224.930 -33.310 2226.110 -32.130 ;
        RECT 2226.530 -33.310 2227.710 -32.130 ;
        RECT 2404.930 3551.810 2406.110 3552.990 ;
        RECT 2406.530 3551.810 2407.710 3552.990 ;
        RECT 2404.930 3550.210 2406.110 3551.390 ;
        RECT 2406.530 3550.210 2407.710 3551.390 ;
        RECT 2404.930 3491.890 2406.110 3493.070 ;
        RECT 2406.530 3491.890 2407.710 3493.070 ;
        RECT 2404.930 3490.290 2406.110 3491.470 ;
        RECT 2406.530 3490.290 2407.710 3491.470 ;
        RECT 2404.930 3311.890 2406.110 3313.070 ;
        RECT 2406.530 3311.890 2407.710 3313.070 ;
        RECT 2404.930 3310.290 2406.110 3311.470 ;
        RECT 2406.530 3310.290 2407.710 3311.470 ;
        RECT 2404.930 3131.890 2406.110 3133.070 ;
        RECT 2406.530 3131.890 2407.710 3133.070 ;
        RECT 2404.930 3130.290 2406.110 3131.470 ;
        RECT 2406.530 3130.290 2407.710 3131.470 ;
        RECT 2404.930 2951.890 2406.110 2953.070 ;
        RECT 2406.530 2951.890 2407.710 2953.070 ;
        RECT 2404.930 2950.290 2406.110 2951.470 ;
        RECT 2406.530 2950.290 2407.710 2951.470 ;
        RECT 2404.930 2771.890 2406.110 2773.070 ;
        RECT 2406.530 2771.890 2407.710 2773.070 ;
        RECT 2404.930 2770.290 2406.110 2771.470 ;
        RECT 2406.530 2770.290 2407.710 2771.470 ;
        RECT 2404.930 2591.890 2406.110 2593.070 ;
        RECT 2406.530 2591.890 2407.710 2593.070 ;
        RECT 2404.930 2590.290 2406.110 2591.470 ;
        RECT 2406.530 2590.290 2407.710 2591.470 ;
        RECT 2404.930 2411.890 2406.110 2413.070 ;
        RECT 2406.530 2411.890 2407.710 2413.070 ;
        RECT 2404.930 2410.290 2406.110 2411.470 ;
        RECT 2406.530 2410.290 2407.710 2411.470 ;
        RECT 2404.930 2231.890 2406.110 2233.070 ;
        RECT 2406.530 2231.890 2407.710 2233.070 ;
        RECT 2404.930 2230.290 2406.110 2231.470 ;
        RECT 2406.530 2230.290 2407.710 2231.470 ;
        RECT 2404.930 2051.890 2406.110 2053.070 ;
        RECT 2406.530 2051.890 2407.710 2053.070 ;
        RECT 2404.930 2050.290 2406.110 2051.470 ;
        RECT 2406.530 2050.290 2407.710 2051.470 ;
        RECT 2404.930 1871.890 2406.110 1873.070 ;
        RECT 2406.530 1871.890 2407.710 1873.070 ;
        RECT 2404.930 1870.290 2406.110 1871.470 ;
        RECT 2406.530 1870.290 2407.710 1871.470 ;
        RECT 2404.930 1691.890 2406.110 1693.070 ;
        RECT 2406.530 1691.890 2407.710 1693.070 ;
        RECT 2404.930 1690.290 2406.110 1691.470 ;
        RECT 2406.530 1690.290 2407.710 1691.470 ;
        RECT 2404.930 1511.890 2406.110 1513.070 ;
        RECT 2406.530 1511.890 2407.710 1513.070 ;
        RECT 2404.930 1510.290 2406.110 1511.470 ;
        RECT 2406.530 1510.290 2407.710 1511.470 ;
        RECT 2404.930 1331.890 2406.110 1333.070 ;
        RECT 2406.530 1331.890 2407.710 1333.070 ;
        RECT 2404.930 1330.290 2406.110 1331.470 ;
        RECT 2406.530 1330.290 2407.710 1331.470 ;
        RECT 2404.930 1151.890 2406.110 1153.070 ;
        RECT 2406.530 1151.890 2407.710 1153.070 ;
        RECT 2404.930 1150.290 2406.110 1151.470 ;
        RECT 2406.530 1150.290 2407.710 1151.470 ;
        RECT 2404.930 971.890 2406.110 973.070 ;
        RECT 2406.530 971.890 2407.710 973.070 ;
        RECT 2404.930 970.290 2406.110 971.470 ;
        RECT 2406.530 970.290 2407.710 971.470 ;
        RECT 2404.930 791.890 2406.110 793.070 ;
        RECT 2406.530 791.890 2407.710 793.070 ;
        RECT 2404.930 790.290 2406.110 791.470 ;
        RECT 2406.530 790.290 2407.710 791.470 ;
        RECT 2404.930 611.890 2406.110 613.070 ;
        RECT 2406.530 611.890 2407.710 613.070 ;
        RECT 2404.930 610.290 2406.110 611.470 ;
        RECT 2406.530 610.290 2407.710 611.470 ;
        RECT 2404.930 431.890 2406.110 433.070 ;
        RECT 2406.530 431.890 2407.710 433.070 ;
        RECT 2404.930 430.290 2406.110 431.470 ;
        RECT 2406.530 430.290 2407.710 431.470 ;
        RECT 2404.930 251.890 2406.110 253.070 ;
        RECT 2406.530 251.890 2407.710 253.070 ;
        RECT 2404.930 250.290 2406.110 251.470 ;
        RECT 2406.530 250.290 2407.710 251.470 ;
        RECT 2404.930 71.890 2406.110 73.070 ;
        RECT 2406.530 71.890 2407.710 73.070 ;
        RECT 2404.930 70.290 2406.110 71.470 ;
        RECT 2406.530 70.290 2407.710 71.470 ;
        RECT 2404.930 -31.710 2406.110 -30.530 ;
        RECT 2406.530 -31.710 2407.710 -30.530 ;
        RECT 2404.930 -33.310 2406.110 -32.130 ;
        RECT 2406.530 -33.310 2407.710 -32.130 ;
        RECT 2584.930 3551.810 2586.110 3552.990 ;
        RECT 2586.530 3551.810 2587.710 3552.990 ;
        RECT 2584.930 3550.210 2586.110 3551.390 ;
        RECT 2586.530 3550.210 2587.710 3551.390 ;
        RECT 2584.930 3491.890 2586.110 3493.070 ;
        RECT 2586.530 3491.890 2587.710 3493.070 ;
        RECT 2584.930 3490.290 2586.110 3491.470 ;
        RECT 2586.530 3490.290 2587.710 3491.470 ;
        RECT 2584.930 3311.890 2586.110 3313.070 ;
        RECT 2586.530 3311.890 2587.710 3313.070 ;
        RECT 2584.930 3310.290 2586.110 3311.470 ;
        RECT 2586.530 3310.290 2587.710 3311.470 ;
        RECT 2584.930 3131.890 2586.110 3133.070 ;
        RECT 2586.530 3131.890 2587.710 3133.070 ;
        RECT 2584.930 3130.290 2586.110 3131.470 ;
        RECT 2586.530 3130.290 2587.710 3131.470 ;
        RECT 2584.930 2951.890 2586.110 2953.070 ;
        RECT 2586.530 2951.890 2587.710 2953.070 ;
        RECT 2584.930 2950.290 2586.110 2951.470 ;
        RECT 2586.530 2950.290 2587.710 2951.470 ;
        RECT 2584.930 2771.890 2586.110 2773.070 ;
        RECT 2586.530 2771.890 2587.710 2773.070 ;
        RECT 2584.930 2770.290 2586.110 2771.470 ;
        RECT 2586.530 2770.290 2587.710 2771.470 ;
        RECT 2584.930 2591.890 2586.110 2593.070 ;
        RECT 2586.530 2591.890 2587.710 2593.070 ;
        RECT 2584.930 2590.290 2586.110 2591.470 ;
        RECT 2586.530 2590.290 2587.710 2591.470 ;
        RECT 2584.930 2411.890 2586.110 2413.070 ;
        RECT 2586.530 2411.890 2587.710 2413.070 ;
        RECT 2584.930 2410.290 2586.110 2411.470 ;
        RECT 2586.530 2410.290 2587.710 2411.470 ;
        RECT 2584.930 2231.890 2586.110 2233.070 ;
        RECT 2586.530 2231.890 2587.710 2233.070 ;
        RECT 2584.930 2230.290 2586.110 2231.470 ;
        RECT 2586.530 2230.290 2587.710 2231.470 ;
        RECT 2584.930 2051.890 2586.110 2053.070 ;
        RECT 2586.530 2051.890 2587.710 2053.070 ;
        RECT 2584.930 2050.290 2586.110 2051.470 ;
        RECT 2586.530 2050.290 2587.710 2051.470 ;
        RECT 2584.930 1871.890 2586.110 1873.070 ;
        RECT 2586.530 1871.890 2587.710 1873.070 ;
        RECT 2584.930 1870.290 2586.110 1871.470 ;
        RECT 2586.530 1870.290 2587.710 1871.470 ;
        RECT 2584.930 1691.890 2586.110 1693.070 ;
        RECT 2586.530 1691.890 2587.710 1693.070 ;
        RECT 2584.930 1690.290 2586.110 1691.470 ;
        RECT 2586.530 1690.290 2587.710 1691.470 ;
        RECT 2584.930 1511.890 2586.110 1513.070 ;
        RECT 2586.530 1511.890 2587.710 1513.070 ;
        RECT 2584.930 1510.290 2586.110 1511.470 ;
        RECT 2586.530 1510.290 2587.710 1511.470 ;
        RECT 2584.930 1331.890 2586.110 1333.070 ;
        RECT 2586.530 1331.890 2587.710 1333.070 ;
        RECT 2584.930 1330.290 2586.110 1331.470 ;
        RECT 2586.530 1330.290 2587.710 1331.470 ;
        RECT 2584.930 1151.890 2586.110 1153.070 ;
        RECT 2586.530 1151.890 2587.710 1153.070 ;
        RECT 2584.930 1150.290 2586.110 1151.470 ;
        RECT 2586.530 1150.290 2587.710 1151.470 ;
        RECT 2584.930 971.890 2586.110 973.070 ;
        RECT 2586.530 971.890 2587.710 973.070 ;
        RECT 2584.930 970.290 2586.110 971.470 ;
        RECT 2586.530 970.290 2587.710 971.470 ;
        RECT 2584.930 791.890 2586.110 793.070 ;
        RECT 2586.530 791.890 2587.710 793.070 ;
        RECT 2584.930 790.290 2586.110 791.470 ;
        RECT 2586.530 790.290 2587.710 791.470 ;
        RECT 2584.930 611.890 2586.110 613.070 ;
        RECT 2586.530 611.890 2587.710 613.070 ;
        RECT 2584.930 610.290 2586.110 611.470 ;
        RECT 2586.530 610.290 2587.710 611.470 ;
        RECT 2584.930 431.890 2586.110 433.070 ;
        RECT 2586.530 431.890 2587.710 433.070 ;
        RECT 2584.930 430.290 2586.110 431.470 ;
        RECT 2586.530 430.290 2587.710 431.470 ;
        RECT 2584.930 251.890 2586.110 253.070 ;
        RECT 2586.530 251.890 2587.710 253.070 ;
        RECT 2584.930 250.290 2586.110 251.470 ;
        RECT 2586.530 250.290 2587.710 251.470 ;
        RECT 2584.930 71.890 2586.110 73.070 ;
        RECT 2586.530 71.890 2587.710 73.070 ;
        RECT 2584.930 70.290 2586.110 71.470 ;
        RECT 2586.530 70.290 2587.710 71.470 ;
        RECT 2584.930 -31.710 2586.110 -30.530 ;
        RECT 2586.530 -31.710 2587.710 -30.530 ;
        RECT 2584.930 -33.310 2586.110 -32.130 ;
        RECT 2586.530 -33.310 2587.710 -32.130 ;
        RECT 2764.930 3551.810 2766.110 3552.990 ;
        RECT 2766.530 3551.810 2767.710 3552.990 ;
        RECT 2764.930 3550.210 2766.110 3551.390 ;
        RECT 2766.530 3550.210 2767.710 3551.390 ;
        RECT 2764.930 3491.890 2766.110 3493.070 ;
        RECT 2766.530 3491.890 2767.710 3493.070 ;
        RECT 2764.930 3490.290 2766.110 3491.470 ;
        RECT 2766.530 3490.290 2767.710 3491.470 ;
        RECT 2764.930 3311.890 2766.110 3313.070 ;
        RECT 2766.530 3311.890 2767.710 3313.070 ;
        RECT 2764.930 3310.290 2766.110 3311.470 ;
        RECT 2766.530 3310.290 2767.710 3311.470 ;
        RECT 2764.930 3131.890 2766.110 3133.070 ;
        RECT 2766.530 3131.890 2767.710 3133.070 ;
        RECT 2764.930 3130.290 2766.110 3131.470 ;
        RECT 2766.530 3130.290 2767.710 3131.470 ;
        RECT 2764.930 2951.890 2766.110 2953.070 ;
        RECT 2766.530 2951.890 2767.710 2953.070 ;
        RECT 2764.930 2950.290 2766.110 2951.470 ;
        RECT 2766.530 2950.290 2767.710 2951.470 ;
        RECT 2764.930 2771.890 2766.110 2773.070 ;
        RECT 2766.530 2771.890 2767.710 2773.070 ;
        RECT 2764.930 2770.290 2766.110 2771.470 ;
        RECT 2766.530 2770.290 2767.710 2771.470 ;
        RECT 2764.930 2591.890 2766.110 2593.070 ;
        RECT 2766.530 2591.890 2767.710 2593.070 ;
        RECT 2764.930 2590.290 2766.110 2591.470 ;
        RECT 2766.530 2590.290 2767.710 2591.470 ;
        RECT 2764.930 2411.890 2766.110 2413.070 ;
        RECT 2766.530 2411.890 2767.710 2413.070 ;
        RECT 2764.930 2410.290 2766.110 2411.470 ;
        RECT 2766.530 2410.290 2767.710 2411.470 ;
        RECT 2764.930 2231.890 2766.110 2233.070 ;
        RECT 2766.530 2231.890 2767.710 2233.070 ;
        RECT 2764.930 2230.290 2766.110 2231.470 ;
        RECT 2766.530 2230.290 2767.710 2231.470 ;
        RECT 2764.930 2051.890 2766.110 2053.070 ;
        RECT 2766.530 2051.890 2767.710 2053.070 ;
        RECT 2764.930 2050.290 2766.110 2051.470 ;
        RECT 2766.530 2050.290 2767.710 2051.470 ;
        RECT 2764.930 1871.890 2766.110 1873.070 ;
        RECT 2766.530 1871.890 2767.710 1873.070 ;
        RECT 2764.930 1870.290 2766.110 1871.470 ;
        RECT 2766.530 1870.290 2767.710 1871.470 ;
        RECT 2764.930 1691.890 2766.110 1693.070 ;
        RECT 2766.530 1691.890 2767.710 1693.070 ;
        RECT 2764.930 1690.290 2766.110 1691.470 ;
        RECT 2766.530 1690.290 2767.710 1691.470 ;
        RECT 2764.930 1511.890 2766.110 1513.070 ;
        RECT 2766.530 1511.890 2767.710 1513.070 ;
        RECT 2764.930 1510.290 2766.110 1511.470 ;
        RECT 2766.530 1510.290 2767.710 1511.470 ;
        RECT 2764.930 1331.890 2766.110 1333.070 ;
        RECT 2766.530 1331.890 2767.710 1333.070 ;
        RECT 2764.930 1330.290 2766.110 1331.470 ;
        RECT 2766.530 1330.290 2767.710 1331.470 ;
        RECT 2764.930 1151.890 2766.110 1153.070 ;
        RECT 2766.530 1151.890 2767.710 1153.070 ;
        RECT 2764.930 1150.290 2766.110 1151.470 ;
        RECT 2766.530 1150.290 2767.710 1151.470 ;
        RECT 2764.930 971.890 2766.110 973.070 ;
        RECT 2766.530 971.890 2767.710 973.070 ;
        RECT 2764.930 970.290 2766.110 971.470 ;
        RECT 2766.530 970.290 2767.710 971.470 ;
        RECT 2764.930 791.890 2766.110 793.070 ;
        RECT 2766.530 791.890 2767.710 793.070 ;
        RECT 2764.930 790.290 2766.110 791.470 ;
        RECT 2766.530 790.290 2767.710 791.470 ;
        RECT 2764.930 611.890 2766.110 613.070 ;
        RECT 2766.530 611.890 2767.710 613.070 ;
        RECT 2764.930 610.290 2766.110 611.470 ;
        RECT 2766.530 610.290 2767.710 611.470 ;
        RECT 2764.930 431.890 2766.110 433.070 ;
        RECT 2766.530 431.890 2767.710 433.070 ;
        RECT 2764.930 430.290 2766.110 431.470 ;
        RECT 2766.530 430.290 2767.710 431.470 ;
        RECT 2764.930 251.890 2766.110 253.070 ;
        RECT 2766.530 251.890 2767.710 253.070 ;
        RECT 2764.930 250.290 2766.110 251.470 ;
        RECT 2766.530 250.290 2767.710 251.470 ;
        RECT 2764.930 71.890 2766.110 73.070 ;
        RECT 2766.530 71.890 2767.710 73.070 ;
        RECT 2764.930 70.290 2766.110 71.470 ;
        RECT 2766.530 70.290 2767.710 71.470 ;
        RECT 2764.930 -31.710 2766.110 -30.530 ;
        RECT 2766.530 -31.710 2767.710 -30.530 ;
        RECT 2764.930 -33.310 2766.110 -32.130 ;
        RECT 2766.530 -33.310 2767.710 -32.130 ;
        RECT 2955.510 3551.810 2956.690 3552.990 ;
        RECT 2957.110 3551.810 2958.290 3552.990 ;
        RECT 2955.510 3550.210 2956.690 3551.390 ;
        RECT 2957.110 3550.210 2958.290 3551.390 ;
        RECT 2955.510 3491.890 2956.690 3493.070 ;
        RECT 2957.110 3491.890 2958.290 3493.070 ;
        RECT 2955.510 3490.290 2956.690 3491.470 ;
        RECT 2957.110 3490.290 2958.290 3491.470 ;
        RECT 2955.510 3311.890 2956.690 3313.070 ;
        RECT 2957.110 3311.890 2958.290 3313.070 ;
        RECT 2955.510 3310.290 2956.690 3311.470 ;
        RECT 2957.110 3310.290 2958.290 3311.470 ;
        RECT 2955.510 3131.890 2956.690 3133.070 ;
        RECT 2957.110 3131.890 2958.290 3133.070 ;
        RECT 2955.510 3130.290 2956.690 3131.470 ;
        RECT 2957.110 3130.290 2958.290 3131.470 ;
        RECT 2955.510 2951.890 2956.690 2953.070 ;
        RECT 2957.110 2951.890 2958.290 2953.070 ;
        RECT 2955.510 2950.290 2956.690 2951.470 ;
        RECT 2957.110 2950.290 2958.290 2951.470 ;
        RECT 2955.510 2771.890 2956.690 2773.070 ;
        RECT 2957.110 2771.890 2958.290 2773.070 ;
        RECT 2955.510 2770.290 2956.690 2771.470 ;
        RECT 2957.110 2770.290 2958.290 2771.470 ;
        RECT 2955.510 2591.890 2956.690 2593.070 ;
        RECT 2957.110 2591.890 2958.290 2593.070 ;
        RECT 2955.510 2590.290 2956.690 2591.470 ;
        RECT 2957.110 2590.290 2958.290 2591.470 ;
        RECT 2955.510 2411.890 2956.690 2413.070 ;
        RECT 2957.110 2411.890 2958.290 2413.070 ;
        RECT 2955.510 2410.290 2956.690 2411.470 ;
        RECT 2957.110 2410.290 2958.290 2411.470 ;
        RECT 2955.510 2231.890 2956.690 2233.070 ;
        RECT 2957.110 2231.890 2958.290 2233.070 ;
        RECT 2955.510 2230.290 2956.690 2231.470 ;
        RECT 2957.110 2230.290 2958.290 2231.470 ;
        RECT 2955.510 2051.890 2956.690 2053.070 ;
        RECT 2957.110 2051.890 2958.290 2053.070 ;
        RECT 2955.510 2050.290 2956.690 2051.470 ;
        RECT 2957.110 2050.290 2958.290 2051.470 ;
        RECT 2955.510 1871.890 2956.690 1873.070 ;
        RECT 2957.110 1871.890 2958.290 1873.070 ;
        RECT 2955.510 1870.290 2956.690 1871.470 ;
        RECT 2957.110 1870.290 2958.290 1871.470 ;
        RECT 2955.510 1691.890 2956.690 1693.070 ;
        RECT 2957.110 1691.890 2958.290 1693.070 ;
        RECT 2955.510 1690.290 2956.690 1691.470 ;
        RECT 2957.110 1690.290 2958.290 1691.470 ;
        RECT 2955.510 1511.890 2956.690 1513.070 ;
        RECT 2957.110 1511.890 2958.290 1513.070 ;
        RECT 2955.510 1510.290 2956.690 1511.470 ;
        RECT 2957.110 1510.290 2958.290 1511.470 ;
        RECT 2955.510 1331.890 2956.690 1333.070 ;
        RECT 2957.110 1331.890 2958.290 1333.070 ;
        RECT 2955.510 1330.290 2956.690 1331.470 ;
        RECT 2957.110 1330.290 2958.290 1331.470 ;
        RECT 2955.510 1151.890 2956.690 1153.070 ;
        RECT 2957.110 1151.890 2958.290 1153.070 ;
        RECT 2955.510 1150.290 2956.690 1151.470 ;
        RECT 2957.110 1150.290 2958.290 1151.470 ;
        RECT 2955.510 971.890 2956.690 973.070 ;
        RECT 2957.110 971.890 2958.290 973.070 ;
        RECT 2955.510 970.290 2956.690 971.470 ;
        RECT 2957.110 970.290 2958.290 971.470 ;
        RECT 2955.510 791.890 2956.690 793.070 ;
        RECT 2957.110 791.890 2958.290 793.070 ;
        RECT 2955.510 790.290 2956.690 791.470 ;
        RECT 2957.110 790.290 2958.290 791.470 ;
        RECT 2955.510 611.890 2956.690 613.070 ;
        RECT 2957.110 611.890 2958.290 613.070 ;
        RECT 2955.510 610.290 2956.690 611.470 ;
        RECT 2957.110 610.290 2958.290 611.470 ;
        RECT 2955.510 431.890 2956.690 433.070 ;
        RECT 2957.110 431.890 2958.290 433.070 ;
        RECT 2955.510 430.290 2956.690 431.470 ;
        RECT 2957.110 430.290 2958.290 431.470 ;
        RECT 2955.510 251.890 2956.690 253.070 ;
        RECT 2957.110 251.890 2958.290 253.070 ;
        RECT 2955.510 250.290 2956.690 251.470 ;
        RECT 2957.110 250.290 2958.290 251.470 ;
        RECT 2955.510 71.890 2956.690 73.070 ;
        RECT 2957.110 71.890 2958.290 73.070 ;
        RECT 2955.510 70.290 2956.690 71.470 ;
        RECT 2957.110 70.290 2958.290 71.470 ;
        RECT 2955.510 -31.710 2956.690 -30.530 ;
        RECT 2957.110 -31.710 2958.290 -30.530 ;
        RECT 2955.510 -33.310 2956.690 -32.130 ;
        RECT 2957.110 -33.310 2958.290 -32.130 ;
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
        RECT -43.630 970.130 2963.250 973.230 ;
        RECT -43.630 790.130 2963.250 793.230 ;
        RECT -43.630 610.130 2963.250 613.230 ;
        RECT -43.630 430.130 2963.250 433.230 ;
        RECT -43.630 250.130 2963.250 253.230 ;
        RECT -43.630 70.130 2963.250 73.230 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
        RECT 316.170 1010.000 319.270 3548.350 ;
        RECT 496.170 1010.000 499.270 3548.350 ;
        RECT 676.170 1010.000 679.270 3548.350 ;
        RECT 856.170 1010.000 859.270 3548.350 ;
        RECT 1036.170 1010.000 1039.270 3548.350 ;
        RECT 316.170 -28.670 319.270 390.000 ;
        RECT 496.170 -28.670 499.270 390.000 ;
        RECT 676.170 -28.670 679.270 390.000 ;
        RECT 856.170 -28.670 859.270 390.000 ;
        RECT 1036.170 -28.670 1039.270 390.000 ;
        RECT 1216.170 -28.670 1219.270 3548.350 ;
        RECT 1396.170 -28.670 1399.270 3548.350 ;
        RECT 1576.170 -28.670 1579.270 3548.350 ;
        RECT 1756.170 -28.670 1759.270 3548.350 ;
        RECT 1936.170 -28.670 1939.270 3548.350 ;
        RECT 2116.170 -28.670 2119.270 3548.350 ;
        RECT 2296.170 -28.670 2299.270 3548.350 ;
        RECT 2476.170 -28.670 2479.270 3548.350 ;
        RECT 2656.170 -28.670 2659.270 3548.350 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
      LAYER via4 ;
        RECT -33.870 3547.010 -32.690 3548.190 ;
        RECT -32.270 3547.010 -31.090 3548.190 ;
        RECT -33.870 3545.410 -32.690 3546.590 ;
        RECT -32.270 3545.410 -31.090 3546.590 ;
        RECT -33.870 3383.290 -32.690 3384.470 ;
        RECT -32.270 3383.290 -31.090 3384.470 ;
        RECT -33.870 3381.690 -32.690 3382.870 ;
        RECT -32.270 3381.690 -31.090 3382.870 ;
        RECT -33.870 3203.290 -32.690 3204.470 ;
        RECT -32.270 3203.290 -31.090 3204.470 ;
        RECT -33.870 3201.690 -32.690 3202.870 ;
        RECT -32.270 3201.690 -31.090 3202.870 ;
        RECT -33.870 3023.290 -32.690 3024.470 ;
        RECT -32.270 3023.290 -31.090 3024.470 ;
        RECT -33.870 3021.690 -32.690 3022.870 ;
        RECT -32.270 3021.690 -31.090 3022.870 ;
        RECT -33.870 2843.290 -32.690 2844.470 ;
        RECT -32.270 2843.290 -31.090 2844.470 ;
        RECT -33.870 2841.690 -32.690 2842.870 ;
        RECT -32.270 2841.690 -31.090 2842.870 ;
        RECT -33.870 2663.290 -32.690 2664.470 ;
        RECT -32.270 2663.290 -31.090 2664.470 ;
        RECT -33.870 2661.690 -32.690 2662.870 ;
        RECT -32.270 2661.690 -31.090 2662.870 ;
        RECT -33.870 2483.290 -32.690 2484.470 ;
        RECT -32.270 2483.290 -31.090 2484.470 ;
        RECT -33.870 2481.690 -32.690 2482.870 ;
        RECT -32.270 2481.690 -31.090 2482.870 ;
        RECT -33.870 2303.290 -32.690 2304.470 ;
        RECT -32.270 2303.290 -31.090 2304.470 ;
        RECT -33.870 2301.690 -32.690 2302.870 ;
        RECT -32.270 2301.690 -31.090 2302.870 ;
        RECT -33.870 2123.290 -32.690 2124.470 ;
        RECT -32.270 2123.290 -31.090 2124.470 ;
        RECT -33.870 2121.690 -32.690 2122.870 ;
        RECT -32.270 2121.690 -31.090 2122.870 ;
        RECT -33.870 1943.290 -32.690 1944.470 ;
        RECT -32.270 1943.290 -31.090 1944.470 ;
        RECT -33.870 1941.690 -32.690 1942.870 ;
        RECT -32.270 1941.690 -31.090 1942.870 ;
        RECT -33.870 1763.290 -32.690 1764.470 ;
        RECT -32.270 1763.290 -31.090 1764.470 ;
        RECT -33.870 1761.690 -32.690 1762.870 ;
        RECT -32.270 1761.690 -31.090 1762.870 ;
        RECT -33.870 1583.290 -32.690 1584.470 ;
        RECT -32.270 1583.290 -31.090 1584.470 ;
        RECT -33.870 1581.690 -32.690 1582.870 ;
        RECT -32.270 1581.690 -31.090 1582.870 ;
        RECT -33.870 1403.290 -32.690 1404.470 ;
        RECT -32.270 1403.290 -31.090 1404.470 ;
        RECT -33.870 1401.690 -32.690 1402.870 ;
        RECT -32.270 1401.690 -31.090 1402.870 ;
        RECT -33.870 1223.290 -32.690 1224.470 ;
        RECT -32.270 1223.290 -31.090 1224.470 ;
        RECT -33.870 1221.690 -32.690 1222.870 ;
        RECT -32.270 1221.690 -31.090 1222.870 ;
        RECT -33.870 1043.290 -32.690 1044.470 ;
        RECT -32.270 1043.290 -31.090 1044.470 ;
        RECT -33.870 1041.690 -32.690 1042.870 ;
        RECT -32.270 1041.690 -31.090 1042.870 ;
        RECT -33.870 863.290 -32.690 864.470 ;
        RECT -32.270 863.290 -31.090 864.470 ;
        RECT -33.870 861.690 -32.690 862.870 ;
        RECT -32.270 861.690 -31.090 862.870 ;
        RECT -33.870 683.290 -32.690 684.470 ;
        RECT -32.270 683.290 -31.090 684.470 ;
        RECT -33.870 681.690 -32.690 682.870 ;
        RECT -32.270 681.690 -31.090 682.870 ;
        RECT -33.870 503.290 -32.690 504.470 ;
        RECT -32.270 503.290 -31.090 504.470 ;
        RECT -33.870 501.690 -32.690 502.870 ;
        RECT -32.270 501.690 -31.090 502.870 ;
        RECT -33.870 323.290 -32.690 324.470 ;
        RECT -32.270 323.290 -31.090 324.470 ;
        RECT -33.870 321.690 -32.690 322.870 ;
        RECT -32.270 321.690 -31.090 322.870 ;
        RECT -33.870 143.290 -32.690 144.470 ;
        RECT -32.270 143.290 -31.090 144.470 ;
        RECT -33.870 141.690 -32.690 142.870 ;
        RECT -32.270 141.690 -31.090 142.870 ;
        RECT -33.870 -26.910 -32.690 -25.730 ;
        RECT -32.270 -26.910 -31.090 -25.730 ;
        RECT -33.870 -28.510 -32.690 -27.330 ;
        RECT -32.270 -28.510 -31.090 -27.330 ;
        RECT 136.330 3547.010 137.510 3548.190 ;
        RECT 137.930 3547.010 139.110 3548.190 ;
        RECT 136.330 3545.410 137.510 3546.590 ;
        RECT 137.930 3545.410 139.110 3546.590 ;
        RECT 136.330 3383.290 137.510 3384.470 ;
        RECT 137.930 3383.290 139.110 3384.470 ;
        RECT 136.330 3381.690 137.510 3382.870 ;
        RECT 137.930 3381.690 139.110 3382.870 ;
        RECT 136.330 3203.290 137.510 3204.470 ;
        RECT 137.930 3203.290 139.110 3204.470 ;
        RECT 136.330 3201.690 137.510 3202.870 ;
        RECT 137.930 3201.690 139.110 3202.870 ;
        RECT 136.330 3023.290 137.510 3024.470 ;
        RECT 137.930 3023.290 139.110 3024.470 ;
        RECT 136.330 3021.690 137.510 3022.870 ;
        RECT 137.930 3021.690 139.110 3022.870 ;
        RECT 136.330 2843.290 137.510 2844.470 ;
        RECT 137.930 2843.290 139.110 2844.470 ;
        RECT 136.330 2841.690 137.510 2842.870 ;
        RECT 137.930 2841.690 139.110 2842.870 ;
        RECT 136.330 2663.290 137.510 2664.470 ;
        RECT 137.930 2663.290 139.110 2664.470 ;
        RECT 136.330 2661.690 137.510 2662.870 ;
        RECT 137.930 2661.690 139.110 2662.870 ;
        RECT 136.330 2483.290 137.510 2484.470 ;
        RECT 137.930 2483.290 139.110 2484.470 ;
        RECT 136.330 2481.690 137.510 2482.870 ;
        RECT 137.930 2481.690 139.110 2482.870 ;
        RECT 136.330 2303.290 137.510 2304.470 ;
        RECT 137.930 2303.290 139.110 2304.470 ;
        RECT 136.330 2301.690 137.510 2302.870 ;
        RECT 137.930 2301.690 139.110 2302.870 ;
        RECT 136.330 2123.290 137.510 2124.470 ;
        RECT 137.930 2123.290 139.110 2124.470 ;
        RECT 136.330 2121.690 137.510 2122.870 ;
        RECT 137.930 2121.690 139.110 2122.870 ;
        RECT 136.330 1943.290 137.510 1944.470 ;
        RECT 137.930 1943.290 139.110 1944.470 ;
        RECT 136.330 1941.690 137.510 1942.870 ;
        RECT 137.930 1941.690 139.110 1942.870 ;
        RECT 136.330 1763.290 137.510 1764.470 ;
        RECT 137.930 1763.290 139.110 1764.470 ;
        RECT 136.330 1761.690 137.510 1762.870 ;
        RECT 137.930 1761.690 139.110 1762.870 ;
        RECT 136.330 1583.290 137.510 1584.470 ;
        RECT 137.930 1583.290 139.110 1584.470 ;
        RECT 136.330 1581.690 137.510 1582.870 ;
        RECT 137.930 1581.690 139.110 1582.870 ;
        RECT 136.330 1403.290 137.510 1404.470 ;
        RECT 137.930 1403.290 139.110 1404.470 ;
        RECT 136.330 1401.690 137.510 1402.870 ;
        RECT 137.930 1401.690 139.110 1402.870 ;
        RECT 136.330 1223.290 137.510 1224.470 ;
        RECT 137.930 1223.290 139.110 1224.470 ;
        RECT 136.330 1221.690 137.510 1222.870 ;
        RECT 137.930 1221.690 139.110 1222.870 ;
        RECT 136.330 1043.290 137.510 1044.470 ;
        RECT 137.930 1043.290 139.110 1044.470 ;
        RECT 136.330 1041.690 137.510 1042.870 ;
        RECT 137.930 1041.690 139.110 1042.870 ;
        RECT 316.330 3547.010 317.510 3548.190 ;
        RECT 317.930 3547.010 319.110 3548.190 ;
        RECT 316.330 3545.410 317.510 3546.590 ;
        RECT 317.930 3545.410 319.110 3546.590 ;
        RECT 316.330 3383.290 317.510 3384.470 ;
        RECT 317.930 3383.290 319.110 3384.470 ;
        RECT 316.330 3381.690 317.510 3382.870 ;
        RECT 317.930 3381.690 319.110 3382.870 ;
        RECT 316.330 3203.290 317.510 3204.470 ;
        RECT 317.930 3203.290 319.110 3204.470 ;
        RECT 316.330 3201.690 317.510 3202.870 ;
        RECT 317.930 3201.690 319.110 3202.870 ;
        RECT 316.330 3023.290 317.510 3024.470 ;
        RECT 317.930 3023.290 319.110 3024.470 ;
        RECT 316.330 3021.690 317.510 3022.870 ;
        RECT 317.930 3021.690 319.110 3022.870 ;
        RECT 316.330 2843.290 317.510 2844.470 ;
        RECT 317.930 2843.290 319.110 2844.470 ;
        RECT 316.330 2841.690 317.510 2842.870 ;
        RECT 317.930 2841.690 319.110 2842.870 ;
        RECT 316.330 2663.290 317.510 2664.470 ;
        RECT 317.930 2663.290 319.110 2664.470 ;
        RECT 316.330 2661.690 317.510 2662.870 ;
        RECT 317.930 2661.690 319.110 2662.870 ;
        RECT 316.330 2483.290 317.510 2484.470 ;
        RECT 317.930 2483.290 319.110 2484.470 ;
        RECT 316.330 2481.690 317.510 2482.870 ;
        RECT 317.930 2481.690 319.110 2482.870 ;
        RECT 316.330 2303.290 317.510 2304.470 ;
        RECT 317.930 2303.290 319.110 2304.470 ;
        RECT 316.330 2301.690 317.510 2302.870 ;
        RECT 317.930 2301.690 319.110 2302.870 ;
        RECT 316.330 2123.290 317.510 2124.470 ;
        RECT 317.930 2123.290 319.110 2124.470 ;
        RECT 316.330 2121.690 317.510 2122.870 ;
        RECT 317.930 2121.690 319.110 2122.870 ;
        RECT 316.330 1943.290 317.510 1944.470 ;
        RECT 317.930 1943.290 319.110 1944.470 ;
        RECT 316.330 1941.690 317.510 1942.870 ;
        RECT 317.930 1941.690 319.110 1942.870 ;
        RECT 316.330 1763.290 317.510 1764.470 ;
        RECT 317.930 1763.290 319.110 1764.470 ;
        RECT 316.330 1761.690 317.510 1762.870 ;
        RECT 317.930 1761.690 319.110 1762.870 ;
        RECT 316.330 1583.290 317.510 1584.470 ;
        RECT 317.930 1583.290 319.110 1584.470 ;
        RECT 316.330 1581.690 317.510 1582.870 ;
        RECT 317.930 1581.690 319.110 1582.870 ;
        RECT 316.330 1403.290 317.510 1404.470 ;
        RECT 317.930 1403.290 319.110 1404.470 ;
        RECT 316.330 1401.690 317.510 1402.870 ;
        RECT 317.930 1401.690 319.110 1402.870 ;
        RECT 316.330 1223.290 317.510 1224.470 ;
        RECT 317.930 1223.290 319.110 1224.470 ;
        RECT 316.330 1221.690 317.510 1222.870 ;
        RECT 317.930 1221.690 319.110 1222.870 ;
        RECT 316.330 1043.290 317.510 1044.470 ;
        RECT 317.930 1043.290 319.110 1044.470 ;
        RECT 316.330 1041.690 317.510 1042.870 ;
        RECT 317.930 1041.690 319.110 1042.870 ;
        RECT 496.330 3547.010 497.510 3548.190 ;
        RECT 497.930 3547.010 499.110 3548.190 ;
        RECT 496.330 3545.410 497.510 3546.590 ;
        RECT 497.930 3545.410 499.110 3546.590 ;
        RECT 496.330 3383.290 497.510 3384.470 ;
        RECT 497.930 3383.290 499.110 3384.470 ;
        RECT 496.330 3381.690 497.510 3382.870 ;
        RECT 497.930 3381.690 499.110 3382.870 ;
        RECT 496.330 3203.290 497.510 3204.470 ;
        RECT 497.930 3203.290 499.110 3204.470 ;
        RECT 496.330 3201.690 497.510 3202.870 ;
        RECT 497.930 3201.690 499.110 3202.870 ;
        RECT 496.330 3023.290 497.510 3024.470 ;
        RECT 497.930 3023.290 499.110 3024.470 ;
        RECT 496.330 3021.690 497.510 3022.870 ;
        RECT 497.930 3021.690 499.110 3022.870 ;
        RECT 496.330 2843.290 497.510 2844.470 ;
        RECT 497.930 2843.290 499.110 2844.470 ;
        RECT 496.330 2841.690 497.510 2842.870 ;
        RECT 497.930 2841.690 499.110 2842.870 ;
        RECT 496.330 2663.290 497.510 2664.470 ;
        RECT 497.930 2663.290 499.110 2664.470 ;
        RECT 496.330 2661.690 497.510 2662.870 ;
        RECT 497.930 2661.690 499.110 2662.870 ;
        RECT 496.330 2483.290 497.510 2484.470 ;
        RECT 497.930 2483.290 499.110 2484.470 ;
        RECT 496.330 2481.690 497.510 2482.870 ;
        RECT 497.930 2481.690 499.110 2482.870 ;
        RECT 496.330 2303.290 497.510 2304.470 ;
        RECT 497.930 2303.290 499.110 2304.470 ;
        RECT 496.330 2301.690 497.510 2302.870 ;
        RECT 497.930 2301.690 499.110 2302.870 ;
        RECT 496.330 2123.290 497.510 2124.470 ;
        RECT 497.930 2123.290 499.110 2124.470 ;
        RECT 496.330 2121.690 497.510 2122.870 ;
        RECT 497.930 2121.690 499.110 2122.870 ;
        RECT 496.330 1943.290 497.510 1944.470 ;
        RECT 497.930 1943.290 499.110 1944.470 ;
        RECT 496.330 1941.690 497.510 1942.870 ;
        RECT 497.930 1941.690 499.110 1942.870 ;
        RECT 496.330 1763.290 497.510 1764.470 ;
        RECT 497.930 1763.290 499.110 1764.470 ;
        RECT 496.330 1761.690 497.510 1762.870 ;
        RECT 497.930 1761.690 499.110 1762.870 ;
        RECT 496.330 1583.290 497.510 1584.470 ;
        RECT 497.930 1583.290 499.110 1584.470 ;
        RECT 496.330 1581.690 497.510 1582.870 ;
        RECT 497.930 1581.690 499.110 1582.870 ;
        RECT 496.330 1403.290 497.510 1404.470 ;
        RECT 497.930 1403.290 499.110 1404.470 ;
        RECT 496.330 1401.690 497.510 1402.870 ;
        RECT 497.930 1401.690 499.110 1402.870 ;
        RECT 496.330 1223.290 497.510 1224.470 ;
        RECT 497.930 1223.290 499.110 1224.470 ;
        RECT 496.330 1221.690 497.510 1222.870 ;
        RECT 497.930 1221.690 499.110 1222.870 ;
        RECT 496.330 1043.290 497.510 1044.470 ;
        RECT 497.930 1043.290 499.110 1044.470 ;
        RECT 496.330 1041.690 497.510 1042.870 ;
        RECT 497.930 1041.690 499.110 1042.870 ;
        RECT 676.330 3547.010 677.510 3548.190 ;
        RECT 677.930 3547.010 679.110 3548.190 ;
        RECT 676.330 3545.410 677.510 3546.590 ;
        RECT 677.930 3545.410 679.110 3546.590 ;
        RECT 676.330 3383.290 677.510 3384.470 ;
        RECT 677.930 3383.290 679.110 3384.470 ;
        RECT 676.330 3381.690 677.510 3382.870 ;
        RECT 677.930 3381.690 679.110 3382.870 ;
        RECT 676.330 3203.290 677.510 3204.470 ;
        RECT 677.930 3203.290 679.110 3204.470 ;
        RECT 676.330 3201.690 677.510 3202.870 ;
        RECT 677.930 3201.690 679.110 3202.870 ;
        RECT 676.330 3023.290 677.510 3024.470 ;
        RECT 677.930 3023.290 679.110 3024.470 ;
        RECT 676.330 3021.690 677.510 3022.870 ;
        RECT 677.930 3021.690 679.110 3022.870 ;
        RECT 676.330 2843.290 677.510 2844.470 ;
        RECT 677.930 2843.290 679.110 2844.470 ;
        RECT 676.330 2841.690 677.510 2842.870 ;
        RECT 677.930 2841.690 679.110 2842.870 ;
        RECT 676.330 2663.290 677.510 2664.470 ;
        RECT 677.930 2663.290 679.110 2664.470 ;
        RECT 676.330 2661.690 677.510 2662.870 ;
        RECT 677.930 2661.690 679.110 2662.870 ;
        RECT 676.330 2483.290 677.510 2484.470 ;
        RECT 677.930 2483.290 679.110 2484.470 ;
        RECT 676.330 2481.690 677.510 2482.870 ;
        RECT 677.930 2481.690 679.110 2482.870 ;
        RECT 676.330 2303.290 677.510 2304.470 ;
        RECT 677.930 2303.290 679.110 2304.470 ;
        RECT 676.330 2301.690 677.510 2302.870 ;
        RECT 677.930 2301.690 679.110 2302.870 ;
        RECT 676.330 2123.290 677.510 2124.470 ;
        RECT 677.930 2123.290 679.110 2124.470 ;
        RECT 676.330 2121.690 677.510 2122.870 ;
        RECT 677.930 2121.690 679.110 2122.870 ;
        RECT 676.330 1943.290 677.510 1944.470 ;
        RECT 677.930 1943.290 679.110 1944.470 ;
        RECT 676.330 1941.690 677.510 1942.870 ;
        RECT 677.930 1941.690 679.110 1942.870 ;
        RECT 676.330 1763.290 677.510 1764.470 ;
        RECT 677.930 1763.290 679.110 1764.470 ;
        RECT 676.330 1761.690 677.510 1762.870 ;
        RECT 677.930 1761.690 679.110 1762.870 ;
        RECT 676.330 1583.290 677.510 1584.470 ;
        RECT 677.930 1583.290 679.110 1584.470 ;
        RECT 676.330 1581.690 677.510 1582.870 ;
        RECT 677.930 1581.690 679.110 1582.870 ;
        RECT 676.330 1403.290 677.510 1404.470 ;
        RECT 677.930 1403.290 679.110 1404.470 ;
        RECT 676.330 1401.690 677.510 1402.870 ;
        RECT 677.930 1401.690 679.110 1402.870 ;
        RECT 676.330 1223.290 677.510 1224.470 ;
        RECT 677.930 1223.290 679.110 1224.470 ;
        RECT 676.330 1221.690 677.510 1222.870 ;
        RECT 677.930 1221.690 679.110 1222.870 ;
        RECT 676.330 1043.290 677.510 1044.470 ;
        RECT 677.930 1043.290 679.110 1044.470 ;
        RECT 676.330 1041.690 677.510 1042.870 ;
        RECT 677.930 1041.690 679.110 1042.870 ;
        RECT 856.330 3547.010 857.510 3548.190 ;
        RECT 857.930 3547.010 859.110 3548.190 ;
        RECT 856.330 3545.410 857.510 3546.590 ;
        RECT 857.930 3545.410 859.110 3546.590 ;
        RECT 856.330 3383.290 857.510 3384.470 ;
        RECT 857.930 3383.290 859.110 3384.470 ;
        RECT 856.330 3381.690 857.510 3382.870 ;
        RECT 857.930 3381.690 859.110 3382.870 ;
        RECT 856.330 3203.290 857.510 3204.470 ;
        RECT 857.930 3203.290 859.110 3204.470 ;
        RECT 856.330 3201.690 857.510 3202.870 ;
        RECT 857.930 3201.690 859.110 3202.870 ;
        RECT 856.330 3023.290 857.510 3024.470 ;
        RECT 857.930 3023.290 859.110 3024.470 ;
        RECT 856.330 3021.690 857.510 3022.870 ;
        RECT 857.930 3021.690 859.110 3022.870 ;
        RECT 856.330 2843.290 857.510 2844.470 ;
        RECT 857.930 2843.290 859.110 2844.470 ;
        RECT 856.330 2841.690 857.510 2842.870 ;
        RECT 857.930 2841.690 859.110 2842.870 ;
        RECT 856.330 2663.290 857.510 2664.470 ;
        RECT 857.930 2663.290 859.110 2664.470 ;
        RECT 856.330 2661.690 857.510 2662.870 ;
        RECT 857.930 2661.690 859.110 2662.870 ;
        RECT 856.330 2483.290 857.510 2484.470 ;
        RECT 857.930 2483.290 859.110 2484.470 ;
        RECT 856.330 2481.690 857.510 2482.870 ;
        RECT 857.930 2481.690 859.110 2482.870 ;
        RECT 856.330 2303.290 857.510 2304.470 ;
        RECT 857.930 2303.290 859.110 2304.470 ;
        RECT 856.330 2301.690 857.510 2302.870 ;
        RECT 857.930 2301.690 859.110 2302.870 ;
        RECT 856.330 2123.290 857.510 2124.470 ;
        RECT 857.930 2123.290 859.110 2124.470 ;
        RECT 856.330 2121.690 857.510 2122.870 ;
        RECT 857.930 2121.690 859.110 2122.870 ;
        RECT 856.330 1943.290 857.510 1944.470 ;
        RECT 857.930 1943.290 859.110 1944.470 ;
        RECT 856.330 1941.690 857.510 1942.870 ;
        RECT 857.930 1941.690 859.110 1942.870 ;
        RECT 856.330 1763.290 857.510 1764.470 ;
        RECT 857.930 1763.290 859.110 1764.470 ;
        RECT 856.330 1761.690 857.510 1762.870 ;
        RECT 857.930 1761.690 859.110 1762.870 ;
        RECT 856.330 1583.290 857.510 1584.470 ;
        RECT 857.930 1583.290 859.110 1584.470 ;
        RECT 856.330 1581.690 857.510 1582.870 ;
        RECT 857.930 1581.690 859.110 1582.870 ;
        RECT 856.330 1403.290 857.510 1404.470 ;
        RECT 857.930 1403.290 859.110 1404.470 ;
        RECT 856.330 1401.690 857.510 1402.870 ;
        RECT 857.930 1401.690 859.110 1402.870 ;
        RECT 856.330 1223.290 857.510 1224.470 ;
        RECT 857.930 1223.290 859.110 1224.470 ;
        RECT 856.330 1221.690 857.510 1222.870 ;
        RECT 857.930 1221.690 859.110 1222.870 ;
        RECT 856.330 1043.290 857.510 1044.470 ;
        RECT 857.930 1043.290 859.110 1044.470 ;
        RECT 856.330 1041.690 857.510 1042.870 ;
        RECT 857.930 1041.690 859.110 1042.870 ;
        RECT 1036.330 3547.010 1037.510 3548.190 ;
        RECT 1037.930 3547.010 1039.110 3548.190 ;
        RECT 1036.330 3545.410 1037.510 3546.590 ;
        RECT 1037.930 3545.410 1039.110 3546.590 ;
        RECT 1036.330 3383.290 1037.510 3384.470 ;
        RECT 1037.930 3383.290 1039.110 3384.470 ;
        RECT 1036.330 3381.690 1037.510 3382.870 ;
        RECT 1037.930 3381.690 1039.110 3382.870 ;
        RECT 1036.330 3203.290 1037.510 3204.470 ;
        RECT 1037.930 3203.290 1039.110 3204.470 ;
        RECT 1036.330 3201.690 1037.510 3202.870 ;
        RECT 1037.930 3201.690 1039.110 3202.870 ;
        RECT 1036.330 3023.290 1037.510 3024.470 ;
        RECT 1037.930 3023.290 1039.110 3024.470 ;
        RECT 1036.330 3021.690 1037.510 3022.870 ;
        RECT 1037.930 3021.690 1039.110 3022.870 ;
        RECT 1036.330 2843.290 1037.510 2844.470 ;
        RECT 1037.930 2843.290 1039.110 2844.470 ;
        RECT 1036.330 2841.690 1037.510 2842.870 ;
        RECT 1037.930 2841.690 1039.110 2842.870 ;
        RECT 1036.330 2663.290 1037.510 2664.470 ;
        RECT 1037.930 2663.290 1039.110 2664.470 ;
        RECT 1036.330 2661.690 1037.510 2662.870 ;
        RECT 1037.930 2661.690 1039.110 2662.870 ;
        RECT 1036.330 2483.290 1037.510 2484.470 ;
        RECT 1037.930 2483.290 1039.110 2484.470 ;
        RECT 1036.330 2481.690 1037.510 2482.870 ;
        RECT 1037.930 2481.690 1039.110 2482.870 ;
        RECT 1036.330 2303.290 1037.510 2304.470 ;
        RECT 1037.930 2303.290 1039.110 2304.470 ;
        RECT 1036.330 2301.690 1037.510 2302.870 ;
        RECT 1037.930 2301.690 1039.110 2302.870 ;
        RECT 1036.330 2123.290 1037.510 2124.470 ;
        RECT 1037.930 2123.290 1039.110 2124.470 ;
        RECT 1036.330 2121.690 1037.510 2122.870 ;
        RECT 1037.930 2121.690 1039.110 2122.870 ;
        RECT 1036.330 1943.290 1037.510 1944.470 ;
        RECT 1037.930 1943.290 1039.110 1944.470 ;
        RECT 1036.330 1941.690 1037.510 1942.870 ;
        RECT 1037.930 1941.690 1039.110 1942.870 ;
        RECT 1036.330 1763.290 1037.510 1764.470 ;
        RECT 1037.930 1763.290 1039.110 1764.470 ;
        RECT 1036.330 1761.690 1037.510 1762.870 ;
        RECT 1037.930 1761.690 1039.110 1762.870 ;
        RECT 1036.330 1583.290 1037.510 1584.470 ;
        RECT 1037.930 1583.290 1039.110 1584.470 ;
        RECT 1036.330 1581.690 1037.510 1582.870 ;
        RECT 1037.930 1581.690 1039.110 1582.870 ;
        RECT 1036.330 1403.290 1037.510 1404.470 ;
        RECT 1037.930 1403.290 1039.110 1404.470 ;
        RECT 1036.330 1401.690 1037.510 1402.870 ;
        RECT 1037.930 1401.690 1039.110 1402.870 ;
        RECT 1036.330 1223.290 1037.510 1224.470 ;
        RECT 1037.930 1223.290 1039.110 1224.470 ;
        RECT 1036.330 1221.690 1037.510 1222.870 ;
        RECT 1037.930 1221.690 1039.110 1222.870 ;
        RECT 1036.330 1043.290 1037.510 1044.470 ;
        RECT 1037.930 1043.290 1039.110 1044.470 ;
        RECT 1036.330 1041.690 1037.510 1042.870 ;
        RECT 1037.930 1041.690 1039.110 1042.870 ;
        RECT 1216.330 3547.010 1217.510 3548.190 ;
        RECT 1217.930 3547.010 1219.110 3548.190 ;
        RECT 1216.330 3545.410 1217.510 3546.590 ;
        RECT 1217.930 3545.410 1219.110 3546.590 ;
        RECT 1216.330 3383.290 1217.510 3384.470 ;
        RECT 1217.930 3383.290 1219.110 3384.470 ;
        RECT 1216.330 3381.690 1217.510 3382.870 ;
        RECT 1217.930 3381.690 1219.110 3382.870 ;
        RECT 1216.330 3203.290 1217.510 3204.470 ;
        RECT 1217.930 3203.290 1219.110 3204.470 ;
        RECT 1216.330 3201.690 1217.510 3202.870 ;
        RECT 1217.930 3201.690 1219.110 3202.870 ;
        RECT 1216.330 3023.290 1217.510 3024.470 ;
        RECT 1217.930 3023.290 1219.110 3024.470 ;
        RECT 1216.330 3021.690 1217.510 3022.870 ;
        RECT 1217.930 3021.690 1219.110 3022.870 ;
        RECT 1216.330 2843.290 1217.510 2844.470 ;
        RECT 1217.930 2843.290 1219.110 2844.470 ;
        RECT 1216.330 2841.690 1217.510 2842.870 ;
        RECT 1217.930 2841.690 1219.110 2842.870 ;
        RECT 1216.330 2663.290 1217.510 2664.470 ;
        RECT 1217.930 2663.290 1219.110 2664.470 ;
        RECT 1216.330 2661.690 1217.510 2662.870 ;
        RECT 1217.930 2661.690 1219.110 2662.870 ;
        RECT 1216.330 2483.290 1217.510 2484.470 ;
        RECT 1217.930 2483.290 1219.110 2484.470 ;
        RECT 1216.330 2481.690 1217.510 2482.870 ;
        RECT 1217.930 2481.690 1219.110 2482.870 ;
        RECT 1216.330 2303.290 1217.510 2304.470 ;
        RECT 1217.930 2303.290 1219.110 2304.470 ;
        RECT 1216.330 2301.690 1217.510 2302.870 ;
        RECT 1217.930 2301.690 1219.110 2302.870 ;
        RECT 1216.330 2123.290 1217.510 2124.470 ;
        RECT 1217.930 2123.290 1219.110 2124.470 ;
        RECT 1216.330 2121.690 1217.510 2122.870 ;
        RECT 1217.930 2121.690 1219.110 2122.870 ;
        RECT 1216.330 1943.290 1217.510 1944.470 ;
        RECT 1217.930 1943.290 1219.110 1944.470 ;
        RECT 1216.330 1941.690 1217.510 1942.870 ;
        RECT 1217.930 1941.690 1219.110 1942.870 ;
        RECT 1216.330 1763.290 1217.510 1764.470 ;
        RECT 1217.930 1763.290 1219.110 1764.470 ;
        RECT 1216.330 1761.690 1217.510 1762.870 ;
        RECT 1217.930 1761.690 1219.110 1762.870 ;
        RECT 1216.330 1583.290 1217.510 1584.470 ;
        RECT 1217.930 1583.290 1219.110 1584.470 ;
        RECT 1216.330 1581.690 1217.510 1582.870 ;
        RECT 1217.930 1581.690 1219.110 1582.870 ;
        RECT 1216.330 1403.290 1217.510 1404.470 ;
        RECT 1217.930 1403.290 1219.110 1404.470 ;
        RECT 1216.330 1401.690 1217.510 1402.870 ;
        RECT 1217.930 1401.690 1219.110 1402.870 ;
        RECT 1216.330 1223.290 1217.510 1224.470 ;
        RECT 1217.930 1223.290 1219.110 1224.470 ;
        RECT 1216.330 1221.690 1217.510 1222.870 ;
        RECT 1217.930 1221.690 1219.110 1222.870 ;
        RECT 1216.330 1043.290 1217.510 1044.470 ;
        RECT 1217.930 1043.290 1219.110 1044.470 ;
        RECT 1216.330 1041.690 1217.510 1042.870 ;
        RECT 1217.930 1041.690 1219.110 1042.870 ;
        RECT 136.330 863.290 137.510 864.470 ;
        RECT 137.930 863.290 139.110 864.470 ;
        RECT 136.330 861.690 137.510 862.870 ;
        RECT 137.930 861.690 139.110 862.870 ;
        RECT 136.330 683.290 137.510 684.470 ;
        RECT 137.930 683.290 139.110 684.470 ;
        RECT 136.330 681.690 137.510 682.870 ;
        RECT 137.930 681.690 139.110 682.870 ;
        RECT 136.330 503.290 137.510 504.470 ;
        RECT 137.930 503.290 139.110 504.470 ;
        RECT 136.330 501.690 137.510 502.870 ;
        RECT 137.930 501.690 139.110 502.870 ;
        RECT 1216.330 863.290 1217.510 864.470 ;
        RECT 1217.930 863.290 1219.110 864.470 ;
        RECT 1216.330 861.690 1217.510 862.870 ;
        RECT 1217.930 861.690 1219.110 862.870 ;
        RECT 1216.330 683.290 1217.510 684.470 ;
        RECT 1217.930 683.290 1219.110 684.470 ;
        RECT 1216.330 681.690 1217.510 682.870 ;
        RECT 1217.930 681.690 1219.110 682.870 ;
        RECT 1216.330 503.290 1217.510 504.470 ;
        RECT 1217.930 503.290 1219.110 504.470 ;
        RECT 1216.330 501.690 1217.510 502.870 ;
        RECT 1217.930 501.690 1219.110 502.870 ;
        RECT 136.330 323.290 137.510 324.470 ;
        RECT 137.930 323.290 139.110 324.470 ;
        RECT 136.330 321.690 137.510 322.870 ;
        RECT 137.930 321.690 139.110 322.870 ;
        RECT 136.330 143.290 137.510 144.470 ;
        RECT 137.930 143.290 139.110 144.470 ;
        RECT 136.330 141.690 137.510 142.870 ;
        RECT 137.930 141.690 139.110 142.870 ;
        RECT 136.330 -26.910 137.510 -25.730 ;
        RECT 137.930 -26.910 139.110 -25.730 ;
        RECT 136.330 -28.510 137.510 -27.330 ;
        RECT 137.930 -28.510 139.110 -27.330 ;
        RECT 316.330 323.290 317.510 324.470 ;
        RECT 317.930 323.290 319.110 324.470 ;
        RECT 316.330 321.690 317.510 322.870 ;
        RECT 317.930 321.690 319.110 322.870 ;
        RECT 316.330 143.290 317.510 144.470 ;
        RECT 317.930 143.290 319.110 144.470 ;
        RECT 316.330 141.690 317.510 142.870 ;
        RECT 317.930 141.690 319.110 142.870 ;
        RECT 316.330 -26.910 317.510 -25.730 ;
        RECT 317.930 -26.910 319.110 -25.730 ;
        RECT 316.330 -28.510 317.510 -27.330 ;
        RECT 317.930 -28.510 319.110 -27.330 ;
        RECT 496.330 323.290 497.510 324.470 ;
        RECT 497.930 323.290 499.110 324.470 ;
        RECT 496.330 321.690 497.510 322.870 ;
        RECT 497.930 321.690 499.110 322.870 ;
        RECT 496.330 143.290 497.510 144.470 ;
        RECT 497.930 143.290 499.110 144.470 ;
        RECT 496.330 141.690 497.510 142.870 ;
        RECT 497.930 141.690 499.110 142.870 ;
        RECT 496.330 -26.910 497.510 -25.730 ;
        RECT 497.930 -26.910 499.110 -25.730 ;
        RECT 496.330 -28.510 497.510 -27.330 ;
        RECT 497.930 -28.510 499.110 -27.330 ;
        RECT 676.330 323.290 677.510 324.470 ;
        RECT 677.930 323.290 679.110 324.470 ;
        RECT 676.330 321.690 677.510 322.870 ;
        RECT 677.930 321.690 679.110 322.870 ;
        RECT 676.330 143.290 677.510 144.470 ;
        RECT 677.930 143.290 679.110 144.470 ;
        RECT 676.330 141.690 677.510 142.870 ;
        RECT 677.930 141.690 679.110 142.870 ;
        RECT 676.330 -26.910 677.510 -25.730 ;
        RECT 677.930 -26.910 679.110 -25.730 ;
        RECT 676.330 -28.510 677.510 -27.330 ;
        RECT 677.930 -28.510 679.110 -27.330 ;
        RECT 856.330 323.290 857.510 324.470 ;
        RECT 857.930 323.290 859.110 324.470 ;
        RECT 856.330 321.690 857.510 322.870 ;
        RECT 857.930 321.690 859.110 322.870 ;
        RECT 856.330 143.290 857.510 144.470 ;
        RECT 857.930 143.290 859.110 144.470 ;
        RECT 856.330 141.690 857.510 142.870 ;
        RECT 857.930 141.690 859.110 142.870 ;
        RECT 856.330 -26.910 857.510 -25.730 ;
        RECT 857.930 -26.910 859.110 -25.730 ;
        RECT 856.330 -28.510 857.510 -27.330 ;
        RECT 857.930 -28.510 859.110 -27.330 ;
        RECT 1036.330 323.290 1037.510 324.470 ;
        RECT 1037.930 323.290 1039.110 324.470 ;
        RECT 1036.330 321.690 1037.510 322.870 ;
        RECT 1037.930 321.690 1039.110 322.870 ;
        RECT 1036.330 143.290 1037.510 144.470 ;
        RECT 1037.930 143.290 1039.110 144.470 ;
        RECT 1036.330 141.690 1037.510 142.870 ;
        RECT 1037.930 141.690 1039.110 142.870 ;
        RECT 1036.330 -26.910 1037.510 -25.730 ;
        RECT 1037.930 -26.910 1039.110 -25.730 ;
        RECT 1036.330 -28.510 1037.510 -27.330 ;
        RECT 1037.930 -28.510 1039.110 -27.330 ;
        RECT 1216.330 323.290 1217.510 324.470 ;
        RECT 1217.930 323.290 1219.110 324.470 ;
        RECT 1216.330 321.690 1217.510 322.870 ;
        RECT 1217.930 321.690 1219.110 322.870 ;
        RECT 1216.330 143.290 1217.510 144.470 ;
        RECT 1217.930 143.290 1219.110 144.470 ;
        RECT 1216.330 141.690 1217.510 142.870 ;
        RECT 1217.930 141.690 1219.110 142.870 ;
        RECT 1216.330 -26.910 1217.510 -25.730 ;
        RECT 1217.930 -26.910 1219.110 -25.730 ;
        RECT 1216.330 -28.510 1217.510 -27.330 ;
        RECT 1217.930 -28.510 1219.110 -27.330 ;
        RECT 1396.330 3547.010 1397.510 3548.190 ;
        RECT 1397.930 3547.010 1399.110 3548.190 ;
        RECT 1396.330 3545.410 1397.510 3546.590 ;
        RECT 1397.930 3545.410 1399.110 3546.590 ;
        RECT 1396.330 3383.290 1397.510 3384.470 ;
        RECT 1397.930 3383.290 1399.110 3384.470 ;
        RECT 1396.330 3381.690 1397.510 3382.870 ;
        RECT 1397.930 3381.690 1399.110 3382.870 ;
        RECT 1396.330 3203.290 1397.510 3204.470 ;
        RECT 1397.930 3203.290 1399.110 3204.470 ;
        RECT 1396.330 3201.690 1397.510 3202.870 ;
        RECT 1397.930 3201.690 1399.110 3202.870 ;
        RECT 1396.330 3023.290 1397.510 3024.470 ;
        RECT 1397.930 3023.290 1399.110 3024.470 ;
        RECT 1396.330 3021.690 1397.510 3022.870 ;
        RECT 1397.930 3021.690 1399.110 3022.870 ;
        RECT 1396.330 2843.290 1397.510 2844.470 ;
        RECT 1397.930 2843.290 1399.110 2844.470 ;
        RECT 1396.330 2841.690 1397.510 2842.870 ;
        RECT 1397.930 2841.690 1399.110 2842.870 ;
        RECT 1396.330 2663.290 1397.510 2664.470 ;
        RECT 1397.930 2663.290 1399.110 2664.470 ;
        RECT 1396.330 2661.690 1397.510 2662.870 ;
        RECT 1397.930 2661.690 1399.110 2662.870 ;
        RECT 1396.330 2483.290 1397.510 2484.470 ;
        RECT 1397.930 2483.290 1399.110 2484.470 ;
        RECT 1396.330 2481.690 1397.510 2482.870 ;
        RECT 1397.930 2481.690 1399.110 2482.870 ;
        RECT 1396.330 2303.290 1397.510 2304.470 ;
        RECT 1397.930 2303.290 1399.110 2304.470 ;
        RECT 1396.330 2301.690 1397.510 2302.870 ;
        RECT 1397.930 2301.690 1399.110 2302.870 ;
        RECT 1396.330 2123.290 1397.510 2124.470 ;
        RECT 1397.930 2123.290 1399.110 2124.470 ;
        RECT 1396.330 2121.690 1397.510 2122.870 ;
        RECT 1397.930 2121.690 1399.110 2122.870 ;
        RECT 1396.330 1943.290 1397.510 1944.470 ;
        RECT 1397.930 1943.290 1399.110 1944.470 ;
        RECT 1396.330 1941.690 1397.510 1942.870 ;
        RECT 1397.930 1941.690 1399.110 1942.870 ;
        RECT 1396.330 1763.290 1397.510 1764.470 ;
        RECT 1397.930 1763.290 1399.110 1764.470 ;
        RECT 1396.330 1761.690 1397.510 1762.870 ;
        RECT 1397.930 1761.690 1399.110 1762.870 ;
        RECT 1396.330 1583.290 1397.510 1584.470 ;
        RECT 1397.930 1583.290 1399.110 1584.470 ;
        RECT 1396.330 1581.690 1397.510 1582.870 ;
        RECT 1397.930 1581.690 1399.110 1582.870 ;
        RECT 1396.330 1403.290 1397.510 1404.470 ;
        RECT 1397.930 1403.290 1399.110 1404.470 ;
        RECT 1396.330 1401.690 1397.510 1402.870 ;
        RECT 1397.930 1401.690 1399.110 1402.870 ;
        RECT 1396.330 1223.290 1397.510 1224.470 ;
        RECT 1397.930 1223.290 1399.110 1224.470 ;
        RECT 1396.330 1221.690 1397.510 1222.870 ;
        RECT 1397.930 1221.690 1399.110 1222.870 ;
        RECT 1396.330 1043.290 1397.510 1044.470 ;
        RECT 1397.930 1043.290 1399.110 1044.470 ;
        RECT 1396.330 1041.690 1397.510 1042.870 ;
        RECT 1397.930 1041.690 1399.110 1042.870 ;
        RECT 1396.330 863.290 1397.510 864.470 ;
        RECT 1397.930 863.290 1399.110 864.470 ;
        RECT 1396.330 861.690 1397.510 862.870 ;
        RECT 1397.930 861.690 1399.110 862.870 ;
        RECT 1396.330 683.290 1397.510 684.470 ;
        RECT 1397.930 683.290 1399.110 684.470 ;
        RECT 1396.330 681.690 1397.510 682.870 ;
        RECT 1397.930 681.690 1399.110 682.870 ;
        RECT 1396.330 503.290 1397.510 504.470 ;
        RECT 1397.930 503.290 1399.110 504.470 ;
        RECT 1396.330 501.690 1397.510 502.870 ;
        RECT 1397.930 501.690 1399.110 502.870 ;
        RECT 1396.330 323.290 1397.510 324.470 ;
        RECT 1397.930 323.290 1399.110 324.470 ;
        RECT 1396.330 321.690 1397.510 322.870 ;
        RECT 1397.930 321.690 1399.110 322.870 ;
        RECT 1396.330 143.290 1397.510 144.470 ;
        RECT 1397.930 143.290 1399.110 144.470 ;
        RECT 1396.330 141.690 1397.510 142.870 ;
        RECT 1397.930 141.690 1399.110 142.870 ;
        RECT 1396.330 -26.910 1397.510 -25.730 ;
        RECT 1397.930 -26.910 1399.110 -25.730 ;
        RECT 1396.330 -28.510 1397.510 -27.330 ;
        RECT 1397.930 -28.510 1399.110 -27.330 ;
        RECT 1576.330 3547.010 1577.510 3548.190 ;
        RECT 1577.930 3547.010 1579.110 3548.190 ;
        RECT 1576.330 3545.410 1577.510 3546.590 ;
        RECT 1577.930 3545.410 1579.110 3546.590 ;
        RECT 1576.330 3383.290 1577.510 3384.470 ;
        RECT 1577.930 3383.290 1579.110 3384.470 ;
        RECT 1576.330 3381.690 1577.510 3382.870 ;
        RECT 1577.930 3381.690 1579.110 3382.870 ;
        RECT 1576.330 3203.290 1577.510 3204.470 ;
        RECT 1577.930 3203.290 1579.110 3204.470 ;
        RECT 1576.330 3201.690 1577.510 3202.870 ;
        RECT 1577.930 3201.690 1579.110 3202.870 ;
        RECT 1576.330 3023.290 1577.510 3024.470 ;
        RECT 1577.930 3023.290 1579.110 3024.470 ;
        RECT 1576.330 3021.690 1577.510 3022.870 ;
        RECT 1577.930 3021.690 1579.110 3022.870 ;
        RECT 1576.330 2843.290 1577.510 2844.470 ;
        RECT 1577.930 2843.290 1579.110 2844.470 ;
        RECT 1576.330 2841.690 1577.510 2842.870 ;
        RECT 1577.930 2841.690 1579.110 2842.870 ;
        RECT 1576.330 2663.290 1577.510 2664.470 ;
        RECT 1577.930 2663.290 1579.110 2664.470 ;
        RECT 1576.330 2661.690 1577.510 2662.870 ;
        RECT 1577.930 2661.690 1579.110 2662.870 ;
        RECT 1576.330 2483.290 1577.510 2484.470 ;
        RECT 1577.930 2483.290 1579.110 2484.470 ;
        RECT 1576.330 2481.690 1577.510 2482.870 ;
        RECT 1577.930 2481.690 1579.110 2482.870 ;
        RECT 1576.330 2303.290 1577.510 2304.470 ;
        RECT 1577.930 2303.290 1579.110 2304.470 ;
        RECT 1576.330 2301.690 1577.510 2302.870 ;
        RECT 1577.930 2301.690 1579.110 2302.870 ;
        RECT 1576.330 2123.290 1577.510 2124.470 ;
        RECT 1577.930 2123.290 1579.110 2124.470 ;
        RECT 1576.330 2121.690 1577.510 2122.870 ;
        RECT 1577.930 2121.690 1579.110 2122.870 ;
        RECT 1576.330 1943.290 1577.510 1944.470 ;
        RECT 1577.930 1943.290 1579.110 1944.470 ;
        RECT 1576.330 1941.690 1577.510 1942.870 ;
        RECT 1577.930 1941.690 1579.110 1942.870 ;
        RECT 1576.330 1763.290 1577.510 1764.470 ;
        RECT 1577.930 1763.290 1579.110 1764.470 ;
        RECT 1576.330 1761.690 1577.510 1762.870 ;
        RECT 1577.930 1761.690 1579.110 1762.870 ;
        RECT 1576.330 1583.290 1577.510 1584.470 ;
        RECT 1577.930 1583.290 1579.110 1584.470 ;
        RECT 1576.330 1581.690 1577.510 1582.870 ;
        RECT 1577.930 1581.690 1579.110 1582.870 ;
        RECT 1576.330 1403.290 1577.510 1404.470 ;
        RECT 1577.930 1403.290 1579.110 1404.470 ;
        RECT 1576.330 1401.690 1577.510 1402.870 ;
        RECT 1577.930 1401.690 1579.110 1402.870 ;
        RECT 1576.330 1223.290 1577.510 1224.470 ;
        RECT 1577.930 1223.290 1579.110 1224.470 ;
        RECT 1576.330 1221.690 1577.510 1222.870 ;
        RECT 1577.930 1221.690 1579.110 1222.870 ;
        RECT 1576.330 1043.290 1577.510 1044.470 ;
        RECT 1577.930 1043.290 1579.110 1044.470 ;
        RECT 1576.330 1041.690 1577.510 1042.870 ;
        RECT 1577.930 1041.690 1579.110 1042.870 ;
        RECT 1576.330 863.290 1577.510 864.470 ;
        RECT 1577.930 863.290 1579.110 864.470 ;
        RECT 1576.330 861.690 1577.510 862.870 ;
        RECT 1577.930 861.690 1579.110 862.870 ;
        RECT 1576.330 683.290 1577.510 684.470 ;
        RECT 1577.930 683.290 1579.110 684.470 ;
        RECT 1576.330 681.690 1577.510 682.870 ;
        RECT 1577.930 681.690 1579.110 682.870 ;
        RECT 1576.330 503.290 1577.510 504.470 ;
        RECT 1577.930 503.290 1579.110 504.470 ;
        RECT 1576.330 501.690 1577.510 502.870 ;
        RECT 1577.930 501.690 1579.110 502.870 ;
        RECT 1576.330 323.290 1577.510 324.470 ;
        RECT 1577.930 323.290 1579.110 324.470 ;
        RECT 1576.330 321.690 1577.510 322.870 ;
        RECT 1577.930 321.690 1579.110 322.870 ;
        RECT 1576.330 143.290 1577.510 144.470 ;
        RECT 1577.930 143.290 1579.110 144.470 ;
        RECT 1576.330 141.690 1577.510 142.870 ;
        RECT 1577.930 141.690 1579.110 142.870 ;
        RECT 1576.330 -26.910 1577.510 -25.730 ;
        RECT 1577.930 -26.910 1579.110 -25.730 ;
        RECT 1576.330 -28.510 1577.510 -27.330 ;
        RECT 1577.930 -28.510 1579.110 -27.330 ;
        RECT 1756.330 3547.010 1757.510 3548.190 ;
        RECT 1757.930 3547.010 1759.110 3548.190 ;
        RECT 1756.330 3545.410 1757.510 3546.590 ;
        RECT 1757.930 3545.410 1759.110 3546.590 ;
        RECT 1756.330 3383.290 1757.510 3384.470 ;
        RECT 1757.930 3383.290 1759.110 3384.470 ;
        RECT 1756.330 3381.690 1757.510 3382.870 ;
        RECT 1757.930 3381.690 1759.110 3382.870 ;
        RECT 1756.330 3203.290 1757.510 3204.470 ;
        RECT 1757.930 3203.290 1759.110 3204.470 ;
        RECT 1756.330 3201.690 1757.510 3202.870 ;
        RECT 1757.930 3201.690 1759.110 3202.870 ;
        RECT 1756.330 3023.290 1757.510 3024.470 ;
        RECT 1757.930 3023.290 1759.110 3024.470 ;
        RECT 1756.330 3021.690 1757.510 3022.870 ;
        RECT 1757.930 3021.690 1759.110 3022.870 ;
        RECT 1756.330 2843.290 1757.510 2844.470 ;
        RECT 1757.930 2843.290 1759.110 2844.470 ;
        RECT 1756.330 2841.690 1757.510 2842.870 ;
        RECT 1757.930 2841.690 1759.110 2842.870 ;
        RECT 1756.330 2663.290 1757.510 2664.470 ;
        RECT 1757.930 2663.290 1759.110 2664.470 ;
        RECT 1756.330 2661.690 1757.510 2662.870 ;
        RECT 1757.930 2661.690 1759.110 2662.870 ;
        RECT 1756.330 2483.290 1757.510 2484.470 ;
        RECT 1757.930 2483.290 1759.110 2484.470 ;
        RECT 1756.330 2481.690 1757.510 2482.870 ;
        RECT 1757.930 2481.690 1759.110 2482.870 ;
        RECT 1756.330 2303.290 1757.510 2304.470 ;
        RECT 1757.930 2303.290 1759.110 2304.470 ;
        RECT 1756.330 2301.690 1757.510 2302.870 ;
        RECT 1757.930 2301.690 1759.110 2302.870 ;
        RECT 1756.330 2123.290 1757.510 2124.470 ;
        RECT 1757.930 2123.290 1759.110 2124.470 ;
        RECT 1756.330 2121.690 1757.510 2122.870 ;
        RECT 1757.930 2121.690 1759.110 2122.870 ;
        RECT 1756.330 1943.290 1757.510 1944.470 ;
        RECT 1757.930 1943.290 1759.110 1944.470 ;
        RECT 1756.330 1941.690 1757.510 1942.870 ;
        RECT 1757.930 1941.690 1759.110 1942.870 ;
        RECT 1756.330 1763.290 1757.510 1764.470 ;
        RECT 1757.930 1763.290 1759.110 1764.470 ;
        RECT 1756.330 1761.690 1757.510 1762.870 ;
        RECT 1757.930 1761.690 1759.110 1762.870 ;
        RECT 1756.330 1583.290 1757.510 1584.470 ;
        RECT 1757.930 1583.290 1759.110 1584.470 ;
        RECT 1756.330 1581.690 1757.510 1582.870 ;
        RECT 1757.930 1581.690 1759.110 1582.870 ;
        RECT 1756.330 1403.290 1757.510 1404.470 ;
        RECT 1757.930 1403.290 1759.110 1404.470 ;
        RECT 1756.330 1401.690 1757.510 1402.870 ;
        RECT 1757.930 1401.690 1759.110 1402.870 ;
        RECT 1756.330 1223.290 1757.510 1224.470 ;
        RECT 1757.930 1223.290 1759.110 1224.470 ;
        RECT 1756.330 1221.690 1757.510 1222.870 ;
        RECT 1757.930 1221.690 1759.110 1222.870 ;
        RECT 1756.330 1043.290 1757.510 1044.470 ;
        RECT 1757.930 1043.290 1759.110 1044.470 ;
        RECT 1756.330 1041.690 1757.510 1042.870 ;
        RECT 1757.930 1041.690 1759.110 1042.870 ;
        RECT 1756.330 863.290 1757.510 864.470 ;
        RECT 1757.930 863.290 1759.110 864.470 ;
        RECT 1756.330 861.690 1757.510 862.870 ;
        RECT 1757.930 861.690 1759.110 862.870 ;
        RECT 1756.330 683.290 1757.510 684.470 ;
        RECT 1757.930 683.290 1759.110 684.470 ;
        RECT 1756.330 681.690 1757.510 682.870 ;
        RECT 1757.930 681.690 1759.110 682.870 ;
        RECT 1756.330 503.290 1757.510 504.470 ;
        RECT 1757.930 503.290 1759.110 504.470 ;
        RECT 1756.330 501.690 1757.510 502.870 ;
        RECT 1757.930 501.690 1759.110 502.870 ;
        RECT 1756.330 323.290 1757.510 324.470 ;
        RECT 1757.930 323.290 1759.110 324.470 ;
        RECT 1756.330 321.690 1757.510 322.870 ;
        RECT 1757.930 321.690 1759.110 322.870 ;
        RECT 1756.330 143.290 1757.510 144.470 ;
        RECT 1757.930 143.290 1759.110 144.470 ;
        RECT 1756.330 141.690 1757.510 142.870 ;
        RECT 1757.930 141.690 1759.110 142.870 ;
        RECT 1756.330 -26.910 1757.510 -25.730 ;
        RECT 1757.930 -26.910 1759.110 -25.730 ;
        RECT 1756.330 -28.510 1757.510 -27.330 ;
        RECT 1757.930 -28.510 1759.110 -27.330 ;
        RECT 1936.330 3547.010 1937.510 3548.190 ;
        RECT 1937.930 3547.010 1939.110 3548.190 ;
        RECT 1936.330 3545.410 1937.510 3546.590 ;
        RECT 1937.930 3545.410 1939.110 3546.590 ;
        RECT 1936.330 3383.290 1937.510 3384.470 ;
        RECT 1937.930 3383.290 1939.110 3384.470 ;
        RECT 1936.330 3381.690 1937.510 3382.870 ;
        RECT 1937.930 3381.690 1939.110 3382.870 ;
        RECT 1936.330 3203.290 1937.510 3204.470 ;
        RECT 1937.930 3203.290 1939.110 3204.470 ;
        RECT 1936.330 3201.690 1937.510 3202.870 ;
        RECT 1937.930 3201.690 1939.110 3202.870 ;
        RECT 1936.330 3023.290 1937.510 3024.470 ;
        RECT 1937.930 3023.290 1939.110 3024.470 ;
        RECT 1936.330 3021.690 1937.510 3022.870 ;
        RECT 1937.930 3021.690 1939.110 3022.870 ;
        RECT 1936.330 2843.290 1937.510 2844.470 ;
        RECT 1937.930 2843.290 1939.110 2844.470 ;
        RECT 1936.330 2841.690 1937.510 2842.870 ;
        RECT 1937.930 2841.690 1939.110 2842.870 ;
        RECT 1936.330 2663.290 1937.510 2664.470 ;
        RECT 1937.930 2663.290 1939.110 2664.470 ;
        RECT 1936.330 2661.690 1937.510 2662.870 ;
        RECT 1937.930 2661.690 1939.110 2662.870 ;
        RECT 1936.330 2483.290 1937.510 2484.470 ;
        RECT 1937.930 2483.290 1939.110 2484.470 ;
        RECT 1936.330 2481.690 1937.510 2482.870 ;
        RECT 1937.930 2481.690 1939.110 2482.870 ;
        RECT 1936.330 2303.290 1937.510 2304.470 ;
        RECT 1937.930 2303.290 1939.110 2304.470 ;
        RECT 1936.330 2301.690 1937.510 2302.870 ;
        RECT 1937.930 2301.690 1939.110 2302.870 ;
        RECT 1936.330 2123.290 1937.510 2124.470 ;
        RECT 1937.930 2123.290 1939.110 2124.470 ;
        RECT 1936.330 2121.690 1937.510 2122.870 ;
        RECT 1937.930 2121.690 1939.110 2122.870 ;
        RECT 1936.330 1943.290 1937.510 1944.470 ;
        RECT 1937.930 1943.290 1939.110 1944.470 ;
        RECT 1936.330 1941.690 1937.510 1942.870 ;
        RECT 1937.930 1941.690 1939.110 1942.870 ;
        RECT 1936.330 1763.290 1937.510 1764.470 ;
        RECT 1937.930 1763.290 1939.110 1764.470 ;
        RECT 1936.330 1761.690 1937.510 1762.870 ;
        RECT 1937.930 1761.690 1939.110 1762.870 ;
        RECT 1936.330 1583.290 1937.510 1584.470 ;
        RECT 1937.930 1583.290 1939.110 1584.470 ;
        RECT 1936.330 1581.690 1937.510 1582.870 ;
        RECT 1937.930 1581.690 1939.110 1582.870 ;
        RECT 1936.330 1403.290 1937.510 1404.470 ;
        RECT 1937.930 1403.290 1939.110 1404.470 ;
        RECT 1936.330 1401.690 1937.510 1402.870 ;
        RECT 1937.930 1401.690 1939.110 1402.870 ;
        RECT 1936.330 1223.290 1937.510 1224.470 ;
        RECT 1937.930 1223.290 1939.110 1224.470 ;
        RECT 1936.330 1221.690 1937.510 1222.870 ;
        RECT 1937.930 1221.690 1939.110 1222.870 ;
        RECT 1936.330 1043.290 1937.510 1044.470 ;
        RECT 1937.930 1043.290 1939.110 1044.470 ;
        RECT 1936.330 1041.690 1937.510 1042.870 ;
        RECT 1937.930 1041.690 1939.110 1042.870 ;
        RECT 1936.330 863.290 1937.510 864.470 ;
        RECT 1937.930 863.290 1939.110 864.470 ;
        RECT 1936.330 861.690 1937.510 862.870 ;
        RECT 1937.930 861.690 1939.110 862.870 ;
        RECT 1936.330 683.290 1937.510 684.470 ;
        RECT 1937.930 683.290 1939.110 684.470 ;
        RECT 1936.330 681.690 1937.510 682.870 ;
        RECT 1937.930 681.690 1939.110 682.870 ;
        RECT 1936.330 503.290 1937.510 504.470 ;
        RECT 1937.930 503.290 1939.110 504.470 ;
        RECT 1936.330 501.690 1937.510 502.870 ;
        RECT 1937.930 501.690 1939.110 502.870 ;
        RECT 1936.330 323.290 1937.510 324.470 ;
        RECT 1937.930 323.290 1939.110 324.470 ;
        RECT 1936.330 321.690 1937.510 322.870 ;
        RECT 1937.930 321.690 1939.110 322.870 ;
        RECT 1936.330 143.290 1937.510 144.470 ;
        RECT 1937.930 143.290 1939.110 144.470 ;
        RECT 1936.330 141.690 1937.510 142.870 ;
        RECT 1937.930 141.690 1939.110 142.870 ;
        RECT 1936.330 -26.910 1937.510 -25.730 ;
        RECT 1937.930 -26.910 1939.110 -25.730 ;
        RECT 1936.330 -28.510 1937.510 -27.330 ;
        RECT 1937.930 -28.510 1939.110 -27.330 ;
        RECT 2116.330 3547.010 2117.510 3548.190 ;
        RECT 2117.930 3547.010 2119.110 3548.190 ;
        RECT 2116.330 3545.410 2117.510 3546.590 ;
        RECT 2117.930 3545.410 2119.110 3546.590 ;
        RECT 2116.330 3383.290 2117.510 3384.470 ;
        RECT 2117.930 3383.290 2119.110 3384.470 ;
        RECT 2116.330 3381.690 2117.510 3382.870 ;
        RECT 2117.930 3381.690 2119.110 3382.870 ;
        RECT 2116.330 3203.290 2117.510 3204.470 ;
        RECT 2117.930 3203.290 2119.110 3204.470 ;
        RECT 2116.330 3201.690 2117.510 3202.870 ;
        RECT 2117.930 3201.690 2119.110 3202.870 ;
        RECT 2116.330 3023.290 2117.510 3024.470 ;
        RECT 2117.930 3023.290 2119.110 3024.470 ;
        RECT 2116.330 3021.690 2117.510 3022.870 ;
        RECT 2117.930 3021.690 2119.110 3022.870 ;
        RECT 2116.330 2843.290 2117.510 2844.470 ;
        RECT 2117.930 2843.290 2119.110 2844.470 ;
        RECT 2116.330 2841.690 2117.510 2842.870 ;
        RECT 2117.930 2841.690 2119.110 2842.870 ;
        RECT 2116.330 2663.290 2117.510 2664.470 ;
        RECT 2117.930 2663.290 2119.110 2664.470 ;
        RECT 2116.330 2661.690 2117.510 2662.870 ;
        RECT 2117.930 2661.690 2119.110 2662.870 ;
        RECT 2116.330 2483.290 2117.510 2484.470 ;
        RECT 2117.930 2483.290 2119.110 2484.470 ;
        RECT 2116.330 2481.690 2117.510 2482.870 ;
        RECT 2117.930 2481.690 2119.110 2482.870 ;
        RECT 2116.330 2303.290 2117.510 2304.470 ;
        RECT 2117.930 2303.290 2119.110 2304.470 ;
        RECT 2116.330 2301.690 2117.510 2302.870 ;
        RECT 2117.930 2301.690 2119.110 2302.870 ;
        RECT 2116.330 2123.290 2117.510 2124.470 ;
        RECT 2117.930 2123.290 2119.110 2124.470 ;
        RECT 2116.330 2121.690 2117.510 2122.870 ;
        RECT 2117.930 2121.690 2119.110 2122.870 ;
        RECT 2116.330 1943.290 2117.510 1944.470 ;
        RECT 2117.930 1943.290 2119.110 1944.470 ;
        RECT 2116.330 1941.690 2117.510 1942.870 ;
        RECT 2117.930 1941.690 2119.110 1942.870 ;
        RECT 2116.330 1763.290 2117.510 1764.470 ;
        RECT 2117.930 1763.290 2119.110 1764.470 ;
        RECT 2116.330 1761.690 2117.510 1762.870 ;
        RECT 2117.930 1761.690 2119.110 1762.870 ;
        RECT 2116.330 1583.290 2117.510 1584.470 ;
        RECT 2117.930 1583.290 2119.110 1584.470 ;
        RECT 2116.330 1581.690 2117.510 1582.870 ;
        RECT 2117.930 1581.690 2119.110 1582.870 ;
        RECT 2116.330 1403.290 2117.510 1404.470 ;
        RECT 2117.930 1403.290 2119.110 1404.470 ;
        RECT 2116.330 1401.690 2117.510 1402.870 ;
        RECT 2117.930 1401.690 2119.110 1402.870 ;
        RECT 2116.330 1223.290 2117.510 1224.470 ;
        RECT 2117.930 1223.290 2119.110 1224.470 ;
        RECT 2116.330 1221.690 2117.510 1222.870 ;
        RECT 2117.930 1221.690 2119.110 1222.870 ;
        RECT 2116.330 1043.290 2117.510 1044.470 ;
        RECT 2117.930 1043.290 2119.110 1044.470 ;
        RECT 2116.330 1041.690 2117.510 1042.870 ;
        RECT 2117.930 1041.690 2119.110 1042.870 ;
        RECT 2116.330 863.290 2117.510 864.470 ;
        RECT 2117.930 863.290 2119.110 864.470 ;
        RECT 2116.330 861.690 2117.510 862.870 ;
        RECT 2117.930 861.690 2119.110 862.870 ;
        RECT 2116.330 683.290 2117.510 684.470 ;
        RECT 2117.930 683.290 2119.110 684.470 ;
        RECT 2116.330 681.690 2117.510 682.870 ;
        RECT 2117.930 681.690 2119.110 682.870 ;
        RECT 2116.330 503.290 2117.510 504.470 ;
        RECT 2117.930 503.290 2119.110 504.470 ;
        RECT 2116.330 501.690 2117.510 502.870 ;
        RECT 2117.930 501.690 2119.110 502.870 ;
        RECT 2116.330 323.290 2117.510 324.470 ;
        RECT 2117.930 323.290 2119.110 324.470 ;
        RECT 2116.330 321.690 2117.510 322.870 ;
        RECT 2117.930 321.690 2119.110 322.870 ;
        RECT 2116.330 143.290 2117.510 144.470 ;
        RECT 2117.930 143.290 2119.110 144.470 ;
        RECT 2116.330 141.690 2117.510 142.870 ;
        RECT 2117.930 141.690 2119.110 142.870 ;
        RECT 2116.330 -26.910 2117.510 -25.730 ;
        RECT 2117.930 -26.910 2119.110 -25.730 ;
        RECT 2116.330 -28.510 2117.510 -27.330 ;
        RECT 2117.930 -28.510 2119.110 -27.330 ;
        RECT 2296.330 3547.010 2297.510 3548.190 ;
        RECT 2297.930 3547.010 2299.110 3548.190 ;
        RECT 2296.330 3545.410 2297.510 3546.590 ;
        RECT 2297.930 3545.410 2299.110 3546.590 ;
        RECT 2296.330 3383.290 2297.510 3384.470 ;
        RECT 2297.930 3383.290 2299.110 3384.470 ;
        RECT 2296.330 3381.690 2297.510 3382.870 ;
        RECT 2297.930 3381.690 2299.110 3382.870 ;
        RECT 2296.330 3203.290 2297.510 3204.470 ;
        RECT 2297.930 3203.290 2299.110 3204.470 ;
        RECT 2296.330 3201.690 2297.510 3202.870 ;
        RECT 2297.930 3201.690 2299.110 3202.870 ;
        RECT 2296.330 3023.290 2297.510 3024.470 ;
        RECT 2297.930 3023.290 2299.110 3024.470 ;
        RECT 2296.330 3021.690 2297.510 3022.870 ;
        RECT 2297.930 3021.690 2299.110 3022.870 ;
        RECT 2296.330 2843.290 2297.510 2844.470 ;
        RECT 2297.930 2843.290 2299.110 2844.470 ;
        RECT 2296.330 2841.690 2297.510 2842.870 ;
        RECT 2297.930 2841.690 2299.110 2842.870 ;
        RECT 2296.330 2663.290 2297.510 2664.470 ;
        RECT 2297.930 2663.290 2299.110 2664.470 ;
        RECT 2296.330 2661.690 2297.510 2662.870 ;
        RECT 2297.930 2661.690 2299.110 2662.870 ;
        RECT 2296.330 2483.290 2297.510 2484.470 ;
        RECT 2297.930 2483.290 2299.110 2484.470 ;
        RECT 2296.330 2481.690 2297.510 2482.870 ;
        RECT 2297.930 2481.690 2299.110 2482.870 ;
        RECT 2296.330 2303.290 2297.510 2304.470 ;
        RECT 2297.930 2303.290 2299.110 2304.470 ;
        RECT 2296.330 2301.690 2297.510 2302.870 ;
        RECT 2297.930 2301.690 2299.110 2302.870 ;
        RECT 2296.330 2123.290 2297.510 2124.470 ;
        RECT 2297.930 2123.290 2299.110 2124.470 ;
        RECT 2296.330 2121.690 2297.510 2122.870 ;
        RECT 2297.930 2121.690 2299.110 2122.870 ;
        RECT 2296.330 1943.290 2297.510 1944.470 ;
        RECT 2297.930 1943.290 2299.110 1944.470 ;
        RECT 2296.330 1941.690 2297.510 1942.870 ;
        RECT 2297.930 1941.690 2299.110 1942.870 ;
        RECT 2296.330 1763.290 2297.510 1764.470 ;
        RECT 2297.930 1763.290 2299.110 1764.470 ;
        RECT 2296.330 1761.690 2297.510 1762.870 ;
        RECT 2297.930 1761.690 2299.110 1762.870 ;
        RECT 2296.330 1583.290 2297.510 1584.470 ;
        RECT 2297.930 1583.290 2299.110 1584.470 ;
        RECT 2296.330 1581.690 2297.510 1582.870 ;
        RECT 2297.930 1581.690 2299.110 1582.870 ;
        RECT 2296.330 1403.290 2297.510 1404.470 ;
        RECT 2297.930 1403.290 2299.110 1404.470 ;
        RECT 2296.330 1401.690 2297.510 1402.870 ;
        RECT 2297.930 1401.690 2299.110 1402.870 ;
        RECT 2296.330 1223.290 2297.510 1224.470 ;
        RECT 2297.930 1223.290 2299.110 1224.470 ;
        RECT 2296.330 1221.690 2297.510 1222.870 ;
        RECT 2297.930 1221.690 2299.110 1222.870 ;
        RECT 2296.330 1043.290 2297.510 1044.470 ;
        RECT 2297.930 1043.290 2299.110 1044.470 ;
        RECT 2296.330 1041.690 2297.510 1042.870 ;
        RECT 2297.930 1041.690 2299.110 1042.870 ;
        RECT 2296.330 863.290 2297.510 864.470 ;
        RECT 2297.930 863.290 2299.110 864.470 ;
        RECT 2296.330 861.690 2297.510 862.870 ;
        RECT 2297.930 861.690 2299.110 862.870 ;
        RECT 2296.330 683.290 2297.510 684.470 ;
        RECT 2297.930 683.290 2299.110 684.470 ;
        RECT 2296.330 681.690 2297.510 682.870 ;
        RECT 2297.930 681.690 2299.110 682.870 ;
        RECT 2296.330 503.290 2297.510 504.470 ;
        RECT 2297.930 503.290 2299.110 504.470 ;
        RECT 2296.330 501.690 2297.510 502.870 ;
        RECT 2297.930 501.690 2299.110 502.870 ;
        RECT 2296.330 323.290 2297.510 324.470 ;
        RECT 2297.930 323.290 2299.110 324.470 ;
        RECT 2296.330 321.690 2297.510 322.870 ;
        RECT 2297.930 321.690 2299.110 322.870 ;
        RECT 2296.330 143.290 2297.510 144.470 ;
        RECT 2297.930 143.290 2299.110 144.470 ;
        RECT 2296.330 141.690 2297.510 142.870 ;
        RECT 2297.930 141.690 2299.110 142.870 ;
        RECT 2296.330 -26.910 2297.510 -25.730 ;
        RECT 2297.930 -26.910 2299.110 -25.730 ;
        RECT 2296.330 -28.510 2297.510 -27.330 ;
        RECT 2297.930 -28.510 2299.110 -27.330 ;
        RECT 2476.330 3547.010 2477.510 3548.190 ;
        RECT 2477.930 3547.010 2479.110 3548.190 ;
        RECT 2476.330 3545.410 2477.510 3546.590 ;
        RECT 2477.930 3545.410 2479.110 3546.590 ;
        RECT 2476.330 3383.290 2477.510 3384.470 ;
        RECT 2477.930 3383.290 2479.110 3384.470 ;
        RECT 2476.330 3381.690 2477.510 3382.870 ;
        RECT 2477.930 3381.690 2479.110 3382.870 ;
        RECT 2476.330 3203.290 2477.510 3204.470 ;
        RECT 2477.930 3203.290 2479.110 3204.470 ;
        RECT 2476.330 3201.690 2477.510 3202.870 ;
        RECT 2477.930 3201.690 2479.110 3202.870 ;
        RECT 2476.330 3023.290 2477.510 3024.470 ;
        RECT 2477.930 3023.290 2479.110 3024.470 ;
        RECT 2476.330 3021.690 2477.510 3022.870 ;
        RECT 2477.930 3021.690 2479.110 3022.870 ;
        RECT 2476.330 2843.290 2477.510 2844.470 ;
        RECT 2477.930 2843.290 2479.110 2844.470 ;
        RECT 2476.330 2841.690 2477.510 2842.870 ;
        RECT 2477.930 2841.690 2479.110 2842.870 ;
        RECT 2476.330 2663.290 2477.510 2664.470 ;
        RECT 2477.930 2663.290 2479.110 2664.470 ;
        RECT 2476.330 2661.690 2477.510 2662.870 ;
        RECT 2477.930 2661.690 2479.110 2662.870 ;
        RECT 2476.330 2483.290 2477.510 2484.470 ;
        RECT 2477.930 2483.290 2479.110 2484.470 ;
        RECT 2476.330 2481.690 2477.510 2482.870 ;
        RECT 2477.930 2481.690 2479.110 2482.870 ;
        RECT 2476.330 2303.290 2477.510 2304.470 ;
        RECT 2477.930 2303.290 2479.110 2304.470 ;
        RECT 2476.330 2301.690 2477.510 2302.870 ;
        RECT 2477.930 2301.690 2479.110 2302.870 ;
        RECT 2476.330 2123.290 2477.510 2124.470 ;
        RECT 2477.930 2123.290 2479.110 2124.470 ;
        RECT 2476.330 2121.690 2477.510 2122.870 ;
        RECT 2477.930 2121.690 2479.110 2122.870 ;
        RECT 2476.330 1943.290 2477.510 1944.470 ;
        RECT 2477.930 1943.290 2479.110 1944.470 ;
        RECT 2476.330 1941.690 2477.510 1942.870 ;
        RECT 2477.930 1941.690 2479.110 1942.870 ;
        RECT 2476.330 1763.290 2477.510 1764.470 ;
        RECT 2477.930 1763.290 2479.110 1764.470 ;
        RECT 2476.330 1761.690 2477.510 1762.870 ;
        RECT 2477.930 1761.690 2479.110 1762.870 ;
        RECT 2476.330 1583.290 2477.510 1584.470 ;
        RECT 2477.930 1583.290 2479.110 1584.470 ;
        RECT 2476.330 1581.690 2477.510 1582.870 ;
        RECT 2477.930 1581.690 2479.110 1582.870 ;
        RECT 2476.330 1403.290 2477.510 1404.470 ;
        RECT 2477.930 1403.290 2479.110 1404.470 ;
        RECT 2476.330 1401.690 2477.510 1402.870 ;
        RECT 2477.930 1401.690 2479.110 1402.870 ;
        RECT 2476.330 1223.290 2477.510 1224.470 ;
        RECT 2477.930 1223.290 2479.110 1224.470 ;
        RECT 2476.330 1221.690 2477.510 1222.870 ;
        RECT 2477.930 1221.690 2479.110 1222.870 ;
        RECT 2476.330 1043.290 2477.510 1044.470 ;
        RECT 2477.930 1043.290 2479.110 1044.470 ;
        RECT 2476.330 1041.690 2477.510 1042.870 ;
        RECT 2477.930 1041.690 2479.110 1042.870 ;
        RECT 2476.330 863.290 2477.510 864.470 ;
        RECT 2477.930 863.290 2479.110 864.470 ;
        RECT 2476.330 861.690 2477.510 862.870 ;
        RECT 2477.930 861.690 2479.110 862.870 ;
        RECT 2476.330 683.290 2477.510 684.470 ;
        RECT 2477.930 683.290 2479.110 684.470 ;
        RECT 2476.330 681.690 2477.510 682.870 ;
        RECT 2477.930 681.690 2479.110 682.870 ;
        RECT 2476.330 503.290 2477.510 504.470 ;
        RECT 2477.930 503.290 2479.110 504.470 ;
        RECT 2476.330 501.690 2477.510 502.870 ;
        RECT 2477.930 501.690 2479.110 502.870 ;
        RECT 2476.330 323.290 2477.510 324.470 ;
        RECT 2477.930 323.290 2479.110 324.470 ;
        RECT 2476.330 321.690 2477.510 322.870 ;
        RECT 2477.930 321.690 2479.110 322.870 ;
        RECT 2476.330 143.290 2477.510 144.470 ;
        RECT 2477.930 143.290 2479.110 144.470 ;
        RECT 2476.330 141.690 2477.510 142.870 ;
        RECT 2477.930 141.690 2479.110 142.870 ;
        RECT 2476.330 -26.910 2477.510 -25.730 ;
        RECT 2477.930 -26.910 2479.110 -25.730 ;
        RECT 2476.330 -28.510 2477.510 -27.330 ;
        RECT 2477.930 -28.510 2479.110 -27.330 ;
        RECT 2656.330 3547.010 2657.510 3548.190 ;
        RECT 2657.930 3547.010 2659.110 3548.190 ;
        RECT 2656.330 3545.410 2657.510 3546.590 ;
        RECT 2657.930 3545.410 2659.110 3546.590 ;
        RECT 2656.330 3383.290 2657.510 3384.470 ;
        RECT 2657.930 3383.290 2659.110 3384.470 ;
        RECT 2656.330 3381.690 2657.510 3382.870 ;
        RECT 2657.930 3381.690 2659.110 3382.870 ;
        RECT 2656.330 3203.290 2657.510 3204.470 ;
        RECT 2657.930 3203.290 2659.110 3204.470 ;
        RECT 2656.330 3201.690 2657.510 3202.870 ;
        RECT 2657.930 3201.690 2659.110 3202.870 ;
        RECT 2656.330 3023.290 2657.510 3024.470 ;
        RECT 2657.930 3023.290 2659.110 3024.470 ;
        RECT 2656.330 3021.690 2657.510 3022.870 ;
        RECT 2657.930 3021.690 2659.110 3022.870 ;
        RECT 2656.330 2843.290 2657.510 2844.470 ;
        RECT 2657.930 2843.290 2659.110 2844.470 ;
        RECT 2656.330 2841.690 2657.510 2842.870 ;
        RECT 2657.930 2841.690 2659.110 2842.870 ;
        RECT 2656.330 2663.290 2657.510 2664.470 ;
        RECT 2657.930 2663.290 2659.110 2664.470 ;
        RECT 2656.330 2661.690 2657.510 2662.870 ;
        RECT 2657.930 2661.690 2659.110 2662.870 ;
        RECT 2656.330 2483.290 2657.510 2484.470 ;
        RECT 2657.930 2483.290 2659.110 2484.470 ;
        RECT 2656.330 2481.690 2657.510 2482.870 ;
        RECT 2657.930 2481.690 2659.110 2482.870 ;
        RECT 2656.330 2303.290 2657.510 2304.470 ;
        RECT 2657.930 2303.290 2659.110 2304.470 ;
        RECT 2656.330 2301.690 2657.510 2302.870 ;
        RECT 2657.930 2301.690 2659.110 2302.870 ;
        RECT 2656.330 2123.290 2657.510 2124.470 ;
        RECT 2657.930 2123.290 2659.110 2124.470 ;
        RECT 2656.330 2121.690 2657.510 2122.870 ;
        RECT 2657.930 2121.690 2659.110 2122.870 ;
        RECT 2656.330 1943.290 2657.510 1944.470 ;
        RECT 2657.930 1943.290 2659.110 1944.470 ;
        RECT 2656.330 1941.690 2657.510 1942.870 ;
        RECT 2657.930 1941.690 2659.110 1942.870 ;
        RECT 2656.330 1763.290 2657.510 1764.470 ;
        RECT 2657.930 1763.290 2659.110 1764.470 ;
        RECT 2656.330 1761.690 2657.510 1762.870 ;
        RECT 2657.930 1761.690 2659.110 1762.870 ;
        RECT 2656.330 1583.290 2657.510 1584.470 ;
        RECT 2657.930 1583.290 2659.110 1584.470 ;
        RECT 2656.330 1581.690 2657.510 1582.870 ;
        RECT 2657.930 1581.690 2659.110 1582.870 ;
        RECT 2656.330 1403.290 2657.510 1404.470 ;
        RECT 2657.930 1403.290 2659.110 1404.470 ;
        RECT 2656.330 1401.690 2657.510 1402.870 ;
        RECT 2657.930 1401.690 2659.110 1402.870 ;
        RECT 2656.330 1223.290 2657.510 1224.470 ;
        RECT 2657.930 1223.290 2659.110 1224.470 ;
        RECT 2656.330 1221.690 2657.510 1222.870 ;
        RECT 2657.930 1221.690 2659.110 1222.870 ;
        RECT 2656.330 1043.290 2657.510 1044.470 ;
        RECT 2657.930 1043.290 2659.110 1044.470 ;
        RECT 2656.330 1041.690 2657.510 1042.870 ;
        RECT 2657.930 1041.690 2659.110 1042.870 ;
        RECT 2656.330 863.290 2657.510 864.470 ;
        RECT 2657.930 863.290 2659.110 864.470 ;
        RECT 2656.330 861.690 2657.510 862.870 ;
        RECT 2657.930 861.690 2659.110 862.870 ;
        RECT 2656.330 683.290 2657.510 684.470 ;
        RECT 2657.930 683.290 2659.110 684.470 ;
        RECT 2656.330 681.690 2657.510 682.870 ;
        RECT 2657.930 681.690 2659.110 682.870 ;
        RECT 2656.330 503.290 2657.510 504.470 ;
        RECT 2657.930 503.290 2659.110 504.470 ;
        RECT 2656.330 501.690 2657.510 502.870 ;
        RECT 2657.930 501.690 2659.110 502.870 ;
        RECT 2656.330 323.290 2657.510 324.470 ;
        RECT 2657.930 323.290 2659.110 324.470 ;
        RECT 2656.330 321.690 2657.510 322.870 ;
        RECT 2657.930 321.690 2659.110 322.870 ;
        RECT 2656.330 143.290 2657.510 144.470 ;
        RECT 2657.930 143.290 2659.110 144.470 ;
        RECT 2656.330 141.690 2657.510 142.870 ;
        RECT 2657.930 141.690 2659.110 142.870 ;
        RECT 2656.330 -26.910 2657.510 -25.730 ;
        RECT 2657.930 -26.910 2659.110 -25.730 ;
        RECT 2656.330 -28.510 2657.510 -27.330 ;
        RECT 2657.930 -28.510 2659.110 -27.330 ;
        RECT 2836.330 3547.010 2837.510 3548.190 ;
        RECT 2837.930 3547.010 2839.110 3548.190 ;
        RECT 2836.330 3545.410 2837.510 3546.590 ;
        RECT 2837.930 3545.410 2839.110 3546.590 ;
        RECT 2836.330 3383.290 2837.510 3384.470 ;
        RECT 2837.930 3383.290 2839.110 3384.470 ;
        RECT 2836.330 3381.690 2837.510 3382.870 ;
        RECT 2837.930 3381.690 2839.110 3382.870 ;
        RECT 2836.330 3203.290 2837.510 3204.470 ;
        RECT 2837.930 3203.290 2839.110 3204.470 ;
        RECT 2836.330 3201.690 2837.510 3202.870 ;
        RECT 2837.930 3201.690 2839.110 3202.870 ;
        RECT 2836.330 3023.290 2837.510 3024.470 ;
        RECT 2837.930 3023.290 2839.110 3024.470 ;
        RECT 2836.330 3021.690 2837.510 3022.870 ;
        RECT 2837.930 3021.690 2839.110 3022.870 ;
        RECT 2836.330 2843.290 2837.510 2844.470 ;
        RECT 2837.930 2843.290 2839.110 2844.470 ;
        RECT 2836.330 2841.690 2837.510 2842.870 ;
        RECT 2837.930 2841.690 2839.110 2842.870 ;
        RECT 2836.330 2663.290 2837.510 2664.470 ;
        RECT 2837.930 2663.290 2839.110 2664.470 ;
        RECT 2836.330 2661.690 2837.510 2662.870 ;
        RECT 2837.930 2661.690 2839.110 2662.870 ;
        RECT 2836.330 2483.290 2837.510 2484.470 ;
        RECT 2837.930 2483.290 2839.110 2484.470 ;
        RECT 2836.330 2481.690 2837.510 2482.870 ;
        RECT 2837.930 2481.690 2839.110 2482.870 ;
        RECT 2836.330 2303.290 2837.510 2304.470 ;
        RECT 2837.930 2303.290 2839.110 2304.470 ;
        RECT 2836.330 2301.690 2837.510 2302.870 ;
        RECT 2837.930 2301.690 2839.110 2302.870 ;
        RECT 2836.330 2123.290 2837.510 2124.470 ;
        RECT 2837.930 2123.290 2839.110 2124.470 ;
        RECT 2836.330 2121.690 2837.510 2122.870 ;
        RECT 2837.930 2121.690 2839.110 2122.870 ;
        RECT 2836.330 1943.290 2837.510 1944.470 ;
        RECT 2837.930 1943.290 2839.110 1944.470 ;
        RECT 2836.330 1941.690 2837.510 1942.870 ;
        RECT 2837.930 1941.690 2839.110 1942.870 ;
        RECT 2836.330 1763.290 2837.510 1764.470 ;
        RECT 2837.930 1763.290 2839.110 1764.470 ;
        RECT 2836.330 1761.690 2837.510 1762.870 ;
        RECT 2837.930 1761.690 2839.110 1762.870 ;
        RECT 2836.330 1583.290 2837.510 1584.470 ;
        RECT 2837.930 1583.290 2839.110 1584.470 ;
        RECT 2836.330 1581.690 2837.510 1582.870 ;
        RECT 2837.930 1581.690 2839.110 1582.870 ;
        RECT 2836.330 1403.290 2837.510 1404.470 ;
        RECT 2837.930 1403.290 2839.110 1404.470 ;
        RECT 2836.330 1401.690 2837.510 1402.870 ;
        RECT 2837.930 1401.690 2839.110 1402.870 ;
        RECT 2836.330 1223.290 2837.510 1224.470 ;
        RECT 2837.930 1223.290 2839.110 1224.470 ;
        RECT 2836.330 1221.690 2837.510 1222.870 ;
        RECT 2837.930 1221.690 2839.110 1222.870 ;
        RECT 2836.330 1043.290 2837.510 1044.470 ;
        RECT 2837.930 1043.290 2839.110 1044.470 ;
        RECT 2836.330 1041.690 2837.510 1042.870 ;
        RECT 2837.930 1041.690 2839.110 1042.870 ;
        RECT 2836.330 863.290 2837.510 864.470 ;
        RECT 2837.930 863.290 2839.110 864.470 ;
        RECT 2836.330 861.690 2837.510 862.870 ;
        RECT 2837.930 861.690 2839.110 862.870 ;
        RECT 2836.330 683.290 2837.510 684.470 ;
        RECT 2837.930 683.290 2839.110 684.470 ;
        RECT 2836.330 681.690 2837.510 682.870 ;
        RECT 2837.930 681.690 2839.110 682.870 ;
        RECT 2836.330 503.290 2837.510 504.470 ;
        RECT 2837.930 503.290 2839.110 504.470 ;
        RECT 2836.330 501.690 2837.510 502.870 ;
        RECT 2837.930 501.690 2839.110 502.870 ;
        RECT 2836.330 323.290 2837.510 324.470 ;
        RECT 2837.930 323.290 2839.110 324.470 ;
        RECT 2836.330 321.690 2837.510 322.870 ;
        RECT 2837.930 321.690 2839.110 322.870 ;
        RECT 2836.330 143.290 2837.510 144.470 ;
        RECT 2837.930 143.290 2839.110 144.470 ;
        RECT 2836.330 141.690 2837.510 142.870 ;
        RECT 2837.930 141.690 2839.110 142.870 ;
        RECT 2836.330 -26.910 2837.510 -25.730 ;
        RECT 2837.930 -26.910 2839.110 -25.730 ;
        RECT 2836.330 -28.510 2837.510 -27.330 ;
        RECT 2837.930 -28.510 2839.110 -27.330 ;
        RECT 2950.710 3547.010 2951.890 3548.190 ;
        RECT 2952.310 3547.010 2953.490 3548.190 ;
        RECT 2950.710 3545.410 2951.890 3546.590 ;
        RECT 2952.310 3545.410 2953.490 3546.590 ;
        RECT 2950.710 3383.290 2951.890 3384.470 ;
        RECT 2952.310 3383.290 2953.490 3384.470 ;
        RECT 2950.710 3381.690 2951.890 3382.870 ;
        RECT 2952.310 3381.690 2953.490 3382.870 ;
        RECT 2950.710 3203.290 2951.890 3204.470 ;
        RECT 2952.310 3203.290 2953.490 3204.470 ;
        RECT 2950.710 3201.690 2951.890 3202.870 ;
        RECT 2952.310 3201.690 2953.490 3202.870 ;
        RECT 2950.710 3023.290 2951.890 3024.470 ;
        RECT 2952.310 3023.290 2953.490 3024.470 ;
        RECT 2950.710 3021.690 2951.890 3022.870 ;
        RECT 2952.310 3021.690 2953.490 3022.870 ;
        RECT 2950.710 2843.290 2951.890 2844.470 ;
        RECT 2952.310 2843.290 2953.490 2844.470 ;
        RECT 2950.710 2841.690 2951.890 2842.870 ;
        RECT 2952.310 2841.690 2953.490 2842.870 ;
        RECT 2950.710 2663.290 2951.890 2664.470 ;
        RECT 2952.310 2663.290 2953.490 2664.470 ;
        RECT 2950.710 2661.690 2951.890 2662.870 ;
        RECT 2952.310 2661.690 2953.490 2662.870 ;
        RECT 2950.710 2483.290 2951.890 2484.470 ;
        RECT 2952.310 2483.290 2953.490 2484.470 ;
        RECT 2950.710 2481.690 2951.890 2482.870 ;
        RECT 2952.310 2481.690 2953.490 2482.870 ;
        RECT 2950.710 2303.290 2951.890 2304.470 ;
        RECT 2952.310 2303.290 2953.490 2304.470 ;
        RECT 2950.710 2301.690 2951.890 2302.870 ;
        RECT 2952.310 2301.690 2953.490 2302.870 ;
        RECT 2950.710 2123.290 2951.890 2124.470 ;
        RECT 2952.310 2123.290 2953.490 2124.470 ;
        RECT 2950.710 2121.690 2951.890 2122.870 ;
        RECT 2952.310 2121.690 2953.490 2122.870 ;
        RECT 2950.710 1943.290 2951.890 1944.470 ;
        RECT 2952.310 1943.290 2953.490 1944.470 ;
        RECT 2950.710 1941.690 2951.890 1942.870 ;
        RECT 2952.310 1941.690 2953.490 1942.870 ;
        RECT 2950.710 1763.290 2951.890 1764.470 ;
        RECT 2952.310 1763.290 2953.490 1764.470 ;
        RECT 2950.710 1761.690 2951.890 1762.870 ;
        RECT 2952.310 1761.690 2953.490 1762.870 ;
        RECT 2950.710 1583.290 2951.890 1584.470 ;
        RECT 2952.310 1583.290 2953.490 1584.470 ;
        RECT 2950.710 1581.690 2951.890 1582.870 ;
        RECT 2952.310 1581.690 2953.490 1582.870 ;
        RECT 2950.710 1403.290 2951.890 1404.470 ;
        RECT 2952.310 1403.290 2953.490 1404.470 ;
        RECT 2950.710 1401.690 2951.890 1402.870 ;
        RECT 2952.310 1401.690 2953.490 1402.870 ;
        RECT 2950.710 1223.290 2951.890 1224.470 ;
        RECT 2952.310 1223.290 2953.490 1224.470 ;
        RECT 2950.710 1221.690 2951.890 1222.870 ;
        RECT 2952.310 1221.690 2953.490 1222.870 ;
        RECT 2950.710 1043.290 2951.890 1044.470 ;
        RECT 2952.310 1043.290 2953.490 1044.470 ;
        RECT 2950.710 1041.690 2951.890 1042.870 ;
        RECT 2952.310 1041.690 2953.490 1042.870 ;
        RECT 2950.710 863.290 2951.890 864.470 ;
        RECT 2952.310 863.290 2953.490 864.470 ;
        RECT 2950.710 861.690 2951.890 862.870 ;
        RECT 2952.310 861.690 2953.490 862.870 ;
        RECT 2950.710 683.290 2951.890 684.470 ;
        RECT 2952.310 683.290 2953.490 684.470 ;
        RECT 2950.710 681.690 2951.890 682.870 ;
        RECT 2952.310 681.690 2953.490 682.870 ;
        RECT 2950.710 503.290 2951.890 504.470 ;
        RECT 2952.310 503.290 2953.490 504.470 ;
        RECT 2950.710 501.690 2951.890 502.870 ;
        RECT 2952.310 501.690 2953.490 502.870 ;
        RECT 2950.710 323.290 2951.890 324.470 ;
        RECT 2952.310 323.290 2953.490 324.470 ;
        RECT 2950.710 321.690 2951.890 322.870 ;
        RECT 2952.310 321.690 2953.490 322.870 ;
        RECT 2950.710 143.290 2951.890 144.470 ;
        RECT 2952.310 143.290 2953.490 144.470 ;
        RECT 2950.710 141.690 2951.890 142.870 ;
        RECT 2952.310 141.690 2953.490 142.870 ;
        RECT 2950.710 -26.910 2951.890 -25.730 ;
        RECT 2952.310 -26.910 2953.490 -25.730 ;
        RECT 2950.710 -28.510 2951.890 -27.330 ;
        RECT 2952.310 -28.510 2953.490 -27.330 ;
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
        RECT -34.030 861.530 2953.650 864.630 ;
        RECT -34.030 681.530 2953.650 684.630 ;
        RECT -34.030 501.530 2953.650 504.630 ;
        RECT -34.030 321.530 2953.650 324.630 ;
        RECT -34.030 141.530 2953.650 144.630 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
        RECT 334.770 1010.000 337.870 3557.950 ;
        RECT 514.770 1010.000 517.870 3557.950 ;
        RECT 694.770 1010.000 697.870 3557.950 ;
        RECT 874.770 1010.000 877.870 3557.950 ;
        RECT 1054.770 1010.000 1057.870 3557.950 ;
        RECT 334.770 -38.270 337.870 390.000 ;
        RECT 514.770 -38.270 517.870 390.000 ;
        RECT 694.770 -38.270 697.870 390.000 ;
        RECT 874.770 -38.270 877.870 390.000 ;
        RECT 1054.770 -38.270 1057.870 390.000 ;
        RECT 1234.770 -38.270 1237.870 3557.950 ;
        RECT 1414.770 -38.270 1417.870 3557.950 ;
        RECT 1594.770 -38.270 1597.870 3557.950 ;
        RECT 1774.770 -38.270 1777.870 3557.950 ;
        RECT 1954.770 -38.270 1957.870 3557.950 ;
        RECT 2134.770 -38.270 2137.870 3557.950 ;
        RECT 2314.770 -38.270 2317.870 3557.950 ;
        RECT 2494.770 -38.270 2497.870 3557.950 ;
        RECT 2674.770 -38.270 2677.870 3557.950 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
      LAYER via4 ;
        RECT -43.470 3556.610 -42.290 3557.790 ;
        RECT -41.870 3556.610 -40.690 3557.790 ;
        RECT -43.470 3555.010 -42.290 3556.190 ;
        RECT -41.870 3555.010 -40.690 3556.190 ;
        RECT -43.470 3401.890 -42.290 3403.070 ;
        RECT -41.870 3401.890 -40.690 3403.070 ;
        RECT -43.470 3400.290 -42.290 3401.470 ;
        RECT -41.870 3400.290 -40.690 3401.470 ;
        RECT -43.470 3221.890 -42.290 3223.070 ;
        RECT -41.870 3221.890 -40.690 3223.070 ;
        RECT -43.470 3220.290 -42.290 3221.470 ;
        RECT -41.870 3220.290 -40.690 3221.470 ;
        RECT -43.470 3041.890 -42.290 3043.070 ;
        RECT -41.870 3041.890 -40.690 3043.070 ;
        RECT -43.470 3040.290 -42.290 3041.470 ;
        RECT -41.870 3040.290 -40.690 3041.470 ;
        RECT -43.470 2861.890 -42.290 2863.070 ;
        RECT -41.870 2861.890 -40.690 2863.070 ;
        RECT -43.470 2860.290 -42.290 2861.470 ;
        RECT -41.870 2860.290 -40.690 2861.470 ;
        RECT -43.470 2681.890 -42.290 2683.070 ;
        RECT -41.870 2681.890 -40.690 2683.070 ;
        RECT -43.470 2680.290 -42.290 2681.470 ;
        RECT -41.870 2680.290 -40.690 2681.470 ;
        RECT -43.470 2501.890 -42.290 2503.070 ;
        RECT -41.870 2501.890 -40.690 2503.070 ;
        RECT -43.470 2500.290 -42.290 2501.470 ;
        RECT -41.870 2500.290 -40.690 2501.470 ;
        RECT -43.470 2321.890 -42.290 2323.070 ;
        RECT -41.870 2321.890 -40.690 2323.070 ;
        RECT -43.470 2320.290 -42.290 2321.470 ;
        RECT -41.870 2320.290 -40.690 2321.470 ;
        RECT -43.470 2141.890 -42.290 2143.070 ;
        RECT -41.870 2141.890 -40.690 2143.070 ;
        RECT -43.470 2140.290 -42.290 2141.470 ;
        RECT -41.870 2140.290 -40.690 2141.470 ;
        RECT -43.470 1961.890 -42.290 1963.070 ;
        RECT -41.870 1961.890 -40.690 1963.070 ;
        RECT -43.470 1960.290 -42.290 1961.470 ;
        RECT -41.870 1960.290 -40.690 1961.470 ;
        RECT -43.470 1781.890 -42.290 1783.070 ;
        RECT -41.870 1781.890 -40.690 1783.070 ;
        RECT -43.470 1780.290 -42.290 1781.470 ;
        RECT -41.870 1780.290 -40.690 1781.470 ;
        RECT -43.470 1601.890 -42.290 1603.070 ;
        RECT -41.870 1601.890 -40.690 1603.070 ;
        RECT -43.470 1600.290 -42.290 1601.470 ;
        RECT -41.870 1600.290 -40.690 1601.470 ;
        RECT -43.470 1421.890 -42.290 1423.070 ;
        RECT -41.870 1421.890 -40.690 1423.070 ;
        RECT -43.470 1420.290 -42.290 1421.470 ;
        RECT -41.870 1420.290 -40.690 1421.470 ;
        RECT -43.470 1241.890 -42.290 1243.070 ;
        RECT -41.870 1241.890 -40.690 1243.070 ;
        RECT -43.470 1240.290 -42.290 1241.470 ;
        RECT -41.870 1240.290 -40.690 1241.470 ;
        RECT -43.470 1061.890 -42.290 1063.070 ;
        RECT -41.870 1061.890 -40.690 1063.070 ;
        RECT -43.470 1060.290 -42.290 1061.470 ;
        RECT -41.870 1060.290 -40.690 1061.470 ;
        RECT -43.470 881.890 -42.290 883.070 ;
        RECT -41.870 881.890 -40.690 883.070 ;
        RECT -43.470 880.290 -42.290 881.470 ;
        RECT -41.870 880.290 -40.690 881.470 ;
        RECT -43.470 701.890 -42.290 703.070 ;
        RECT -41.870 701.890 -40.690 703.070 ;
        RECT -43.470 700.290 -42.290 701.470 ;
        RECT -41.870 700.290 -40.690 701.470 ;
        RECT -43.470 521.890 -42.290 523.070 ;
        RECT -41.870 521.890 -40.690 523.070 ;
        RECT -43.470 520.290 -42.290 521.470 ;
        RECT -41.870 520.290 -40.690 521.470 ;
        RECT -43.470 341.890 -42.290 343.070 ;
        RECT -41.870 341.890 -40.690 343.070 ;
        RECT -43.470 340.290 -42.290 341.470 ;
        RECT -41.870 340.290 -40.690 341.470 ;
        RECT -43.470 161.890 -42.290 163.070 ;
        RECT -41.870 161.890 -40.690 163.070 ;
        RECT -43.470 160.290 -42.290 161.470 ;
        RECT -41.870 160.290 -40.690 161.470 ;
        RECT -43.470 -36.510 -42.290 -35.330 ;
        RECT -41.870 -36.510 -40.690 -35.330 ;
        RECT -43.470 -38.110 -42.290 -36.930 ;
        RECT -41.870 -38.110 -40.690 -36.930 ;
        RECT 154.930 3556.610 156.110 3557.790 ;
        RECT 156.530 3556.610 157.710 3557.790 ;
        RECT 154.930 3555.010 156.110 3556.190 ;
        RECT 156.530 3555.010 157.710 3556.190 ;
        RECT 154.930 3401.890 156.110 3403.070 ;
        RECT 156.530 3401.890 157.710 3403.070 ;
        RECT 154.930 3400.290 156.110 3401.470 ;
        RECT 156.530 3400.290 157.710 3401.470 ;
        RECT 154.930 3221.890 156.110 3223.070 ;
        RECT 156.530 3221.890 157.710 3223.070 ;
        RECT 154.930 3220.290 156.110 3221.470 ;
        RECT 156.530 3220.290 157.710 3221.470 ;
        RECT 154.930 3041.890 156.110 3043.070 ;
        RECT 156.530 3041.890 157.710 3043.070 ;
        RECT 154.930 3040.290 156.110 3041.470 ;
        RECT 156.530 3040.290 157.710 3041.470 ;
        RECT 154.930 2861.890 156.110 2863.070 ;
        RECT 156.530 2861.890 157.710 2863.070 ;
        RECT 154.930 2860.290 156.110 2861.470 ;
        RECT 156.530 2860.290 157.710 2861.470 ;
        RECT 154.930 2681.890 156.110 2683.070 ;
        RECT 156.530 2681.890 157.710 2683.070 ;
        RECT 154.930 2680.290 156.110 2681.470 ;
        RECT 156.530 2680.290 157.710 2681.470 ;
        RECT 154.930 2501.890 156.110 2503.070 ;
        RECT 156.530 2501.890 157.710 2503.070 ;
        RECT 154.930 2500.290 156.110 2501.470 ;
        RECT 156.530 2500.290 157.710 2501.470 ;
        RECT 154.930 2321.890 156.110 2323.070 ;
        RECT 156.530 2321.890 157.710 2323.070 ;
        RECT 154.930 2320.290 156.110 2321.470 ;
        RECT 156.530 2320.290 157.710 2321.470 ;
        RECT 154.930 2141.890 156.110 2143.070 ;
        RECT 156.530 2141.890 157.710 2143.070 ;
        RECT 154.930 2140.290 156.110 2141.470 ;
        RECT 156.530 2140.290 157.710 2141.470 ;
        RECT 154.930 1961.890 156.110 1963.070 ;
        RECT 156.530 1961.890 157.710 1963.070 ;
        RECT 154.930 1960.290 156.110 1961.470 ;
        RECT 156.530 1960.290 157.710 1961.470 ;
        RECT 154.930 1781.890 156.110 1783.070 ;
        RECT 156.530 1781.890 157.710 1783.070 ;
        RECT 154.930 1780.290 156.110 1781.470 ;
        RECT 156.530 1780.290 157.710 1781.470 ;
        RECT 154.930 1601.890 156.110 1603.070 ;
        RECT 156.530 1601.890 157.710 1603.070 ;
        RECT 154.930 1600.290 156.110 1601.470 ;
        RECT 156.530 1600.290 157.710 1601.470 ;
        RECT 154.930 1421.890 156.110 1423.070 ;
        RECT 156.530 1421.890 157.710 1423.070 ;
        RECT 154.930 1420.290 156.110 1421.470 ;
        RECT 156.530 1420.290 157.710 1421.470 ;
        RECT 154.930 1241.890 156.110 1243.070 ;
        RECT 156.530 1241.890 157.710 1243.070 ;
        RECT 154.930 1240.290 156.110 1241.470 ;
        RECT 156.530 1240.290 157.710 1241.470 ;
        RECT 154.930 1061.890 156.110 1063.070 ;
        RECT 156.530 1061.890 157.710 1063.070 ;
        RECT 154.930 1060.290 156.110 1061.470 ;
        RECT 156.530 1060.290 157.710 1061.470 ;
        RECT 334.930 3556.610 336.110 3557.790 ;
        RECT 336.530 3556.610 337.710 3557.790 ;
        RECT 334.930 3555.010 336.110 3556.190 ;
        RECT 336.530 3555.010 337.710 3556.190 ;
        RECT 334.930 3401.890 336.110 3403.070 ;
        RECT 336.530 3401.890 337.710 3403.070 ;
        RECT 334.930 3400.290 336.110 3401.470 ;
        RECT 336.530 3400.290 337.710 3401.470 ;
        RECT 334.930 3221.890 336.110 3223.070 ;
        RECT 336.530 3221.890 337.710 3223.070 ;
        RECT 334.930 3220.290 336.110 3221.470 ;
        RECT 336.530 3220.290 337.710 3221.470 ;
        RECT 334.930 3041.890 336.110 3043.070 ;
        RECT 336.530 3041.890 337.710 3043.070 ;
        RECT 334.930 3040.290 336.110 3041.470 ;
        RECT 336.530 3040.290 337.710 3041.470 ;
        RECT 334.930 2861.890 336.110 2863.070 ;
        RECT 336.530 2861.890 337.710 2863.070 ;
        RECT 334.930 2860.290 336.110 2861.470 ;
        RECT 336.530 2860.290 337.710 2861.470 ;
        RECT 334.930 2681.890 336.110 2683.070 ;
        RECT 336.530 2681.890 337.710 2683.070 ;
        RECT 334.930 2680.290 336.110 2681.470 ;
        RECT 336.530 2680.290 337.710 2681.470 ;
        RECT 334.930 2501.890 336.110 2503.070 ;
        RECT 336.530 2501.890 337.710 2503.070 ;
        RECT 334.930 2500.290 336.110 2501.470 ;
        RECT 336.530 2500.290 337.710 2501.470 ;
        RECT 334.930 2321.890 336.110 2323.070 ;
        RECT 336.530 2321.890 337.710 2323.070 ;
        RECT 334.930 2320.290 336.110 2321.470 ;
        RECT 336.530 2320.290 337.710 2321.470 ;
        RECT 334.930 2141.890 336.110 2143.070 ;
        RECT 336.530 2141.890 337.710 2143.070 ;
        RECT 334.930 2140.290 336.110 2141.470 ;
        RECT 336.530 2140.290 337.710 2141.470 ;
        RECT 334.930 1961.890 336.110 1963.070 ;
        RECT 336.530 1961.890 337.710 1963.070 ;
        RECT 334.930 1960.290 336.110 1961.470 ;
        RECT 336.530 1960.290 337.710 1961.470 ;
        RECT 334.930 1781.890 336.110 1783.070 ;
        RECT 336.530 1781.890 337.710 1783.070 ;
        RECT 334.930 1780.290 336.110 1781.470 ;
        RECT 336.530 1780.290 337.710 1781.470 ;
        RECT 334.930 1601.890 336.110 1603.070 ;
        RECT 336.530 1601.890 337.710 1603.070 ;
        RECT 334.930 1600.290 336.110 1601.470 ;
        RECT 336.530 1600.290 337.710 1601.470 ;
        RECT 334.930 1421.890 336.110 1423.070 ;
        RECT 336.530 1421.890 337.710 1423.070 ;
        RECT 334.930 1420.290 336.110 1421.470 ;
        RECT 336.530 1420.290 337.710 1421.470 ;
        RECT 334.930 1241.890 336.110 1243.070 ;
        RECT 336.530 1241.890 337.710 1243.070 ;
        RECT 334.930 1240.290 336.110 1241.470 ;
        RECT 336.530 1240.290 337.710 1241.470 ;
        RECT 334.930 1061.890 336.110 1063.070 ;
        RECT 336.530 1061.890 337.710 1063.070 ;
        RECT 334.930 1060.290 336.110 1061.470 ;
        RECT 336.530 1060.290 337.710 1061.470 ;
        RECT 514.930 3556.610 516.110 3557.790 ;
        RECT 516.530 3556.610 517.710 3557.790 ;
        RECT 514.930 3555.010 516.110 3556.190 ;
        RECT 516.530 3555.010 517.710 3556.190 ;
        RECT 514.930 3401.890 516.110 3403.070 ;
        RECT 516.530 3401.890 517.710 3403.070 ;
        RECT 514.930 3400.290 516.110 3401.470 ;
        RECT 516.530 3400.290 517.710 3401.470 ;
        RECT 514.930 3221.890 516.110 3223.070 ;
        RECT 516.530 3221.890 517.710 3223.070 ;
        RECT 514.930 3220.290 516.110 3221.470 ;
        RECT 516.530 3220.290 517.710 3221.470 ;
        RECT 514.930 3041.890 516.110 3043.070 ;
        RECT 516.530 3041.890 517.710 3043.070 ;
        RECT 514.930 3040.290 516.110 3041.470 ;
        RECT 516.530 3040.290 517.710 3041.470 ;
        RECT 514.930 2861.890 516.110 2863.070 ;
        RECT 516.530 2861.890 517.710 2863.070 ;
        RECT 514.930 2860.290 516.110 2861.470 ;
        RECT 516.530 2860.290 517.710 2861.470 ;
        RECT 514.930 2681.890 516.110 2683.070 ;
        RECT 516.530 2681.890 517.710 2683.070 ;
        RECT 514.930 2680.290 516.110 2681.470 ;
        RECT 516.530 2680.290 517.710 2681.470 ;
        RECT 514.930 2501.890 516.110 2503.070 ;
        RECT 516.530 2501.890 517.710 2503.070 ;
        RECT 514.930 2500.290 516.110 2501.470 ;
        RECT 516.530 2500.290 517.710 2501.470 ;
        RECT 514.930 2321.890 516.110 2323.070 ;
        RECT 516.530 2321.890 517.710 2323.070 ;
        RECT 514.930 2320.290 516.110 2321.470 ;
        RECT 516.530 2320.290 517.710 2321.470 ;
        RECT 514.930 2141.890 516.110 2143.070 ;
        RECT 516.530 2141.890 517.710 2143.070 ;
        RECT 514.930 2140.290 516.110 2141.470 ;
        RECT 516.530 2140.290 517.710 2141.470 ;
        RECT 514.930 1961.890 516.110 1963.070 ;
        RECT 516.530 1961.890 517.710 1963.070 ;
        RECT 514.930 1960.290 516.110 1961.470 ;
        RECT 516.530 1960.290 517.710 1961.470 ;
        RECT 514.930 1781.890 516.110 1783.070 ;
        RECT 516.530 1781.890 517.710 1783.070 ;
        RECT 514.930 1780.290 516.110 1781.470 ;
        RECT 516.530 1780.290 517.710 1781.470 ;
        RECT 514.930 1601.890 516.110 1603.070 ;
        RECT 516.530 1601.890 517.710 1603.070 ;
        RECT 514.930 1600.290 516.110 1601.470 ;
        RECT 516.530 1600.290 517.710 1601.470 ;
        RECT 514.930 1421.890 516.110 1423.070 ;
        RECT 516.530 1421.890 517.710 1423.070 ;
        RECT 514.930 1420.290 516.110 1421.470 ;
        RECT 516.530 1420.290 517.710 1421.470 ;
        RECT 514.930 1241.890 516.110 1243.070 ;
        RECT 516.530 1241.890 517.710 1243.070 ;
        RECT 514.930 1240.290 516.110 1241.470 ;
        RECT 516.530 1240.290 517.710 1241.470 ;
        RECT 514.930 1061.890 516.110 1063.070 ;
        RECT 516.530 1061.890 517.710 1063.070 ;
        RECT 514.930 1060.290 516.110 1061.470 ;
        RECT 516.530 1060.290 517.710 1061.470 ;
        RECT 694.930 3556.610 696.110 3557.790 ;
        RECT 696.530 3556.610 697.710 3557.790 ;
        RECT 694.930 3555.010 696.110 3556.190 ;
        RECT 696.530 3555.010 697.710 3556.190 ;
        RECT 694.930 3401.890 696.110 3403.070 ;
        RECT 696.530 3401.890 697.710 3403.070 ;
        RECT 694.930 3400.290 696.110 3401.470 ;
        RECT 696.530 3400.290 697.710 3401.470 ;
        RECT 694.930 3221.890 696.110 3223.070 ;
        RECT 696.530 3221.890 697.710 3223.070 ;
        RECT 694.930 3220.290 696.110 3221.470 ;
        RECT 696.530 3220.290 697.710 3221.470 ;
        RECT 694.930 3041.890 696.110 3043.070 ;
        RECT 696.530 3041.890 697.710 3043.070 ;
        RECT 694.930 3040.290 696.110 3041.470 ;
        RECT 696.530 3040.290 697.710 3041.470 ;
        RECT 694.930 2861.890 696.110 2863.070 ;
        RECT 696.530 2861.890 697.710 2863.070 ;
        RECT 694.930 2860.290 696.110 2861.470 ;
        RECT 696.530 2860.290 697.710 2861.470 ;
        RECT 694.930 2681.890 696.110 2683.070 ;
        RECT 696.530 2681.890 697.710 2683.070 ;
        RECT 694.930 2680.290 696.110 2681.470 ;
        RECT 696.530 2680.290 697.710 2681.470 ;
        RECT 694.930 2501.890 696.110 2503.070 ;
        RECT 696.530 2501.890 697.710 2503.070 ;
        RECT 694.930 2500.290 696.110 2501.470 ;
        RECT 696.530 2500.290 697.710 2501.470 ;
        RECT 694.930 2321.890 696.110 2323.070 ;
        RECT 696.530 2321.890 697.710 2323.070 ;
        RECT 694.930 2320.290 696.110 2321.470 ;
        RECT 696.530 2320.290 697.710 2321.470 ;
        RECT 694.930 2141.890 696.110 2143.070 ;
        RECT 696.530 2141.890 697.710 2143.070 ;
        RECT 694.930 2140.290 696.110 2141.470 ;
        RECT 696.530 2140.290 697.710 2141.470 ;
        RECT 694.930 1961.890 696.110 1963.070 ;
        RECT 696.530 1961.890 697.710 1963.070 ;
        RECT 694.930 1960.290 696.110 1961.470 ;
        RECT 696.530 1960.290 697.710 1961.470 ;
        RECT 694.930 1781.890 696.110 1783.070 ;
        RECT 696.530 1781.890 697.710 1783.070 ;
        RECT 694.930 1780.290 696.110 1781.470 ;
        RECT 696.530 1780.290 697.710 1781.470 ;
        RECT 694.930 1601.890 696.110 1603.070 ;
        RECT 696.530 1601.890 697.710 1603.070 ;
        RECT 694.930 1600.290 696.110 1601.470 ;
        RECT 696.530 1600.290 697.710 1601.470 ;
        RECT 694.930 1421.890 696.110 1423.070 ;
        RECT 696.530 1421.890 697.710 1423.070 ;
        RECT 694.930 1420.290 696.110 1421.470 ;
        RECT 696.530 1420.290 697.710 1421.470 ;
        RECT 694.930 1241.890 696.110 1243.070 ;
        RECT 696.530 1241.890 697.710 1243.070 ;
        RECT 694.930 1240.290 696.110 1241.470 ;
        RECT 696.530 1240.290 697.710 1241.470 ;
        RECT 694.930 1061.890 696.110 1063.070 ;
        RECT 696.530 1061.890 697.710 1063.070 ;
        RECT 694.930 1060.290 696.110 1061.470 ;
        RECT 696.530 1060.290 697.710 1061.470 ;
        RECT 874.930 3556.610 876.110 3557.790 ;
        RECT 876.530 3556.610 877.710 3557.790 ;
        RECT 874.930 3555.010 876.110 3556.190 ;
        RECT 876.530 3555.010 877.710 3556.190 ;
        RECT 874.930 3401.890 876.110 3403.070 ;
        RECT 876.530 3401.890 877.710 3403.070 ;
        RECT 874.930 3400.290 876.110 3401.470 ;
        RECT 876.530 3400.290 877.710 3401.470 ;
        RECT 874.930 3221.890 876.110 3223.070 ;
        RECT 876.530 3221.890 877.710 3223.070 ;
        RECT 874.930 3220.290 876.110 3221.470 ;
        RECT 876.530 3220.290 877.710 3221.470 ;
        RECT 874.930 3041.890 876.110 3043.070 ;
        RECT 876.530 3041.890 877.710 3043.070 ;
        RECT 874.930 3040.290 876.110 3041.470 ;
        RECT 876.530 3040.290 877.710 3041.470 ;
        RECT 874.930 2861.890 876.110 2863.070 ;
        RECT 876.530 2861.890 877.710 2863.070 ;
        RECT 874.930 2860.290 876.110 2861.470 ;
        RECT 876.530 2860.290 877.710 2861.470 ;
        RECT 874.930 2681.890 876.110 2683.070 ;
        RECT 876.530 2681.890 877.710 2683.070 ;
        RECT 874.930 2680.290 876.110 2681.470 ;
        RECT 876.530 2680.290 877.710 2681.470 ;
        RECT 874.930 2501.890 876.110 2503.070 ;
        RECT 876.530 2501.890 877.710 2503.070 ;
        RECT 874.930 2500.290 876.110 2501.470 ;
        RECT 876.530 2500.290 877.710 2501.470 ;
        RECT 874.930 2321.890 876.110 2323.070 ;
        RECT 876.530 2321.890 877.710 2323.070 ;
        RECT 874.930 2320.290 876.110 2321.470 ;
        RECT 876.530 2320.290 877.710 2321.470 ;
        RECT 874.930 2141.890 876.110 2143.070 ;
        RECT 876.530 2141.890 877.710 2143.070 ;
        RECT 874.930 2140.290 876.110 2141.470 ;
        RECT 876.530 2140.290 877.710 2141.470 ;
        RECT 874.930 1961.890 876.110 1963.070 ;
        RECT 876.530 1961.890 877.710 1963.070 ;
        RECT 874.930 1960.290 876.110 1961.470 ;
        RECT 876.530 1960.290 877.710 1961.470 ;
        RECT 874.930 1781.890 876.110 1783.070 ;
        RECT 876.530 1781.890 877.710 1783.070 ;
        RECT 874.930 1780.290 876.110 1781.470 ;
        RECT 876.530 1780.290 877.710 1781.470 ;
        RECT 874.930 1601.890 876.110 1603.070 ;
        RECT 876.530 1601.890 877.710 1603.070 ;
        RECT 874.930 1600.290 876.110 1601.470 ;
        RECT 876.530 1600.290 877.710 1601.470 ;
        RECT 874.930 1421.890 876.110 1423.070 ;
        RECT 876.530 1421.890 877.710 1423.070 ;
        RECT 874.930 1420.290 876.110 1421.470 ;
        RECT 876.530 1420.290 877.710 1421.470 ;
        RECT 874.930 1241.890 876.110 1243.070 ;
        RECT 876.530 1241.890 877.710 1243.070 ;
        RECT 874.930 1240.290 876.110 1241.470 ;
        RECT 876.530 1240.290 877.710 1241.470 ;
        RECT 874.930 1061.890 876.110 1063.070 ;
        RECT 876.530 1061.890 877.710 1063.070 ;
        RECT 874.930 1060.290 876.110 1061.470 ;
        RECT 876.530 1060.290 877.710 1061.470 ;
        RECT 1054.930 3556.610 1056.110 3557.790 ;
        RECT 1056.530 3556.610 1057.710 3557.790 ;
        RECT 1054.930 3555.010 1056.110 3556.190 ;
        RECT 1056.530 3555.010 1057.710 3556.190 ;
        RECT 1054.930 3401.890 1056.110 3403.070 ;
        RECT 1056.530 3401.890 1057.710 3403.070 ;
        RECT 1054.930 3400.290 1056.110 3401.470 ;
        RECT 1056.530 3400.290 1057.710 3401.470 ;
        RECT 1054.930 3221.890 1056.110 3223.070 ;
        RECT 1056.530 3221.890 1057.710 3223.070 ;
        RECT 1054.930 3220.290 1056.110 3221.470 ;
        RECT 1056.530 3220.290 1057.710 3221.470 ;
        RECT 1054.930 3041.890 1056.110 3043.070 ;
        RECT 1056.530 3041.890 1057.710 3043.070 ;
        RECT 1054.930 3040.290 1056.110 3041.470 ;
        RECT 1056.530 3040.290 1057.710 3041.470 ;
        RECT 1054.930 2861.890 1056.110 2863.070 ;
        RECT 1056.530 2861.890 1057.710 2863.070 ;
        RECT 1054.930 2860.290 1056.110 2861.470 ;
        RECT 1056.530 2860.290 1057.710 2861.470 ;
        RECT 1054.930 2681.890 1056.110 2683.070 ;
        RECT 1056.530 2681.890 1057.710 2683.070 ;
        RECT 1054.930 2680.290 1056.110 2681.470 ;
        RECT 1056.530 2680.290 1057.710 2681.470 ;
        RECT 1054.930 2501.890 1056.110 2503.070 ;
        RECT 1056.530 2501.890 1057.710 2503.070 ;
        RECT 1054.930 2500.290 1056.110 2501.470 ;
        RECT 1056.530 2500.290 1057.710 2501.470 ;
        RECT 1054.930 2321.890 1056.110 2323.070 ;
        RECT 1056.530 2321.890 1057.710 2323.070 ;
        RECT 1054.930 2320.290 1056.110 2321.470 ;
        RECT 1056.530 2320.290 1057.710 2321.470 ;
        RECT 1054.930 2141.890 1056.110 2143.070 ;
        RECT 1056.530 2141.890 1057.710 2143.070 ;
        RECT 1054.930 2140.290 1056.110 2141.470 ;
        RECT 1056.530 2140.290 1057.710 2141.470 ;
        RECT 1054.930 1961.890 1056.110 1963.070 ;
        RECT 1056.530 1961.890 1057.710 1963.070 ;
        RECT 1054.930 1960.290 1056.110 1961.470 ;
        RECT 1056.530 1960.290 1057.710 1961.470 ;
        RECT 1054.930 1781.890 1056.110 1783.070 ;
        RECT 1056.530 1781.890 1057.710 1783.070 ;
        RECT 1054.930 1780.290 1056.110 1781.470 ;
        RECT 1056.530 1780.290 1057.710 1781.470 ;
        RECT 1054.930 1601.890 1056.110 1603.070 ;
        RECT 1056.530 1601.890 1057.710 1603.070 ;
        RECT 1054.930 1600.290 1056.110 1601.470 ;
        RECT 1056.530 1600.290 1057.710 1601.470 ;
        RECT 1054.930 1421.890 1056.110 1423.070 ;
        RECT 1056.530 1421.890 1057.710 1423.070 ;
        RECT 1054.930 1420.290 1056.110 1421.470 ;
        RECT 1056.530 1420.290 1057.710 1421.470 ;
        RECT 1054.930 1241.890 1056.110 1243.070 ;
        RECT 1056.530 1241.890 1057.710 1243.070 ;
        RECT 1054.930 1240.290 1056.110 1241.470 ;
        RECT 1056.530 1240.290 1057.710 1241.470 ;
        RECT 1054.930 1061.890 1056.110 1063.070 ;
        RECT 1056.530 1061.890 1057.710 1063.070 ;
        RECT 1054.930 1060.290 1056.110 1061.470 ;
        RECT 1056.530 1060.290 1057.710 1061.470 ;
        RECT 1234.930 3556.610 1236.110 3557.790 ;
        RECT 1236.530 3556.610 1237.710 3557.790 ;
        RECT 1234.930 3555.010 1236.110 3556.190 ;
        RECT 1236.530 3555.010 1237.710 3556.190 ;
        RECT 1234.930 3401.890 1236.110 3403.070 ;
        RECT 1236.530 3401.890 1237.710 3403.070 ;
        RECT 1234.930 3400.290 1236.110 3401.470 ;
        RECT 1236.530 3400.290 1237.710 3401.470 ;
        RECT 1234.930 3221.890 1236.110 3223.070 ;
        RECT 1236.530 3221.890 1237.710 3223.070 ;
        RECT 1234.930 3220.290 1236.110 3221.470 ;
        RECT 1236.530 3220.290 1237.710 3221.470 ;
        RECT 1234.930 3041.890 1236.110 3043.070 ;
        RECT 1236.530 3041.890 1237.710 3043.070 ;
        RECT 1234.930 3040.290 1236.110 3041.470 ;
        RECT 1236.530 3040.290 1237.710 3041.470 ;
        RECT 1234.930 2861.890 1236.110 2863.070 ;
        RECT 1236.530 2861.890 1237.710 2863.070 ;
        RECT 1234.930 2860.290 1236.110 2861.470 ;
        RECT 1236.530 2860.290 1237.710 2861.470 ;
        RECT 1234.930 2681.890 1236.110 2683.070 ;
        RECT 1236.530 2681.890 1237.710 2683.070 ;
        RECT 1234.930 2680.290 1236.110 2681.470 ;
        RECT 1236.530 2680.290 1237.710 2681.470 ;
        RECT 1234.930 2501.890 1236.110 2503.070 ;
        RECT 1236.530 2501.890 1237.710 2503.070 ;
        RECT 1234.930 2500.290 1236.110 2501.470 ;
        RECT 1236.530 2500.290 1237.710 2501.470 ;
        RECT 1234.930 2321.890 1236.110 2323.070 ;
        RECT 1236.530 2321.890 1237.710 2323.070 ;
        RECT 1234.930 2320.290 1236.110 2321.470 ;
        RECT 1236.530 2320.290 1237.710 2321.470 ;
        RECT 1234.930 2141.890 1236.110 2143.070 ;
        RECT 1236.530 2141.890 1237.710 2143.070 ;
        RECT 1234.930 2140.290 1236.110 2141.470 ;
        RECT 1236.530 2140.290 1237.710 2141.470 ;
        RECT 1234.930 1961.890 1236.110 1963.070 ;
        RECT 1236.530 1961.890 1237.710 1963.070 ;
        RECT 1234.930 1960.290 1236.110 1961.470 ;
        RECT 1236.530 1960.290 1237.710 1961.470 ;
        RECT 1234.930 1781.890 1236.110 1783.070 ;
        RECT 1236.530 1781.890 1237.710 1783.070 ;
        RECT 1234.930 1780.290 1236.110 1781.470 ;
        RECT 1236.530 1780.290 1237.710 1781.470 ;
        RECT 1234.930 1601.890 1236.110 1603.070 ;
        RECT 1236.530 1601.890 1237.710 1603.070 ;
        RECT 1234.930 1600.290 1236.110 1601.470 ;
        RECT 1236.530 1600.290 1237.710 1601.470 ;
        RECT 1234.930 1421.890 1236.110 1423.070 ;
        RECT 1236.530 1421.890 1237.710 1423.070 ;
        RECT 1234.930 1420.290 1236.110 1421.470 ;
        RECT 1236.530 1420.290 1237.710 1421.470 ;
        RECT 1234.930 1241.890 1236.110 1243.070 ;
        RECT 1236.530 1241.890 1237.710 1243.070 ;
        RECT 1234.930 1240.290 1236.110 1241.470 ;
        RECT 1236.530 1240.290 1237.710 1241.470 ;
        RECT 1234.930 1061.890 1236.110 1063.070 ;
        RECT 1236.530 1061.890 1237.710 1063.070 ;
        RECT 1234.930 1060.290 1236.110 1061.470 ;
        RECT 1236.530 1060.290 1237.710 1061.470 ;
        RECT 154.930 881.890 156.110 883.070 ;
        RECT 156.530 881.890 157.710 883.070 ;
        RECT 154.930 880.290 156.110 881.470 ;
        RECT 156.530 880.290 157.710 881.470 ;
        RECT 154.930 701.890 156.110 703.070 ;
        RECT 156.530 701.890 157.710 703.070 ;
        RECT 154.930 700.290 156.110 701.470 ;
        RECT 156.530 700.290 157.710 701.470 ;
        RECT 154.930 521.890 156.110 523.070 ;
        RECT 156.530 521.890 157.710 523.070 ;
        RECT 154.930 520.290 156.110 521.470 ;
        RECT 156.530 520.290 157.710 521.470 ;
        RECT 1234.930 881.890 1236.110 883.070 ;
        RECT 1236.530 881.890 1237.710 883.070 ;
        RECT 1234.930 880.290 1236.110 881.470 ;
        RECT 1236.530 880.290 1237.710 881.470 ;
        RECT 1234.930 701.890 1236.110 703.070 ;
        RECT 1236.530 701.890 1237.710 703.070 ;
        RECT 1234.930 700.290 1236.110 701.470 ;
        RECT 1236.530 700.290 1237.710 701.470 ;
        RECT 1234.930 521.890 1236.110 523.070 ;
        RECT 1236.530 521.890 1237.710 523.070 ;
        RECT 1234.930 520.290 1236.110 521.470 ;
        RECT 1236.530 520.290 1237.710 521.470 ;
        RECT 154.930 341.890 156.110 343.070 ;
        RECT 156.530 341.890 157.710 343.070 ;
        RECT 154.930 340.290 156.110 341.470 ;
        RECT 156.530 340.290 157.710 341.470 ;
        RECT 154.930 161.890 156.110 163.070 ;
        RECT 156.530 161.890 157.710 163.070 ;
        RECT 154.930 160.290 156.110 161.470 ;
        RECT 156.530 160.290 157.710 161.470 ;
        RECT 154.930 -36.510 156.110 -35.330 ;
        RECT 156.530 -36.510 157.710 -35.330 ;
        RECT 154.930 -38.110 156.110 -36.930 ;
        RECT 156.530 -38.110 157.710 -36.930 ;
        RECT 334.930 341.890 336.110 343.070 ;
        RECT 336.530 341.890 337.710 343.070 ;
        RECT 334.930 340.290 336.110 341.470 ;
        RECT 336.530 340.290 337.710 341.470 ;
        RECT 334.930 161.890 336.110 163.070 ;
        RECT 336.530 161.890 337.710 163.070 ;
        RECT 334.930 160.290 336.110 161.470 ;
        RECT 336.530 160.290 337.710 161.470 ;
        RECT 334.930 -36.510 336.110 -35.330 ;
        RECT 336.530 -36.510 337.710 -35.330 ;
        RECT 334.930 -38.110 336.110 -36.930 ;
        RECT 336.530 -38.110 337.710 -36.930 ;
        RECT 514.930 341.890 516.110 343.070 ;
        RECT 516.530 341.890 517.710 343.070 ;
        RECT 514.930 340.290 516.110 341.470 ;
        RECT 516.530 340.290 517.710 341.470 ;
        RECT 514.930 161.890 516.110 163.070 ;
        RECT 516.530 161.890 517.710 163.070 ;
        RECT 514.930 160.290 516.110 161.470 ;
        RECT 516.530 160.290 517.710 161.470 ;
        RECT 514.930 -36.510 516.110 -35.330 ;
        RECT 516.530 -36.510 517.710 -35.330 ;
        RECT 514.930 -38.110 516.110 -36.930 ;
        RECT 516.530 -38.110 517.710 -36.930 ;
        RECT 694.930 341.890 696.110 343.070 ;
        RECT 696.530 341.890 697.710 343.070 ;
        RECT 694.930 340.290 696.110 341.470 ;
        RECT 696.530 340.290 697.710 341.470 ;
        RECT 694.930 161.890 696.110 163.070 ;
        RECT 696.530 161.890 697.710 163.070 ;
        RECT 694.930 160.290 696.110 161.470 ;
        RECT 696.530 160.290 697.710 161.470 ;
        RECT 694.930 -36.510 696.110 -35.330 ;
        RECT 696.530 -36.510 697.710 -35.330 ;
        RECT 694.930 -38.110 696.110 -36.930 ;
        RECT 696.530 -38.110 697.710 -36.930 ;
        RECT 874.930 341.890 876.110 343.070 ;
        RECT 876.530 341.890 877.710 343.070 ;
        RECT 874.930 340.290 876.110 341.470 ;
        RECT 876.530 340.290 877.710 341.470 ;
        RECT 874.930 161.890 876.110 163.070 ;
        RECT 876.530 161.890 877.710 163.070 ;
        RECT 874.930 160.290 876.110 161.470 ;
        RECT 876.530 160.290 877.710 161.470 ;
        RECT 874.930 -36.510 876.110 -35.330 ;
        RECT 876.530 -36.510 877.710 -35.330 ;
        RECT 874.930 -38.110 876.110 -36.930 ;
        RECT 876.530 -38.110 877.710 -36.930 ;
        RECT 1054.930 341.890 1056.110 343.070 ;
        RECT 1056.530 341.890 1057.710 343.070 ;
        RECT 1054.930 340.290 1056.110 341.470 ;
        RECT 1056.530 340.290 1057.710 341.470 ;
        RECT 1054.930 161.890 1056.110 163.070 ;
        RECT 1056.530 161.890 1057.710 163.070 ;
        RECT 1054.930 160.290 1056.110 161.470 ;
        RECT 1056.530 160.290 1057.710 161.470 ;
        RECT 1054.930 -36.510 1056.110 -35.330 ;
        RECT 1056.530 -36.510 1057.710 -35.330 ;
        RECT 1054.930 -38.110 1056.110 -36.930 ;
        RECT 1056.530 -38.110 1057.710 -36.930 ;
        RECT 1234.930 341.890 1236.110 343.070 ;
        RECT 1236.530 341.890 1237.710 343.070 ;
        RECT 1234.930 340.290 1236.110 341.470 ;
        RECT 1236.530 340.290 1237.710 341.470 ;
        RECT 1234.930 161.890 1236.110 163.070 ;
        RECT 1236.530 161.890 1237.710 163.070 ;
        RECT 1234.930 160.290 1236.110 161.470 ;
        RECT 1236.530 160.290 1237.710 161.470 ;
        RECT 1234.930 -36.510 1236.110 -35.330 ;
        RECT 1236.530 -36.510 1237.710 -35.330 ;
        RECT 1234.930 -38.110 1236.110 -36.930 ;
        RECT 1236.530 -38.110 1237.710 -36.930 ;
        RECT 1414.930 3556.610 1416.110 3557.790 ;
        RECT 1416.530 3556.610 1417.710 3557.790 ;
        RECT 1414.930 3555.010 1416.110 3556.190 ;
        RECT 1416.530 3555.010 1417.710 3556.190 ;
        RECT 1414.930 3401.890 1416.110 3403.070 ;
        RECT 1416.530 3401.890 1417.710 3403.070 ;
        RECT 1414.930 3400.290 1416.110 3401.470 ;
        RECT 1416.530 3400.290 1417.710 3401.470 ;
        RECT 1414.930 3221.890 1416.110 3223.070 ;
        RECT 1416.530 3221.890 1417.710 3223.070 ;
        RECT 1414.930 3220.290 1416.110 3221.470 ;
        RECT 1416.530 3220.290 1417.710 3221.470 ;
        RECT 1414.930 3041.890 1416.110 3043.070 ;
        RECT 1416.530 3041.890 1417.710 3043.070 ;
        RECT 1414.930 3040.290 1416.110 3041.470 ;
        RECT 1416.530 3040.290 1417.710 3041.470 ;
        RECT 1414.930 2861.890 1416.110 2863.070 ;
        RECT 1416.530 2861.890 1417.710 2863.070 ;
        RECT 1414.930 2860.290 1416.110 2861.470 ;
        RECT 1416.530 2860.290 1417.710 2861.470 ;
        RECT 1414.930 2681.890 1416.110 2683.070 ;
        RECT 1416.530 2681.890 1417.710 2683.070 ;
        RECT 1414.930 2680.290 1416.110 2681.470 ;
        RECT 1416.530 2680.290 1417.710 2681.470 ;
        RECT 1414.930 2501.890 1416.110 2503.070 ;
        RECT 1416.530 2501.890 1417.710 2503.070 ;
        RECT 1414.930 2500.290 1416.110 2501.470 ;
        RECT 1416.530 2500.290 1417.710 2501.470 ;
        RECT 1414.930 2321.890 1416.110 2323.070 ;
        RECT 1416.530 2321.890 1417.710 2323.070 ;
        RECT 1414.930 2320.290 1416.110 2321.470 ;
        RECT 1416.530 2320.290 1417.710 2321.470 ;
        RECT 1414.930 2141.890 1416.110 2143.070 ;
        RECT 1416.530 2141.890 1417.710 2143.070 ;
        RECT 1414.930 2140.290 1416.110 2141.470 ;
        RECT 1416.530 2140.290 1417.710 2141.470 ;
        RECT 1414.930 1961.890 1416.110 1963.070 ;
        RECT 1416.530 1961.890 1417.710 1963.070 ;
        RECT 1414.930 1960.290 1416.110 1961.470 ;
        RECT 1416.530 1960.290 1417.710 1961.470 ;
        RECT 1414.930 1781.890 1416.110 1783.070 ;
        RECT 1416.530 1781.890 1417.710 1783.070 ;
        RECT 1414.930 1780.290 1416.110 1781.470 ;
        RECT 1416.530 1780.290 1417.710 1781.470 ;
        RECT 1414.930 1601.890 1416.110 1603.070 ;
        RECT 1416.530 1601.890 1417.710 1603.070 ;
        RECT 1414.930 1600.290 1416.110 1601.470 ;
        RECT 1416.530 1600.290 1417.710 1601.470 ;
        RECT 1414.930 1421.890 1416.110 1423.070 ;
        RECT 1416.530 1421.890 1417.710 1423.070 ;
        RECT 1414.930 1420.290 1416.110 1421.470 ;
        RECT 1416.530 1420.290 1417.710 1421.470 ;
        RECT 1414.930 1241.890 1416.110 1243.070 ;
        RECT 1416.530 1241.890 1417.710 1243.070 ;
        RECT 1414.930 1240.290 1416.110 1241.470 ;
        RECT 1416.530 1240.290 1417.710 1241.470 ;
        RECT 1414.930 1061.890 1416.110 1063.070 ;
        RECT 1416.530 1061.890 1417.710 1063.070 ;
        RECT 1414.930 1060.290 1416.110 1061.470 ;
        RECT 1416.530 1060.290 1417.710 1061.470 ;
        RECT 1414.930 881.890 1416.110 883.070 ;
        RECT 1416.530 881.890 1417.710 883.070 ;
        RECT 1414.930 880.290 1416.110 881.470 ;
        RECT 1416.530 880.290 1417.710 881.470 ;
        RECT 1414.930 701.890 1416.110 703.070 ;
        RECT 1416.530 701.890 1417.710 703.070 ;
        RECT 1414.930 700.290 1416.110 701.470 ;
        RECT 1416.530 700.290 1417.710 701.470 ;
        RECT 1414.930 521.890 1416.110 523.070 ;
        RECT 1416.530 521.890 1417.710 523.070 ;
        RECT 1414.930 520.290 1416.110 521.470 ;
        RECT 1416.530 520.290 1417.710 521.470 ;
        RECT 1414.930 341.890 1416.110 343.070 ;
        RECT 1416.530 341.890 1417.710 343.070 ;
        RECT 1414.930 340.290 1416.110 341.470 ;
        RECT 1416.530 340.290 1417.710 341.470 ;
        RECT 1414.930 161.890 1416.110 163.070 ;
        RECT 1416.530 161.890 1417.710 163.070 ;
        RECT 1414.930 160.290 1416.110 161.470 ;
        RECT 1416.530 160.290 1417.710 161.470 ;
        RECT 1414.930 -36.510 1416.110 -35.330 ;
        RECT 1416.530 -36.510 1417.710 -35.330 ;
        RECT 1414.930 -38.110 1416.110 -36.930 ;
        RECT 1416.530 -38.110 1417.710 -36.930 ;
        RECT 1594.930 3556.610 1596.110 3557.790 ;
        RECT 1596.530 3556.610 1597.710 3557.790 ;
        RECT 1594.930 3555.010 1596.110 3556.190 ;
        RECT 1596.530 3555.010 1597.710 3556.190 ;
        RECT 1594.930 3401.890 1596.110 3403.070 ;
        RECT 1596.530 3401.890 1597.710 3403.070 ;
        RECT 1594.930 3400.290 1596.110 3401.470 ;
        RECT 1596.530 3400.290 1597.710 3401.470 ;
        RECT 1594.930 3221.890 1596.110 3223.070 ;
        RECT 1596.530 3221.890 1597.710 3223.070 ;
        RECT 1594.930 3220.290 1596.110 3221.470 ;
        RECT 1596.530 3220.290 1597.710 3221.470 ;
        RECT 1594.930 3041.890 1596.110 3043.070 ;
        RECT 1596.530 3041.890 1597.710 3043.070 ;
        RECT 1594.930 3040.290 1596.110 3041.470 ;
        RECT 1596.530 3040.290 1597.710 3041.470 ;
        RECT 1594.930 2861.890 1596.110 2863.070 ;
        RECT 1596.530 2861.890 1597.710 2863.070 ;
        RECT 1594.930 2860.290 1596.110 2861.470 ;
        RECT 1596.530 2860.290 1597.710 2861.470 ;
        RECT 1594.930 2681.890 1596.110 2683.070 ;
        RECT 1596.530 2681.890 1597.710 2683.070 ;
        RECT 1594.930 2680.290 1596.110 2681.470 ;
        RECT 1596.530 2680.290 1597.710 2681.470 ;
        RECT 1594.930 2501.890 1596.110 2503.070 ;
        RECT 1596.530 2501.890 1597.710 2503.070 ;
        RECT 1594.930 2500.290 1596.110 2501.470 ;
        RECT 1596.530 2500.290 1597.710 2501.470 ;
        RECT 1594.930 2321.890 1596.110 2323.070 ;
        RECT 1596.530 2321.890 1597.710 2323.070 ;
        RECT 1594.930 2320.290 1596.110 2321.470 ;
        RECT 1596.530 2320.290 1597.710 2321.470 ;
        RECT 1594.930 2141.890 1596.110 2143.070 ;
        RECT 1596.530 2141.890 1597.710 2143.070 ;
        RECT 1594.930 2140.290 1596.110 2141.470 ;
        RECT 1596.530 2140.290 1597.710 2141.470 ;
        RECT 1594.930 1961.890 1596.110 1963.070 ;
        RECT 1596.530 1961.890 1597.710 1963.070 ;
        RECT 1594.930 1960.290 1596.110 1961.470 ;
        RECT 1596.530 1960.290 1597.710 1961.470 ;
        RECT 1594.930 1781.890 1596.110 1783.070 ;
        RECT 1596.530 1781.890 1597.710 1783.070 ;
        RECT 1594.930 1780.290 1596.110 1781.470 ;
        RECT 1596.530 1780.290 1597.710 1781.470 ;
        RECT 1594.930 1601.890 1596.110 1603.070 ;
        RECT 1596.530 1601.890 1597.710 1603.070 ;
        RECT 1594.930 1600.290 1596.110 1601.470 ;
        RECT 1596.530 1600.290 1597.710 1601.470 ;
        RECT 1594.930 1421.890 1596.110 1423.070 ;
        RECT 1596.530 1421.890 1597.710 1423.070 ;
        RECT 1594.930 1420.290 1596.110 1421.470 ;
        RECT 1596.530 1420.290 1597.710 1421.470 ;
        RECT 1594.930 1241.890 1596.110 1243.070 ;
        RECT 1596.530 1241.890 1597.710 1243.070 ;
        RECT 1594.930 1240.290 1596.110 1241.470 ;
        RECT 1596.530 1240.290 1597.710 1241.470 ;
        RECT 1594.930 1061.890 1596.110 1063.070 ;
        RECT 1596.530 1061.890 1597.710 1063.070 ;
        RECT 1594.930 1060.290 1596.110 1061.470 ;
        RECT 1596.530 1060.290 1597.710 1061.470 ;
        RECT 1594.930 881.890 1596.110 883.070 ;
        RECT 1596.530 881.890 1597.710 883.070 ;
        RECT 1594.930 880.290 1596.110 881.470 ;
        RECT 1596.530 880.290 1597.710 881.470 ;
        RECT 1594.930 701.890 1596.110 703.070 ;
        RECT 1596.530 701.890 1597.710 703.070 ;
        RECT 1594.930 700.290 1596.110 701.470 ;
        RECT 1596.530 700.290 1597.710 701.470 ;
        RECT 1594.930 521.890 1596.110 523.070 ;
        RECT 1596.530 521.890 1597.710 523.070 ;
        RECT 1594.930 520.290 1596.110 521.470 ;
        RECT 1596.530 520.290 1597.710 521.470 ;
        RECT 1594.930 341.890 1596.110 343.070 ;
        RECT 1596.530 341.890 1597.710 343.070 ;
        RECT 1594.930 340.290 1596.110 341.470 ;
        RECT 1596.530 340.290 1597.710 341.470 ;
        RECT 1594.930 161.890 1596.110 163.070 ;
        RECT 1596.530 161.890 1597.710 163.070 ;
        RECT 1594.930 160.290 1596.110 161.470 ;
        RECT 1596.530 160.290 1597.710 161.470 ;
        RECT 1594.930 -36.510 1596.110 -35.330 ;
        RECT 1596.530 -36.510 1597.710 -35.330 ;
        RECT 1594.930 -38.110 1596.110 -36.930 ;
        RECT 1596.530 -38.110 1597.710 -36.930 ;
        RECT 1774.930 3556.610 1776.110 3557.790 ;
        RECT 1776.530 3556.610 1777.710 3557.790 ;
        RECT 1774.930 3555.010 1776.110 3556.190 ;
        RECT 1776.530 3555.010 1777.710 3556.190 ;
        RECT 1774.930 3401.890 1776.110 3403.070 ;
        RECT 1776.530 3401.890 1777.710 3403.070 ;
        RECT 1774.930 3400.290 1776.110 3401.470 ;
        RECT 1776.530 3400.290 1777.710 3401.470 ;
        RECT 1774.930 3221.890 1776.110 3223.070 ;
        RECT 1776.530 3221.890 1777.710 3223.070 ;
        RECT 1774.930 3220.290 1776.110 3221.470 ;
        RECT 1776.530 3220.290 1777.710 3221.470 ;
        RECT 1774.930 3041.890 1776.110 3043.070 ;
        RECT 1776.530 3041.890 1777.710 3043.070 ;
        RECT 1774.930 3040.290 1776.110 3041.470 ;
        RECT 1776.530 3040.290 1777.710 3041.470 ;
        RECT 1774.930 2861.890 1776.110 2863.070 ;
        RECT 1776.530 2861.890 1777.710 2863.070 ;
        RECT 1774.930 2860.290 1776.110 2861.470 ;
        RECT 1776.530 2860.290 1777.710 2861.470 ;
        RECT 1774.930 2681.890 1776.110 2683.070 ;
        RECT 1776.530 2681.890 1777.710 2683.070 ;
        RECT 1774.930 2680.290 1776.110 2681.470 ;
        RECT 1776.530 2680.290 1777.710 2681.470 ;
        RECT 1774.930 2501.890 1776.110 2503.070 ;
        RECT 1776.530 2501.890 1777.710 2503.070 ;
        RECT 1774.930 2500.290 1776.110 2501.470 ;
        RECT 1776.530 2500.290 1777.710 2501.470 ;
        RECT 1774.930 2321.890 1776.110 2323.070 ;
        RECT 1776.530 2321.890 1777.710 2323.070 ;
        RECT 1774.930 2320.290 1776.110 2321.470 ;
        RECT 1776.530 2320.290 1777.710 2321.470 ;
        RECT 1774.930 2141.890 1776.110 2143.070 ;
        RECT 1776.530 2141.890 1777.710 2143.070 ;
        RECT 1774.930 2140.290 1776.110 2141.470 ;
        RECT 1776.530 2140.290 1777.710 2141.470 ;
        RECT 1774.930 1961.890 1776.110 1963.070 ;
        RECT 1776.530 1961.890 1777.710 1963.070 ;
        RECT 1774.930 1960.290 1776.110 1961.470 ;
        RECT 1776.530 1960.290 1777.710 1961.470 ;
        RECT 1774.930 1781.890 1776.110 1783.070 ;
        RECT 1776.530 1781.890 1777.710 1783.070 ;
        RECT 1774.930 1780.290 1776.110 1781.470 ;
        RECT 1776.530 1780.290 1777.710 1781.470 ;
        RECT 1774.930 1601.890 1776.110 1603.070 ;
        RECT 1776.530 1601.890 1777.710 1603.070 ;
        RECT 1774.930 1600.290 1776.110 1601.470 ;
        RECT 1776.530 1600.290 1777.710 1601.470 ;
        RECT 1774.930 1421.890 1776.110 1423.070 ;
        RECT 1776.530 1421.890 1777.710 1423.070 ;
        RECT 1774.930 1420.290 1776.110 1421.470 ;
        RECT 1776.530 1420.290 1777.710 1421.470 ;
        RECT 1774.930 1241.890 1776.110 1243.070 ;
        RECT 1776.530 1241.890 1777.710 1243.070 ;
        RECT 1774.930 1240.290 1776.110 1241.470 ;
        RECT 1776.530 1240.290 1777.710 1241.470 ;
        RECT 1774.930 1061.890 1776.110 1063.070 ;
        RECT 1776.530 1061.890 1777.710 1063.070 ;
        RECT 1774.930 1060.290 1776.110 1061.470 ;
        RECT 1776.530 1060.290 1777.710 1061.470 ;
        RECT 1774.930 881.890 1776.110 883.070 ;
        RECT 1776.530 881.890 1777.710 883.070 ;
        RECT 1774.930 880.290 1776.110 881.470 ;
        RECT 1776.530 880.290 1777.710 881.470 ;
        RECT 1774.930 701.890 1776.110 703.070 ;
        RECT 1776.530 701.890 1777.710 703.070 ;
        RECT 1774.930 700.290 1776.110 701.470 ;
        RECT 1776.530 700.290 1777.710 701.470 ;
        RECT 1774.930 521.890 1776.110 523.070 ;
        RECT 1776.530 521.890 1777.710 523.070 ;
        RECT 1774.930 520.290 1776.110 521.470 ;
        RECT 1776.530 520.290 1777.710 521.470 ;
        RECT 1774.930 341.890 1776.110 343.070 ;
        RECT 1776.530 341.890 1777.710 343.070 ;
        RECT 1774.930 340.290 1776.110 341.470 ;
        RECT 1776.530 340.290 1777.710 341.470 ;
        RECT 1774.930 161.890 1776.110 163.070 ;
        RECT 1776.530 161.890 1777.710 163.070 ;
        RECT 1774.930 160.290 1776.110 161.470 ;
        RECT 1776.530 160.290 1777.710 161.470 ;
        RECT 1774.930 -36.510 1776.110 -35.330 ;
        RECT 1776.530 -36.510 1777.710 -35.330 ;
        RECT 1774.930 -38.110 1776.110 -36.930 ;
        RECT 1776.530 -38.110 1777.710 -36.930 ;
        RECT 1954.930 3556.610 1956.110 3557.790 ;
        RECT 1956.530 3556.610 1957.710 3557.790 ;
        RECT 1954.930 3555.010 1956.110 3556.190 ;
        RECT 1956.530 3555.010 1957.710 3556.190 ;
        RECT 1954.930 3401.890 1956.110 3403.070 ;
        RECT 1956.530 3401.890 1957.710 3403.070 ;
        RECT 1954.930 3400.290 1956.110 3401.470 ;
        RECT 1956.530 3400.290 1957.710 3401.470 ;
        RECT 1954.930 3221.890 1956.110 3223.070 ;
        RECT 1956.530 3221.890 1957.710 3223.070 ;
        RECT 1954.930 3220.290 1956.110 3221.470 ;
        RECT 1956.530 3220.290 1957.710 3221.470 ;
        RECT 1954.930 3041.890 1956.110 3043.070 ;
        RECT 1956.530 3041.890 1957.710 3043.070 ;
        RECT 1954.930 3040.290 1956.110 3041.470 ;
        RECT 1956.530 3040.290 1957.710 3041.470 ;
        RECT 1954.930 2861.890 1956.110 2863.070 ;
        RECT 1956.530 2861.890 1957.710 2863.070 ;
        RECT 1954.930 2860.290 1956.110 2861.470 ;
        RECT 1956.530 2860.290 1957.710 2861.470 ;
        RECT 1954.930 2681.890 1956.110 2683.070 ;
        RECT 1956.530 2681.890 1957.710 2683.070 ;
        RECT 1954.930 2680.290 1956.110 2681.470 ;
        RECT 1956.530 2680.290 1957.710 2681.470 ;
        RECT 1954.930 2501.890 1956.110 2503.070 ;
        RECT 1956.530 2501.890 1957.710 2503.070 ;
        RECT 1954.930 2500.290 1956.110 2501.470 ;
        RECT 1956.530 2500.290 1957.710 2501.470 ;
        RECT 1954.930 2321.890 1956.110 2323.070 ;
        RECT 1956.530 2321.890 1957.710 2323.070 ;
        RECT 1954.930 2320.290 1956.110 2321.470 ;
        RECT 1956.530 2320.290 1957.710 2321.470 ;
        RECT 1954.930 2141.890 1956.110 2143.070 ;
        RECT 1956.530 2141.890 1957.710 2143.070 ;
        RECT 1954.930 2140.290 1956.110 2141.470 ;
        RECT 1956.530 2140.290 1957.710 2141.470 ;
        RECT 1954.930 1961.890 1956.110 1963.070 ;
        RECT 1956.530 1961.890 1957.710 1963.070 ;
        RECT 1954.930 1960.290 1956.110 1961.470 ;
        RECT 1956.530 1960.290 1957.710 1961.470 ;
        RECT 1954.930 1781.890 1956.110 1783.070 ;
        RECT 1956.530 1781.890 1957.710 1783.070 ;
        RECT 1954.930 1780.290 1956.110 1781.470 ;
        RECT 1956.530 1780.290 1957.710 1781.470 ;
        RECT 1954.930 1601.890 1956.110 1603.070 ;
        RECT 1956.530 1601.890 1957.710 1603.070 ;
        RECT 1954.930 1600.290 1956.110 1601.470 ;
        RECT 1956.530 1600.290 1957.710 1601.470 ;
        RECT 1954.930 1421.890 1956.110 1423.070 ;
        RECT 1956.530 1421.890 1957.710 1423.070 ;
        RECT 1954.930 1420.290 1956.110 1421.470 ;
        RECT 1956.530 1420.290 1957.710 1421.470 ;
        RECT 1954.930 1241.890 1956.110 1243.070 ;
        RECT 1956.530 1241.890 1957.710 1243.070 ;
        RECT 1954.930 1240.290 1956.110 1241.470 ;
        RECT 1956.530 1240.290 1957.710 1241.470 ;
        RECT 1954.930 1061.890 1956.110 1063.070 ;
        RECT 1956.530 1061.890 1957.710 1063.070 ;
        RECT 1954.930 1060.290 1956.110 1061.470 ;
        RECT 1956.530 1060.290 1957.710 1061.470 ;
        RECT 1954.930 881.890 1956.110 883.070 ;
        RECT 1956.530 881.890 1957.710 883.070 ;
        RECT 1954.930 880.290 1956.110 881.470 ;
        RECT 1956.530 880.290 1957.710 881.470 ;
        RECT 1954.930 701.890 1956.110 703.070 ;
        RECT 1956.530 701.890 1957.710 703.070 ;
        RECT 1954.930 700.290 1956.110 701.470 ;
        RECT 1956.530 700.290 1957.710 701.470 ;
        RECT 1954.930 521.890 1956.110 523.070 ;
        RECT 1956.530 521.890 1957.710 523.070 ;
        RECT 1954.930 520.290 1956.110 521.470 ;
        RECT 1956.530 520.290 1957.710 521.470 ;
        RECT 1954.930 341.890 1956.110 343.070 ;
        RECT 1956.530 341.890 1957.710 343.070 ;
        RECT 1954.930 340.290 1956.110 341.470 ;
        RECT 1956.530 340.290 1957.710 341.470 ;
        RECT 1954.930 161.890 1956.110 163.070 ;
        RECT 1956.530 161.890 1957.710 163.070 ;
        RECT 1954.930 160.290 1956.110 161.470 ;
        RECT 1956.530 160.290 1957.710 161.470 ;
        RECT 1954.930 -36.510 1956.110 -35.330 ;
        RECT 1956.530 -36.510 1957.710 -35.330 ;
        RECT 1954.930 -38.110 1956.110 -36.930 ;
        RECT 1956.530 -38.110 1957.710 -36.930 ;
        RECT 2134.930 3556.610 2136.110 3557.790 ;
        RECT 2136.530 3556.610 2137.710 3557.790 ;
        RECT 2134.930 3555.010 2136.110 3556.190 ;
        RECT 2136.530 3555.010 2137.710 3556.190 ;
        RECT 2134.930 3401.890 2136.110 3403.070 ;
        RECT 2136.530 3401.890 2137.710 3403.070 ;
        RECT 2134.930 3400.290 2136.110 3401.470 ;
        RECT 2136.530 3400.290 2137.710 3401.470 ;
        RECT 2134.930 3221.890 2136.110 3223.070 ;
        RECT 2136.530 3221.890 2137.710 3223.070 ;
        RECT 2134.930 3220.290 2136.110 3221.470 ;
        RECT 2136.530 3220.290 2137.710 3221.470 ;
        RECT 2134.930 3041.890 2136.110 3043.070 ;
        RECT 2136.530 3041.890 2137.710 3043.070 ;
        RECT 2134.930 3040.290 2136.110 3041.470 ;
        RECT 2136.530 3040.290 2137.710 3041.470 ;
        RECT 2134.930 2861.890 2136.110 2863.070 ;
        RECT 2136.530 2861.890 2137.710 2863.070 ;
        RECT 2134.930 2860.290 2136.110 2861.470 ;
        RECT 2136.530 2860.290 2137.710 2861.470 ;
        RECT 2134.930 2681.890 2136.110 2683.070 ;
        RECT 2136.530 2681.890 2137.710 2683.070 ;
        RECT 2134.930 2680.290 2136.110 2681.470 ;
        RECT 2136.530 2680.290 2137.710 2681.470 ;
        RECT 2134.930 2501.890 2136.110 2503.070 ;
        RECT 2136.530 2501.890 2137.710 2503.070 ;
        RECT 2134.930 2500.290 2136.110 2501.470 ;
        RECT 2136.530 2500.290 2137.710 2501.470 ;
        RECT 2134.930 2321.890 2136.110 2323.070 ;
        RECT 2136.530 2321.890 2137.710 2323.070 ;
        RECT 2134.930 2320.290 2136.110 2321.470 ;
        RECT 2136.530 2320.290 2137.710 2321.470 ;
        RECT 2134.930 2141.890 2136.110 2143.070 ;
        RECT 2136.530 2141.890 2137.710 2143.070 ;
        RECT 2134.930 2140.290 2136.110 2141.470 ;
        RECT 2136.530 2140.290 2137.710 2141.470 ;
        RECT 2134.930 1961.890 2136.110 1963.070 ;
        RECT 2136.530 1961.890 2137.710 1963.070 ;
        RECT 2134.930 1960.290 2136.110 1961.470 ;
        RECT 2136.530 1960.290 2137.710 1961.470 ;
        RECT 2134.930 1781.890 2136.110 1783.070 ;
        RECT 2136.530 1781.890 2137.710 1783.070 ;
        RECT 2134.930 1780.290 2136.110 1781.470 ;
        RECT 2136.530 1780.290 2137.710 1781.470 ;
        RECT 2134.930 1601.890 2136.110 1603.070 ;
        RECT 2136.530 1601.890 2137.710 1603.070 ;
        RECT 2134.930 1600.290 2136.110 1601.470 ;
        RECT 2136.530 1600.290 2137.710 1601.470 ;
        RECT 2134.930 1421.890 2136.110 1423.070 ;
        RECT 2136.530 1421.890 2137.710 1423.070 ;
        RECT 2134.930 1420.290 2136.110 1421.470 ;
        RECT 2136.530 1420.290 2137.710 1421.470 ;
        RECT 2134.930 1241.890 2136.110 1243.070 ;
        RECT 2136.530 1241.890 2137.710 1243.070 ;
        RECT 2134.930 1240.290 2136.110 1241.470 ;
        RECT 2136.530 1240.290 2137.710 1241.470 ;
        RECT 2134.930 1061.890 2136.110 1063.070 ;
        RECT 2136.530 1061.890 2137.710 1063.070 ;
        RECT 2134.930 1060.290 2136.110 1061.470 ;
        RECT 2136.530 1060.290 2137.710 1061.470 ;
        RECT 2134.930 881.890 2136.110 883.070 ;
        RECT 2136.530 881.890 2137.710 883.070 ;
        RECT 2134.930 880.290 2136.110 881.470 ;
        RECT 2136.530 880.290 2137.710 881.470 ;
        RECT 2134.930 701.890 2136.110 703.070 ;
        RECT 2136.530 701.890 2137.710 703.070 ;
        RECT 2134.930 700.290 2136.110 701.470 ;
        RECT 2136.530 700.290 2137.710 701.470 ;
        RECT 2134.930 521.890 2136.110 523.070 ;
        RECT 2136.530 521.890 2137.710 523.070 ;
        RECT 2134.930 520.290 2136.110 521.470 ;
        RECT 2136.530 520.290 2137.710 521.470 ;
        RECT 2134.930 341.890 2136.110 343.070 ;
        RECT 2136.530 341.890 2137.710 343.070 ;
        RECT 2134.930 340.290 2136.110 341.470 ;
        RECT 2136.530 340.290 2137.710 341.470 ;
        RECT 2134.930 161.890 2136.110 163.070 ;
        RECT 2136.530 161.890 2137.710 163.070 ;
        RECT 2134.930 160.290 2136.110 161.470 ;
        RECT 2136.530 160.290 2137.710 161.470 ;
        RECT 2134.930 -36.510 2136.110 -35.330 ;
        RECT 2136.530 -36.510 2137.710 -35.330 ;
        RECT 2134.930 -38.110 2136.110 -36.930 ;
        RECT 2136.530 -38.110 2137.710 -36.930 ;
        RECT 2314.930 3556.610 2316.110 3557.790 ;
        RECT 2316.530 3556.610 2317.710 3557.790 ;
        RECT 2314.930 3555.010 2316.110 3556.190 ;
        RECT 2316.530 3555.010 2317.710 3556.190 ;
        RECT 2314.930 3401.890 2316.110 3403.070 ;
        RECT 2316.530 3401.890 2317.710 3403.070 ;
        RECT 2314.930 3400.290 2316.110 3401.470 ;
        RECT 2316.530 3400.290 2317.710 3401.470 ;
        RECT 2314.930 3221.890 2316.110 3223.070 ;
        RECT 2316.530 3221.890 2317.710 3223.070 ;
        RECT 2314.930 3220.290 2316.110 3221.470 ;
        RECT 2316.530 3220.290 2317.710 3221.470 ;
        RECT 2314.930 3041.890 2316.110 3043.070 ;
        RECT 2316.530 3041.890 2317.710 3043.070 ;
        RECT 2314.930 3040.290 2316.110 3041.470 ;
        RECT 2316.530 3040.290 2317.710 3041.470 ;
        RECT 2314.930 2861.890 2316.110 2863.070 ;
        RECT 2316.530 2861.890 2317.710 2863.070 ;
        RECT 2314.930 2860.290 2316.110 2861.470 ;
        RECT 2316.530 2860.290 2317.710 2861.470 ;
        RECT 2314.930 2681.890 2316.110 2683.070 ;
        RECT 2316.530 2681.890 2317.710 2683.070 ;
        RECT 2314.930 2680.290 2316.110 2681.470 ;
        RECT 2316.530 2680.290 2317.710 2681.470 ;
        RECT 2314.930 2501.890 2316.110 2503.070 ;
        RECT 2316.530 2501.890 2317.710 2503.070 ;
        RECT 2314.930 2500.290 2316.110 2501.470 ;
        RECT 2316.530 2500.290 2317.710 2501.470 ;
        RECT 2314.930 2321.890 2316.110 2323.070 ;
        RECT 2316.530 2321.890 2317.710 2323.070 ;
        RECT 2314.930 2320.290 2316.110 2321.470 ;
        RECT 2316.530 2320.290 2317.710 2321.470 ;
        RECT 2314.930 2141.890 2316.110 2143.070 ;
        RECT 2316.530 2141.890 2317.710 2143.070 ;
        RECT 2314.930 2140.290 2316.110 2141.470 ;
        RECT 2316.530 2140.290 2317.710 2141.470 ;
        RECT 2314.930 1961.890 2316.110 1963.070 ;
        RECT 2316.530 1961.890 2317.710 1963.070 ;
        RECT 2314.930 1960.290 2316.110 1961.470 ;
        RECT 2316.530 1960.290 2317.710 1961.470 ;
        RECT 2314.930 1781.890 2316.110 1783.070 ;
        RECT 2316.530 1781.890 2317.710 1783.070 ;
        RECT 2314.930 1780.290 2316.110 1781.470 ;
        RECT 2316.530 1780.290 2317.710 1781.470 ;
        RECT 2314.930 1601.890 2316.110 1603.070 ;
        RECT 2316.530 1601.890 2317.710 1603.070 ;
        RECT 2314.930 1600.290 2316.110 1601.470 ;
        RECT 2316.530 1600.290 2317.710 1601.470 ;
        RECT 2314.930 1421.890 2316.110 1423.070 ;
        RECT 2316.530 1421.890 2317.710 1423.070 ;
        RECT 2314.930 1420.290 2316.110 1421.470 ;
        RECT 2316.530 1420.290 2317.710 1421.470 ;
        RECT 2314.930 1241.890 2316.110 1243.070 ;
        RECT 2316.530 1241.890 2317.710 1243.070 ;
        RECT 2314.930 1240.290 2316.110 1241.470 ;
        RECT 2316.530 1240.290 2317.710 1241.470 ;
        RECT 2314.930 1061.890 2316.110 1063.070 ;
        RECT 2316.530 1061.890 2317.710 1063.070 ;
        RECT 2314.930 1060.290 2316.110 1061.470 ;
        RECT 2316.530 1060.290 2317.710 1061.470 ;
        RECT 2314.930 881.890 2316.110 883.070 ;
        RECT 2316.530 881.890 2317.710 883.070 ;
        RECT 2314.930 880.290 2316.110 881.470 ;
        RECT 2316.530 880.290 2317.710 881.470 ;
        RECT 2314.930 701.890 2316.110 703.070 ;
        RECT 2316.530 701.890 2317.710 703.070 ;
        RECT 2314.930 700.290 2316.110 701.470 ;
        RECT 2316.530 700.290 2317.710 701.470 ;
        RECT 2314.930 521.890 2316.110 523.070 ;
        RECT 2316.530 521.890 2317.710 523.070 ;
        RECT 2314.930 520.290 2316.110 521.470 ;
        RECT 2316.530 520.290 2317.710 521.470 ;
        RECT 2314.930 341.890 2316.110 343.070 ;
        RECT 2316.530 341.890 2317.710 343.070 ;
        RECT 2314.930 340.290 2316.110 341.470 ;
        RECT 2316.530 340.290 2317.710 341.470 ;
        RECT 2314.930 161.890 2316.110 163.070 ;
        RECT 2316.530 161.890 2317.710 163.070 ;
        RECT 2314.930 160.290 2316.110 161.470 ;
        RECT 2316.530 160.290 2317.710 161.470 ;
        RECT 2314.930 -36.510 2316.110 -35.330 ;
        RECT 2316.530 -36.510 2317.710 -35.330 ;
        RECT 2314.930 -38.110 2316.110 -36.930 ;
        RECT 2316.530 -38.110 2317.710 -36.930 ;
        RECT 2494.930 3556.610 2496.110 3557.790 ;
        RECT 2496.530 3556.610 2497.710 3557.790 ;
        RECT 2494.930 3555.010 2496.110 3556.190 ;
        RECT 2496.530 3555.010 2497.710 3556.190 ;
        RECT 2494.930 3401.890 2496.110 3403.070 ;
        RECT 2496.530 3401.890 2497.710 3403.070 ;
        RECT 2494.930 3400.290 2496.110 3401.470 ;
        RECT 2496.530 3400.290 2497.710 3401.470 ;
        RECT 2494.930 3221.890 2496.110 3223.070 ;
        RECT 2496.530 3221.890 2497.710 3223.070 ;
        RECT 2494.930 3220.290 2496.110 3221.470 ;
        RECT 2496.530 3220.290 2497.710 3221.470 ;
        RECT 2494.930 3041.890 2496.110 3043.070 ;
        RECT 2496.530 3041.890 2497.710 3043.070 ;
        RECT 2494.930 3040.290 2496.110 3041.470 ;
        RECT 2496.530 3040.290 2497.710 3041.470 ;
        RECT 2494.930 2861.890 2496.110 2863.070 ;
        RECT 2496.530 2861.890 2497.710 2863.070 ;
        RECT 2494.930 2860.290 2496.110 2861.470 ;
        RECT 2496.530 2860.290 2497.710 2861.470 ;
        RECT 2494.930 2681.890 2496.110 2683.070 ;
        RECT 2496.530 2681.890 2497.710 2683.070 ;
        RECT 2494.930 2680.290 2496.110 2681.470 ;
        RECT 2496.530 2680.290 2497.710 2681.470 ;
        RECT 2494.930 2501.890 2496.110 2503.070 ;
        RECT 2496.530 2501.890 2497.710 2503.070 ;
        RECT 2494.930 2500.290 2496.110 2501.470 ;
        RECT 2496.530 2500.290 2497.710 2501.470 ;
        RECT 2494.930 2321.890 2496.110 2323.070 ;
        RECT 2496.530 2321.890 2497.710 2323.070 ;
        RECT 2494.930 2320.290 2496.110 2321.470 ;
        RECT 2496.530 2320.290 2497.710 2321.470 ;
        RECT 2494.930 2141.890 2496.110 2143.070 ;
        RECT 2496.530 2141.890 2497.710 2143.070 ;
        RECT 2494.930 2140.290 2496.110 2141.470 ;
        RECT 2496.530 2140.290 2497.710 2141.470 ;
        RECT 2494.930 1961.890 2496.110 1963.070 ;
        RECT 2496.530 1961.890 2497.710 1963.070 ;
        RECT 2494.930 1960.290 2496.110 1961.470 ;
        RECT 2496.530 1960.290 2497.710 1961.470 ;
        RECT 2494.930 1781.890 2496.110 1783.070 ;
        RECT 2496.530 1781.890 2497.710 1783.070 ;
        RECT 2494.930 1780.290 2496.110 1781.470 ;
        RECT 2496.530 1780.290 2497.710 1781.470 ;
        RECT 2494.930 1601.890 2496.110 1603.070 ;
        RECT 2496.530 1601.890 2497.710 1603.070 ;
        RECT 2494.930 1600.290 2496.110 1601.470 ;
        RECT 2496.530 1600.290 2497.710 1601.470 ;
        RECT 2494.930 1421.890 2496.110 1423.070 ;
        RECT 2496.530 1421.890 2497.710 1423.070 ;
        RECT 2494.930 1420.290 2496.110 1421.470 ;
        RECT 2496.530 1420.290 2497.710 1421.470 ;
        RECT 2494.930 1241.890 2496.110 1243.070 ;
        RECT 2496.530 1241.890 2497.710 1243.070 ;
        RECT 2494.930 1240.290 2496.110 1241.470 ;
        RECT 2496.530 1240.290 2497.710 1241.470 ;
        RECT 2494.930 1061.890 2496.110 1063.070 ;
        RECT 2496.530 1061.890 2497.710 1063.070 ;
        RECT 2494.930 1060.290 2496.110 1061.470 ;
        RECT 2496.530 1060.290 2497.710 1061.470 ;
        RECT 2494.930 881.890 2496.110 883.070 ;
        RECT 2496.530 881.890 2497.710 883.070 ;
        RECT 2494.930 880.290 2496.110 881.470 ;
        RECT 2496.530 880.290 2497.710 881.470 ;
        RECT 2494.930 701.890 2496.110 703.070 ;
        RECT 2496.530 701.890 2497.710 703.070 ;
        RECT 2494.930 700.290 2496.110 701.470 ;
        RECT 2496.530 700.290 2497.710 701.470 ;
        RECT 2494.930 521.890 2496.110 523.070 ;
        RECT 2496.530 521.890 2497.710 523.070 ;
        RECT 2494.930 520.290 2496.110 521.470 ;
        RECT 2496.530 520.290 2497.710 521.470 ;
        RECT 2494.930 341.890 2496.110 343.070 ;
        RECT 2496.530 341.890 2497.710 343.070 ;
        RECT 2494.930 340.290 2496.110 341.470 ;
        RECT 2496.530 340.290 2497.710 341.470 ;
        RECT 2494.930 161.890 2496.110 163.070 ;
        RECT 2496.530 161.890 2497.710 163.070 ;
        RECT 2494.930 160.290 2496.110 161.470 ;
        RECT 2496.530 160.290 2497.710 161.470 ;
        RECT 2494.930 -36.510 2496.110 -35.330 ;
        RECT 2496.530 -36.510 2497.710 -35.330 ;
        RECT 2494.930 -38.110 2496.110 -36.930 ;
        RECT 2496.530 -38.110 2497.710 -36.930 ;
        RECT 2674.930 3556.610 2676.110 3557.790 ;
        RECT 2676.530 3556.610 2677.710 3557.790 ;
        RECT 2674.930 3555.010 2676.110 3556.190 ;
        RECT 2676.530 3555.010 2677.710 3556.190 ;
        RECT 2674.930 3401.890 2676.110 3403.070 ;
        RECT 2676.530 3401.890 2677.710 3403.070 ;
        RECT 2674.930 3400.290 2676.110 3401.470 ;
        RECT 2676.530 3400.290 2677.710 3401.470 ;
        RECT 2674.930 3221.890 2676.110 3223.070 ;
        RECT 2676.530 3221.890 2677.710 3223.070 ;
        RECT 2674.930 3220.290 2676.110 3221.470 ;
        RECT 2676.530 3220.290 2677.710 3221.470 ;
        RECT 2674.930 3041.890 2676.110 3043.070 ;
        RECT 2676.530 3041.890 2677.710 3043.070 ;
        RECT 2674.930 3040.290 2676.110 3041.470 ;
        RECT 2676.530 3040.290 2677.710 3041.470 ;
        RECT 2674.930 2861.890 2676.110 2863.070 ;
        RECT 2676.530 2861.890 2677.710 2863.070 ;
        RECT 2674.930 2860.290 2676.110 2861.470 ;
        RECT 2676.530 2860.290 2677.710 2861.470 ;
        RECT 2674.930 2681.890 2676.110 2683.070 ;
        RECT 2676.530 2681.890 2677.710 2683.070 ;
        RECT 2674.930 2680.290 2676.110 2681.470 ;
        RECT 2676.530 2680.290 2677.710 2681.470 ;
        RECT 2674.930 2501.890 2676.110 2503.070 ;
        RECT 2676.530 2501.890 2677.710 2503.070 ;
        RECT 2674.930 2500.290 2676.110 2501.470 ;
        RECT 2676.530 2500.290 2677.710 2501.470 ;
        RECT 2674.930 2321.890 2676.110 2323.070 ;
        RECT 2676.530 2321.890 2677.710 2323.070 ;
        RECT 2674.930 2320.290 2676.110 2321.470 ;
        RECT 2676.530 2320.290 2677.710 2321.470 ;
        RECT 2674.930 2141.890 2676.110 2143.070 ;
        RECT 2676.530 2141.890 2677.710 2143.070 ;
        RECT 2674.930 2140.290 2676.110 2141.470 ;
        RECT 2676.530 2140.290 2677.710 2141.470 ;
        RECT 2674.930 1961.890 2676.110 1963.070 ;
        RECT 2676.530 1961.890 2677.710 1963.070 ;
        RECT 2674.930 1960.290 2676.110 1961.470 ;
        RECT 2676.530 1960.290 2677.710 1961.470 ;
        RECT 2674.930 1781.890 2676.110 1783.070 ;
        RECT 2676.530 1781.890 2677.710 1783.070 ;
        RECT 2674.930 1780.290 2676.110 1781.470 ;
        RECT 2676.530 1780.290 2677.710 1781.470 ;
        RECT 2674.930 1601.890 2676.110 1603.070 ;
        RECT 2676.530 1601.890 2677.710 1603.070 ;
        RECT 2674.930 1600.290 2676.110 1601.470 ;
        RECT 2676.530 1600.290 2677.710 1601.470 ;
        RECT 2674.930 1421.890 2676.110 1423.070 ;
        RECT 2676.530 1421.890 2677.710 1423.070 ;
        RECT 2674.930 1420.290 2676.110 1421.470 ;
        RECT 2676.530 1420.290 2677.710 1421.470 ;
        RECT 2674.930 1241.890 2676.110 1243.070 ;
        RECT 2676.530 1241.890 2677.710 1243.070 ;
        RECT 2674.930 1240.290 2676.110 1241.470 ;
        RECT 2676.530 1240.290 2677.710 1241.470 ;
        RECT 2674.930 1061.890 2676.110 1063.070 ;
        RECT 2676.530 1061.890 2677.710 1063.070 ;
        RECT 2674.930 1060.290 2676.110 1061.470 ;
        RECT 2676.530 1060.290 2677.710 1061.470 ;
        RECT 2674.930 881.890 2676.110 883.070 ;
        RECT 2676.530 881.890 2677.710 883.070 ;
        RECT 2674.930 880.290 2676.110 881.470 ;
        RECT 2676.530 880.290 2677.710 881.470 ;
        RECT 2674.930 701.890 2676.110 703.070 ;
        RECT 2676.530 701.890 2677.710 703.070 ;
        RECT 2674.930 700.290 2676.110 701.470 ;
        RECT 2676.530 700.290 2677.710 701.470 ;
        RECT 2674.930 521.890 2676.110 523.070 ;
        RECT 2676.530 521.890 2677.710 523.070 ;
        RECT 2674.930 520.290 2676.110 521.470 ;
        RECT 2676.530 520.290 2677.710 521.470 ;
        RECT 2674.930 341.890 2676.110 343.070 ;
        RECT 2676.530 341.890 2677.710 343.070 ;
        RECT 2674.930 340.290 2676.110 341.470 ;
        RECT 2676.530 340.290 2677.710 341.470 ;
        RECT 2674.930 161.890 2676.110 163.070 ;
        RECT 2676.530 161.890 2677.710 163.070 ;
        RECT 2674.930 160.290 2676.110 161.470 ;
        RECT 2676.530 160.290 2677.710 161.470 ;
        RECT 2674.930 -36.510 2676.110 -35.330 ;
        RECT 2676.530 -36.510 2677.710 -35.330 ;
        RECT 2674.930 -38.110 2676.110 -36.930 ;
        RECT 2676.530 -38.110 2677.710 -36.930 ;
        RECT 2854.930 3556.610 2856.110 3557.790 ;
        RECT 2856.530 3556.610 2857.710 3557.790 ;
        RECT 2854.930 3555.010 2856.110 3556.190 ;
        RECT 2856.530 3555.010 2857.710 3556.190 ;
        RECT 2854.930 3401.890 2856.110 3403.070 ;
        RECT 2856.530 3401.890 2857.710 3403.070 ;
        RECT 2854.930 3400.290 2856.110 3401.470 ;
        RECT 2856.530 3400.290 2857.710 3401.470 ;
        RECT 2854.930 3221.890 2856.110 3223.070 ;
        RECT 2856.530 3221.890 2857.710 3223.070 ;
        RECT 2854.930 3220.290 2856.110 3221.470 ;
        RECT 2856.530 3220.290 2857.710 3221.470 ;
        RECT 2854.930 3041.890 2856.110 3043.070 ;
        RECT 2856.530 3041.890 2857.710 3043.070 ;
        RECT 2854.930 3040.290 2856.110 3041.470 ;
        RECT 2856.530 3040.290 2857.710 3041.470 ;
        RECT 2854.930 2861.890 2856.110 2863.070 ;
        RECT 2856.530 2861.890 2857.710 2863.070 ;
        RECT 2854.930 2860.290 2856.110 2861.470 ;
        RECT 2856.530 2860.290 2857.710 2861.470 ;
        RECT 2854.930 2681.890 2856.110 2683.070 ;
        RECT 2856.530 2681.890 2857.710 2683.070 ;
        RECT 2854.930 2680.290 2856.110 2681.470 ;
        RECT 2856.530 2680.290 2857.710 2681.470 ;
        RECT 2854.930 2501.890 2856.110 2503.070 ;
        RECT 2856.530 2501.890 2857.710 2503.070 ;
        RECT 2854.930 2500.290 2856.110 2501.470 ;
        RECT 2856.530 2500.290 2857.710 2501.470 ;
        RECT 2854.930 2321.890 2856.110 2323.070 ;
        RECT 2856.530 2321.890 2857.710 2323.070 ;
        RECT 2854.930 2320.290 2856.110 2321.470 ;
        RECT 2856.530 2320.290 2857.710 2321.470 ;
        RECT 2854.930 2141.890 2856.110 2143.070 ;
        RECT 2856.530 2141.890 2857.710 2143.070 ;
        RECT 2854.930 2140.290 2856.110 2141.470 ;
        RECT 2856.530 2140.290 2857.710 2141.470 ;
        RECT 2854.930 1961.890 2856.110 1963.070 ;
        RECT 2856.530 1961.890 2857.710 1963.070 ;
        RECT 2854.930 1960.290 2856.110 1961.470 ;
        RECT 2856.530 1960.290 2857.710 1961.470 ;
        RECT 2854.930 1781.890 2856.110 1783.070 ;
        RECT 2856.530 1781.890 2857.710 1783.070 ;
        RECT 2854.930 1780.290 2856.110 1781.470 ;
        RECT 2856.530 1780.290 2857.710 1781.470 ;
        RECT 2854.930 1601.890 2856.110 1603.070 ;
        RECT 2856.530 1601.890 2857.710 1603.070 ;
        RECT 2854.930 1600.290 2856.110 1601.470 ;
        RECT 2856.530 1600.290 2857.710 1601.470 ;
        RECT 2854.930 1421.890 2856.110 1423.070 ;
        RECT 2856.530 1421.890 2857.710 1423.070 ;
        RECT 2854.930 1420.290 2856.110 1421.470 ;
        RECT 2856.530 1420.290 2857.710 1421.470 ;
        RECT 2854.930 1241.890 2856.110 1243.070 ;
        RECT 2856.530 1241.890 2857.710 1243.070 ;
        RECT 2854.930 1240.290 2856.110 1241.470 ;
        RECT 2856.530 1240.290 2857.710 1241.470 ;
        RECT 2854.930 1061.890 2856.110 1063.070 ;
        RECT 2856.530 1061.890 2857.710 1063.070 ;
        RECT 2854.930 1060.290 2856.110 1061.470 ;
        RECT 2856.530 1060.290 2857.710 1061.470 ;
        RECT 2854.930 881.890 2856.110 883.070 ;
        RECT 2856.530 881.890 2857.710 883.070 ;
        RECT 2854.930 880.290 2856.110 881.470 ;
        RECT 2856.530 880.290 2857.710 881.470 ;
        RECT 2854.930 701.890 2856.110 703.070 ;
        RECT 2856.530 701.890 2857.710 703.070 ;
        RECT 2854.930 700.290 2856.110 701.470 ;
        RECT 2856.530 700.290 2857.710 701.470 ;
        RECT 2854.930 521.890 2856.110 523.070 ;
        RECT 2856.530 521.890 2857.710 523.070 ;
        RECT 2854.930 520.290 2856.110 521.470 ;
        RECT 2856.530 520.290 2857.710 521.470 ;
        RECT 2854.930 341.890 2856.110 343.070 ;
        RECT 2856.530 341.890 2857.710 343.070 ;
        RECT 2854.930 340.290 2856.110 341.470 ;
        RECT 2856.530 340.290 2857.710 341.470 ;
        RECT 2854.930 161.890 2856.110 163.070 ;
        RECT 2856.530 161.890 2857.710 163.070 ;
        RECT 2854.930 160.290 2856.110 161.470 ;
        RECT 2856.530 160.290 2857.710 161.470 ;
        RECT 2854.930 -36.510 2856.110 -35.330 ;
        RECT 2856.530 -36.510 2857.710 -35.330 ;
        RECT 2854.930 -38.110 2856.110 -36.930 ;
        RECT 2856.530 -38.110 2857.710 -36.930 ;
        RECT 2960.310 3556.610 2961.490 3557.790 ;
        RECT 2961.910 3556.610 2963.090 3557.790 ;
        RECT 2960.310 3555.010 2961.490 3556.190 ;
        RECT 2961.910 3555.010 2963.090 3556.190 ;
        RECT 2960.310 3401.890 2961.490 3403.070 ;
        RECT 2961.910 3401.890 2963.090 3403.070 ;
        RECT 2960.310 3400.290 2961.490 3401.470 ;
        RECT 2961.910 3400.290 2963.090 3401.470 ;
        RECT 2960.310 3221.890 2961.490 3223.070 ;
        RECT 2961.910 3221.890 2963.090 3223.070 ;
        RECT 2960.310 3220.290 2961.490 3221.470 ;
        RECT 2961.910 3220.290 2963.090 3221.470 ;
        RECT 2960.310 3041.890 2961.490 3043.070 ;
        RECT 2961.910 3041.890 2963.090 3043.070 ;
        RECT 2960.310 3040.290 2961.490 3041.470 ;
        RECT 2961.910 3040.290 2963.090 3041.470 ;
        RECT 2960.310 2861.890 2961.490 2863.070 ;
        RECT 2961.910 2861.890 2963.090 2863.070 ;
        RECT 2960.310 2860.290 2961.490 2861.470 ;
        RECT 2961.910 2860.290 2963.090 2861.470 ;
        RECT 2960.310 2681.890 2961.490 2683.070 ;
        RECT 2961.910 2681.890 2963.090 2683.070 ;
        RECT 2960.310 2680.290 2961.490 2681.470 ;
        RECT 2961.910 2680.290 2963.090 2681.470 ;
        RECT 2960.310 2501.890 2961.490 2503.070 ;
        RECT 2961.910 2501.890 2963.090 2503.070 ;
        RECT 2960.310 2500.290 2961.490 2501.470 ;
        RECT 2961.910 2500.290 2963.090 2501.470 ;
        RECT 2960.310 2321.890 2961.490 2323.070 ;
        RECT 2961.910 2321.890 2963.090 2323.070 ;
        RECT 2960.310 2320.290 2961.490 2321.470 ;
        RECT 2961.910 2320.290 2963.090 2321.470 ;
        RECT 2960.310 2141.890 2961.490 2143.070 ;
        RECT 2961.910 2141.890 2963.090 2143.070 ;
        RECT 2960.310 2140.290 2961.490 2141.470 ;
        RECT 2961.910 2140.290 2963.090 2141.470 ;
        RECT 2960.310 1961.890 2961.490 1963.070 ;
        RECT 2961.910 1961.890 2963.090 1963.070 ;
        RECT 2960.310 1960.290 2961.490 1961.470 ;
        RECT 2961.910 1960.290 2963.090 1961.470 ;
        RECT 2960.310 1781.890 2961.490 1783.070 ;
        RECT 2961.910 1781.890 2963.090 1783.070 ;
        RECT 2960.310 1780.290 2961.490 1781.470 ;
        RECT 2961.910 1780.290 2963.090 1781.470 ;
        RECT 2960.310 1601.890 2961.490 1603.070 ;
        RECT 2961.910 1601.890 2963.090 1603.070 ;
        RECT 2960.310 1600.290 2961.490 1601.470 ;
        RECT 2961.910 1600.290 2963.090 1601.470 ;
        RECT 2960.310 1421.890 2961.490 1423.070 ;
        RECT 2961.910 1421.890 2963.090 1423.070 ;
        RECT 2960.310 1420.290 2961.490 1421.470 ;
        RECT 2961.910 1420.290 2963.090 1421.470 ;
        RECT 2960.310 1241.890 2961.490 1243.070 ;
        RECT 2961.910 1241.890 2963.090 1243.070 ;
        RECT 2960.310 1240.290 2961.490 1241.470 ;
        RECT 2961.910 1240.290 2963.090 1241.470 ;
        RECT 2960.310 1061.890 2961.490 1063.070 ;
        RECT 2961.910 1061.890 2963.090 1063.070 ;
        RECT 2960.310 1060.290 2961.490 1061.470 ;
        RECT 2961.910 1060.290 2963.090 1061.470 ;
        RECT 2960.310 881.890 2961.490 883.070 ;
        RECT 2961.910 881.890 2963.090 883.070 ;
        RECT 2960.310 880.290 2961.490 881.470 ;
        RECT 2961.910 880.290 2963.090 881.470 ;
        RECT 2960.310 701.890 2961.490 703.070 ;
        RECT 2961.910 701.890 2963.090 703.070 ;
        RECT 2960.310 700.290 2961.490 701.470 ;
        RECT 2961.910 700.290 2963.090 701.470 ;
        RECT 2960.310 521.890 2961.490 523.070 ;
        RECT 2961.910 521.890 2963.090 523.070 ;
        RECT 2960.310 520.290 2961.490 521.470 ;
        RECT 2961.910 520.290 2963.090 521.470 ;
        RECT 2960.310 341.890 2961.490 343.070 ;
        RECT 2961.910 341.890 2963.090 343.070 ;
        RECT 2960.310 340.290 2961.490 341.470 ;
        RECT 2961.910 340.290 2963.090 341.470 ;
        RECT 2960.310 161.890 2961.490 163.070 ;
        RECT 2961.910 161.890 2963.090 163.070 ;
        RECT 2960.310 160.290 2961.490 161.470 ;
        RECT 2961.910 160.290 2963.090 161.470 ;
        RECT 2960.310 -36.510 2961.490 -35.330 ;
        RECT 2961.910 -36.510 2963.090 -35.330 ;
        RECT 2960.310 -38.110 2961.490 -36.930 ;
        RECT 2961.910 -38.110 2963.090 -36.930 ;
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
        RECT -43.630 880.130 2963.250 883.230 ;
        RECT -43.630 700.130 2963.250 703.230 ;
        RECT -43.630 520.130 2963.250 523.230 ;
        RECT -43.630 340.130 2963.250 343.230 ;
        RECT -43.630 160.130 2963.250 163.230 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
        RECT 278.970 1010.000 282.070 3529.150 ;
        RECT 458.970 1010.000 462.070 3529.150 ;
        RECT 638.970 1010.000 642.070 3529.150 ;
        RECT 818.970 1010.000 822.070 3529.150 ;
        RECT 998.970 1010.000 1002.070 3529.150 ;
        RECT 297.840 410.640 299.440 987.760 ;
        RECT 451.440 410.640 453.040 987.760 ;
        RECT 605.040 410.640 606.640 987.760 ;
        RECT 758.640 410.640 760.240 987.760 ;
        RECT 912.240 410.640 913.840 987.760 ;
        RECT 1065.840 410.640 1067.440 987.760 ;
        RECT 278.970 -9.470 282.070 390.000 ;
        RECT 458.970 -9.470 462.070 390.000 ;
        RECT 638.970 -9.470 642.070 390.000 ;
        RECT 818.970 -9.470 822.070 390.000 ;
        RECT 998.970 -9.470 1002.070 390.000 ;
        RECT 1178.970 -9.470 1182.070 3529.150 ;
        RECT 1358.970 -9.470 1362.070 3529.150 ;
        RECT 1538.970 -9.470 1542.070 3529.150 ;
        RECT 1718.970 -9.470 1722.070 3529.150 ;
        RECT 1898.970 -9.470 1902.070 3529.150 ;
        RECT 2078.970 -9.470 2082.070 3529.150 ;
        RECT 2258.970 -9.470 2262.070 3529.150 ;
        RECT 2438.970 -9.470 2442.070 3529.150 ;
        RECT 2618.970 -9.470 2622.070 3529.150 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
      LAYER via4 ;
        RECT -14.670 3527.810 -13.490 3528.990 ;
        RECT -13.070 3527.810 -11.890 3528.990 ;
        RECT -14.670 3526.210 -13.490 3527.390 ;
        RECT -13.070 3526.210 -11.890 3527.390 ;
        RECT -14.670 3346.090 -13.490 3347.270 ;
        RECT -13.070 3346.090 -11.890 3347.270 ;
        RECT -14.670 3344.490 -13.490 3345.670 ;
        RECT -13.070 3344.490 -11.890 3345.670 ;
        RECT -14.670 3166.090 -13.490 3167.270 ;
        RECT -13.070 3166.090 -11.890 3167.270 ;
        RECT -14.670 3164.490 -13.490 3165.670 ;
        RECT -13.070 3164.490 -11.890 3165.670 ;
        RECT -14.670 2986.090 -13.490 2987.270 ;
        RECT -13.070 2986.090 -11.890 2987.270 ;
        RECT -14.670 2984.490 -13.490 2985.670 ;
        RECT -13.070 2984.490 -11.890 2985.670 ;
        RECT -14.670 2806.090 -13.490 2807.270 ;
        RECT -13.070 2806.090 -11.890 2807.270 ;
        RECT -14.670 2804.490 -13.490 2805.670 ;
        RECT -13.070 2804.490 -11.890 2805.670 ;
        RECT -14.670 2626.090 -13.490 2627.270 ;
        RECT -13.070 2626.090 -11.890 2627.270 ;
        RECT -14.670 2624.490 -13.490 2625.670 ;
        RECT -13.070 2624.490 -11.890 2625.670 ;
        RECT -14.670 2446.090 -13.490 2447.270 ;
        RECT -13.070 2446.090 -11.890 2447.270 ;
        RECT -14.670 2444.490 -13.490 2445.670 ;
        RECT -13.070 2444.490 -11.890 2445.670 ;
        RECT -14.670 2266.090 -13.490 2267.270 ;
        RECT -13.070 2266.090 -11.890 2267.270 ;
        RECT -14.670 2264.490 -13.490 2265.670 ;
        RECT -13.070 2264.490 -11.890 2265.670 ;
        RECT -14.670 2086.090 -13.490 2087.270 ;
        RECT -13.070 2086.090 -11.890 2087.270 ;
        RECT -14.670 2084.490 -13.490 2085.670 ;
        RECT -13.070 2084.490 -11.890 2085.670 ;
        RECT -14.670 1906.090 -13.490 1907.270 ;
        RECT -13.070 1906.090 -11.890 1907.270 ;
        RECT -14.670 1904.490 -13.490 1905.670 ;
        RECT -13.070 1904.490 -11.890 1905.670 ;
        RECT -14.670 1726.090 -13.490 1727.270 ;
        RECT -13.070 1726.090 -11.890 1727.270 ;
        RECT -14.670 1724.490 -13.490 1725.670 ;
        RECT -13.070 1724.490 -11.890 1725.670 ;
        RECT -14.670 1546.090 -13.490 1547.270 ;
        RECT -13.070 1546.090 -11.890 1547.270 ;
        RECT -14.670 1544.490 -13.490 1545.670 ;
        RECT -13.070 1544.490 -11.890 1545.670 ;
        RECT -14.670 1366.090 -13.490 1367.270 ;
        RECT -13.070 1366.090 -11.890 1367.270 ;
        RECT -14.670 1364.490 -13.490 1365.670 ;
        RECT -13.070 1364.490 -11.890 1365.670 ;
        RECT -14.670 1186.090 -13.490 1187.270 ;
        RECT -13.070 1186.090 -11.890 1187.270 ;
        RECT -14.670 1184.490 -13.490 1185.670 ;
        RECT -13.070 1184.490 -11.890 1185.670 ;
        RECT -14.670 1006.090 -13.490 1007.270 ;
        RECT -13.070 1006.090 -11.890 1007.270 ;
        RECT -14.670 1004.490 -13.490 1005.670 ;
        RECT -13.070 1004.490 -11.890 1005.670 ;
        RECT -14.670 826.090 -13.490 827.270 ;
        RECT -13.070 826.090 -11.890 827.270 ;
        RECT -14.670 824.490 -13.490 825.670 ;
        RECT -13.070 824.490 -11.890 825.670 ;
        RECT -14.670 646.090 -13.490 647.270 ;
        RECT -13.070 646.090 -11.890 647.270 ;
        RECT -14.670 644.490 -13.490 645.670 ;
        RECT -13.070 644.490 -11.890 645.670 ;
        RECT -14.670 466.090 -13.490 467.270 ;
        RECT -13.070 466.090 -11.890 467.270 ;
        RECT -14.670 464.490 -13.490 465.670 ;
        RECT -13.070 464.490 -11.890 465.670 ;
        RECT -14.670 286.090 -13.490 287.270 ;
        RECT -13.070 286.090 -11.890 287.270 ;
        RECT -14.670 284.490 -13.490 285.670 ;
        RECT -13.070 284.490 -11.890 285.670 ;
        RECT -14.670 106.090 -13.490 107.270 ;
        RECT -13.070 106.090 -11.890 107.270 ;
        RECT -14.670 104.490 -13.490 105.670 ;
        RECT -13.070 104.490 -11.890 105.670 ;
        RECT -14.670 -7.710 -13.490 -6.530 ;
        RECT -13.070 -7.710 -11.890 -6.530 ;
        RECT -14.670 -9.310 -13.490 -8.130 ;
        RECT -13.070 -9.310 -11.890 -8.130 ;
        RECT 99.130 3527.810 100.310 3528.990 ;
        RECT 100.730 3527.810 101.910 3528.990 ;
        RECT 99.130 3526.210 100.310 3527.390 ;
        RECT 100.730 3526.210 101.910 3527.390 ;
        RECT 99.130 3346.090 100.310 3347.270 ;
        RECT 100.730 3346.090 101.910 3347.270 ;
        RECT 99.130 3344.490 100.310 3345.670 ;
        RECT 100.730 3344.490 101.910 3345.670 ;
        RECT 99.130 3166.090 100.310 3167.270 ;
        RECT 100.730 3166.090 101.910 3167.270 ;
        RECT 99.130 3164.490 100.310 3165.670 ;
        RECT 100.730 3164.490 101.910 3165.670 ;
        RECT 99.130 2986.090 100.310 2987.270 ;
        RECT 100.730 2986.090 101.910 2987.270 ;
        RECT 99.130 2984.490 100.310 2985.670 ;
        RECT 100.730 2984.490 101.910 2985.670 ;
        RECT 99.130 2806.090 100.310 2807.270 ;
        RECT 100.730 2806.090 101.910 2807.270 ;
        RECT 99.130 2804.490 100.310 2805.670 ;
        RECT 100.730 2804.490 101.910 2805.670 ;
        RECT 99.130 2626.090 100.310 2627.270 ;
        RECT 100.730 2626.090 101.910 2627.270 ;
        RECT 99.130 2624.490 100.310 2625.670 ;
        RECT 100.730 2624.490 101.910 2625.670 ;
        RECT 99.130 2446.090 100.310 2447.270 ;
        RECT 100.730 2446.090 101.910 2447.270 ;
        RECT 99.130 2444.490 100.310 2445.670 ;
        RECT 100.730 2444.490 101.910 2445.670 ;
        RECT 99.130 2266.090 100.310 2267.270 ;
        RECT 100.730 2266.090 101.910 2267.270 ;
        RECT 99.130 2264.490 100.310 2265.670 ;
        RECT 100.730 2264.490 101.910 2265.670 ;
        RECT 99.130 2086.090 100.310 2087.270 ;
        RECT 100.730 2086.090 101.910 2087.270 ;
        RECT 99.130 2084.490 100.310 2085.670 ;
        RECT 100.730 2084.490 101.910 2085.670 ;
        RECT 99.130 1906.090 100.310 1907.270 ;
        RECT 100.730 1906.090 101.910 1907.270 ;
        RECT 99.130 1904.490 100.310 1905.670 ;
        RECT 100.730 1904.490 101.910 1905.670 ;
        RECT 99.130 1726.090 100.310 1727.270 ;
        RECT 100.730 1726.090 101.910 1727.270 ;
        RECT 99.130 1724.490 100.310 1725.670 ;
        RECT 100.730 1724.490 101.910 1725.670 ;
        RECT 99.130 1546.090 100.310 1547.270 ;
        RECT 100.730 1546.090 101.910 1547.270 ;
        RECT 99.130 1544.490 100.310 1545.670 ;
        RECT 100.730 1544.490 101.910 1545.670 ;
        RECT 99.130 1366.090 100.310 1367.270 ;
        RECT 100.730 1366.090 101.910 1367.270 ;
        RECT 99.130 1364.490 100.310 1365.670 ;
        RECT 100.730 1364.490 101.910 1365.670 ;
        RECT 99.130 1186.090 100.310 1187.270 ;
        RECT 100.730 1186.090 101.910 1187.270 ;
        RECT 99.130 1184.490 100.310 1185.670 ;
        RECT 100.730 1184.490 101.910 1185.670 ;
        RECT 279.130 3527.810 280.310 3528.990 ;
        RECT 280.730 3527.810 281.910 3528.990 ;
        RECT 279.130 3526.210 280.310 3527.390 ;
        RECT 280.730 3526.210 281.910 3527.390 ;
        RECT 279.130 3346.090 280.310 3347.270 ;
        RECT 280.730 3346.090 281.910 3347.270 ;
        RECT 279.130 3344.490 280.310 3345.670 ;
        RECT 280.730 3344.490 281.910 3345.670 ;
        RECT 279.130 3166.090 280.310 3167.270 ;
        RECT 280.730 3166.090 281.910 3167.270 ;
        RECT 279.130 3164.490 280.310 3165.670 ;
        RECT 280.730 3164.490 281.910 3165.670 ;
        RECT 279.130 2986.090 280.310 2987.270 ;
        RECT 280.730 2986.090 281.910 2987.270 ;
        RECT 279.130 2984.490 280.310 2985.670 ;
        RECT 280.730 2984.490 281.910 2985.670 ;
        RECT 279.130 2806.090 280.310 2807.270 ;
        RECT 280.730 2806.090 281.910 2807.270 ;
        RECT 279.130 2804.490 280.310 2805.670 ;
        RECT 280.730 2804.490 281.910 2805.670 ;
        RECT 279.130 2626.090 280.310 2627.270 ;
        RECT 280.730 2626.090 281.910 2627.270 ;
        RECT 279.130 2624.490 280.310 2625.670 ;
        RECT 280.730 2624.490 281.910 2625.670 ;
        RECT 279.130 2446.090 280.310 2447.270 ;
        RECT 280.730 2446.090 281.910 2447.270 ;
        RECT 279.130 2444.490 280.310 2445.670 ;
        RECT 280.730 2444.490 281.910 2445.670 ;
        RECT 279.130 2266.090 280.310 2267.270 ;
        RECT 280.730 2266.090 281.910 2267.270 ;
        RECT 279.130 2264.490 280.310 2265.670 ;
        RECT 280.730 2264.490 281.910 2265.670 ;
        RECT 279.130 2086.090 280.310 2087.270 ;
        RECT 280.730 2086.090 281.910 2087.270 ;
        RECT 279.130 2084.490 280.310 2085.670 ;
        RECT 280.730 2084.490 281.910 2085.670 ;
        RECT 279.130 1906.090 280.310 1907.270 ;
        RECT 280.730 1906.090 281.910 1907.270 ;
        RECT 279.130 1904.490 280.310 1905.670 ;
        RECT 280.730 1904.490 281.910 1905.670 ;
        RECT 279.130 1726.090 280.310 1727.270 ;
        RECT 280.730 1726.090 281.910 1727.270 ;
        RECT 279.130 1724.490 280.310 1725.670 ;
        RECT 280.730 1724.490 281.910 1725.670 ;
        RECT 279.130 1546.090 280.310 1547.270 ;
        RECT 280.730 1546.090 281.910 1547.270 ;
        RECT 279.130 1544.490 280.310 1545.670 ;
        RECT 280.730 1544.490 281.910 1545.670 ;
        RECT 279.130 1366.090 280.310 1367.270 ;
        RECT 280.730 1366.090 281.910 1367.270 ;
        RECT 279.130 1364.490 280.310 1365.670 ;
        RECT 280.730 1364.490 281.910 1365.670 ;
        RECT 279.130 1186.090 280.310 1187.270 ;
        RECT 280.730 1186.090 281.910 1187.270 ;
        RECT 279.130 1184.490 280.310 1185.670 ;
        RECT 280.730 1184.490 281.910 1185.670 ;
        RECT 459.130 3527.810 460.310 3528.990 ;
        RECT 460.730 3527.810 461.910 3528.990 ;
        RECT 459.130 3526.210 460.310 3527.390 ;
        RECT 460.730 3526.210 461.910 3527.390 ;
        RECT 459.130 3346.090 460.310 3347.270 ;
        RECT 460.730 3346.090 461.910 3347.270 ;
        RECT 459.130 3344.490 460.310 3345.670 ;
        RECT 460.730 3344.490 461.910 3345.670 ;
        RECT 459.130 3166.090 460.310 3167.270 ;
        RECT 460.730 3166.090 461.910 3167.270 ;
        RECT 459.130 3164.490 460.310 3165.670 ;
        RECT 460.730 3164.490 461.910 3165.670 ;
        RECT 459.130 2986.090 460.310 2987.270 ;
        RECT 460.730 2986.090 461.910 2987.270 ;
        RECT 459.130 2984.490 460.310 2985.670 ;
        RECT 460.730 2984.490 461.910 2985.670 ;
        RECT 459.130 2806.090 460.310 2807.270 ;
        RECT 460.730 2806.090 461.910 2807.270 ;
        RECT 459.130 2804.490 460.310 2805.670 ;
        RECT 460.730 2804.490 461.910 2805.670 ;
        RECT 459.130 2626.090 460.310 2627.270 ;
        RECT 460.730 2626.090 461.910 2627.270 ;
        RECT 459.130 2624.490 460.310 2625.670 ;
        RECT 460.730 2624.490 461.910 2625.670 ;
        RECT 459.130 2446.090 460.310 2447.270 ;
        RECT 460.730 2446.090 461.910 2447.270 ;
        RECT 459.130 2444.490 460.310 2445.670 ;
        RECT 460.730 2444.490 461.910 2445.670 ;
        RECT 459.130 2266.090 460.310 2267.270 ;
        RECT 460.730 2266.090 461.910 2267.270 ;
        RECT 459.130 2264.490 460.310 2265.670 ;
        RECT 460.730 2264.490 461.910 2265.670 ;
        RECT 459.130 2086.090 460.310 2087.270 ;
        RECT 460.730 2086.090 461.910 2087.270 ;
        RECT 459.130 2084.490 460.310 2085.670 ;
        RECT 460.730 2084.490 461.910 2085.670 ;
        RECT 459.130 1906.090 460.310 1907.270 ;
        RECT 460.730 1906.090 461.910 1907.270 ;
        RECT 459.130 1904.490 460.310 1905.670 ;
        RECT 460.730 1904.490 461.910 1905.670 ;
        RECT 459.130 1726.090 460.310 1727.270 ;
        RECT 460.730 1726.090 461.910 1727.270 ;
        RECT 459.130 1724.490 460.310 1725.670 ;
        RECT 460.730 1724.490 461.910 1725.670 ;
        RECT 459.130 1546.090 460.310 1547.270 ;
        RECT 460.730 1546.090 461.910 1547.270 ;
        RECT 459.130 1544.490 460.310 1545.670 ;
        RECT 460.730 1544.490 461.910 1545.670 ;
        RECT 459.130 1366.090 460.310 1367.270 ;
        RECT 460.730 1366.090 461.910 1367.270 ;
        RECT 459.130 1364.490 460.310 1365.670 ;
        RECT 460.730 1364.490 461.910 1365.670 ;
        RECT 459.130 1186.090 460.310 1187.270 ;
        RECT 460.730 1186.090 461.910 1187.270 ;
        RECT 459.130 1184.490 460.310 1185.670 ;
        RECT 460.730 1184.490 461.910 1185.670 ;
        RECT 639.130 3527.810 640.310 3528.990 ;
        RECT 640.730 3527.810 641.910 3528.990 ;
        RECT 639.130 3526.210 640.310 3527.390 ;
        RECT 640.730 3526.210 641.910 3527.390 ;
        RECT 639.130 3346.090 640.310 3347.270 ;
        RECT 640.730 3346.090 641.910 3347.270 ;
        RECT 639.130 3344.490 640.310 3345.670 ;
        RECT 640.730 3344.490 641.910 3345.670 ;
        RECT 639.130 3166.090 640.310 3167.270 ;
        RECT 640.730 3166.090 641.910 3167.270 ;
        RECT 639.130 3164.490 640.310 3165.670 ;
        RECT 640.730 3164.490 641.910 3165.670 ;
        RECT 639.130 2986.090 640.310 2987.270 ;
        RECT 640.730 2986.090 641.910 2987.270 ;
        RECT 639.130 2984.490 640.310 2985.670 ;
        RECT 640.730 2984.490 641.910 2985.670 ;
        RECT 639.130 2806.090 640.310 2807.270 ;
        RECT 640.730 2806.090 641.910 2807.270 ;
        RECT 639.130 2804.490 640.310 2805.670 ;
        RECT 640.730 2804.490 641.910 2805.670 ;
        RECT 639.130 2626.090 640.310 2627.270 ;
        RECT 640.730 2626.090 641.910 2627.270 ;
        RECT 639.130 2624.490 640.310 2625.670 ;
        RECT 640.730 2624.490 641.910 2625.670 ;
        RECT 639.130 2446.090 640.310 2447.270 ;
        RECT 640.730 2446.090 641.910 2447.270 ;
        RECT 639.130 2444.490 640.310 2445.670 ;
        RECT 640.730 2444.490 641.910 2445.670 ;
        RECT 639.130 2266.090 640.310 2267.270 ;
        RECT 640.730 2266.090 641.910 2267.270 ;
        RECT 639.130 2264.490 640.310 2265.670 ;
        RECT 640.730 2264.490 641.910 2265.670 ;
        RECT 639.130 2086.090 640.310 2087.270 ;
        RECT 640.730 2086.090 641.910 2087.270 ;
        RECT 639.130 2084.490 640.310 2085.670 ;
        RECT 640.730 2084.490 641.910 2085.670 ;
        RECT 639.130 1906.090 640.310 1907.270 ;
        RECT 640.730 1906.090 641.910 1907.270 ;
        RECT 639.130 1904.490 640.310 1905.670 ;
        RECT 640.730 1904.490 641.910 1905.670 ;
        RECT 639.130 1726.090 640.310 1727.270 ;
        RECT 640.730 1726.090 641.910 1727.270 ;
        RECT 639.130 1724.490 640.310 1725.670 ;
        RECT 640.730 1724.490 641.910 1725.670 ;
        RECT 639.130 1546.090 640.310 1547.270 ;
        RECT 640.730 1546.090 641.910 1547.270 ;
        RECT 639.130 1544.490 640.310 1545.670 ;
        RECT 640.730 1544.490 641.910 1545.670 ;
        RECT 639.130 1366.090 640.310 1367.270 ;
        RECT 640.730 1366.090 641.910 1367.270 ;
        RECT 639.130 1364.490 640.310 1365.670 ;
        RECT 640.730 1364.490 641.910 1365.670 ;
        RECT 639.130 1186.090 640.310 1187.270 ;
        RECT 640.730 1186.090 641.910 1187.270 ;
        RECT 639.130 1184.490 640.310 1185.670 ;
        RECT 640.730 1184.490 641.910 1185.670 ;
        RECT 819.130 3527.810 820.310 3528.990 ;
        RECT 820.730 3527.810 821.910 3528.990 ;
        RECT 819.130 3526.210 820.310 3527.390 ;
        RECT 820.730 3526.210 821.910 3527.390 ;
        RECT 819.130 3346.090 820.310 3347.270 ;
        RECT 820.730 3346.090 821.910 3347.270 ;
        RECT 819.130 3344.490 820.310 3345.670 ;
        RECT 820.730 3344.490 821.910 3345.670 ;
        RECT 819.130 3166.090 820.310 3167.270 ;
        RECT 820.730 3166.090 821.910 3167.270 ;
        RECT 819.130 3164.490 820.310 3165.670 ;
        RECT 820.730 3164.490 821.910 3165.670 ;
        RECT 819.130 2986.090 820.310 2987.270 ;
        RECT 820.730 2986.090 821.910 2987.270 ;
        RECT 819.130 2984.490 820.310 2985.670 ;
        RECT 820.730 2984.490 821.910 2985.670 ;
        RECT 819.130 2806.090 820.310 2807.270 ;
        RECT 820.730 2806.090 821.910 2807.270 ;
        RECT 819.130 2804.490 820.310 2805.670 ;
        RECT 820.730 2804.490 821.910 2805.670 ;
        RECT 819.130 2626.090 820.310 2627.270 ;
        RECT 820.730 2626.090 821.910 2627.270 ;
        RECT 819.130 2624.490 820.310 2625.670 ;
        RECT 820.730 2624.490 821.910 2625.670 ;
        RECT 819.130 2446.090 820.310 2447.270 ;
        RECT 820.730 2446.090 821.910 2447.270 ;
        RECT 819.130 2444.490 820.310 2445.670 ;
        RECT 820.730 2444.490 821.910 2445.670 ;
        RECT 819.130 2266.090 820.310 2267.270 ;
        RECT 820.730 2266.090 821.910 2267.270 ;
        RECT 819.130 2264.490 820.310 2265.670 ;
        RECT 820.730 2264.490 821.910 2265.670 ;
        RECT 819.130 2086.090 820.310 2087.270 ;
        RECT 820.730 2086.090 821.910 2087.270 ;
        RECT 819.130 2084.490 820.310 2085.670 ;
        RECT 820.730 2084.490 821.910 2085.670 ;
        RECT 819.130 1906.090 820.310 1907.270 ;
        RECT 820.730 1906.090 821.910 1907.270 ;
        RECT 819.130 1904.490 820.310 1905.670 ;
        RECT 820.730 1904.490 821.910 1905.670 ;
        RECT 819.130 1726.090 820.310 1727.270 ;
        RECT 820.730 1726.090 821.910 1727.270 ;
        RECT 819.130 1724.490 820.310 1725.670 ;
        RECT 820.730 1724.490 821.910 1725.670 ;
        RECT 819.130 1546.090 820.310 1547.270 ;
        RECT 820.730 1546.090 821.910 1547.270 ;
        RECT 819.130 1544.490 820.310 1545.670 ;
        RECT 820.730 1544.490 821.910 1545.670 ;
        RECT 819.130 1366.090 820.310 1367.270 ;
        RECT 820.730 1366.090 821.910 1367.270 ;
        RECT 819.130 1364.490 820.310 1365.670 ;
        RECT 820.730 1364.490 821.910 1365.670 ;
        RECT 819.130 1186.090 820.310 1187.270 ;
        RECT 820.730 1186.090 821.910 1187.270 ;
        RECT 819.130 1184.490 820.310 1185.670 ;
        RECT 820.730 1184.490 821.910 1185.670 ;
        RECT 999.130 3527.810 1000.310 3528.990 ;
        RECT 1000.730 3527.810 1001.910 3528.990 ;
        RECT 999.130 3526.210 1000.310 3527.390 ;
        RECT 1000.730 3526.210 1001.910 3527.390 ;
        RECT 999.130 3346.090 1000.310 3347.270 ;
        RECT 1000.730 3346.090 1001.910 3347.270 ;
        RECT 999.130 3344.490 1000.310 3345.670 ;
        RECT 1000.730 3344.490 1001.910 3345.670 ;
        RECT 999.130 3166.090 1000.310 3167.270 ;
        RECT 1000.730 3166.090 1001.910 3167.270 ;
        RECT 999.130 3164.490 1000.310 3165.670 ;
        RECT 1000.730 3164.490 1001.910 3165.670 ;
        RECT 999.130 2986.090 1000.310 2987.270 ;
        RECT 1000.730 2986.090 1001.910 2987.270 ;
        RECT 999.130 2984.490 1000.310 2985.670 ;
        RECT 1000.730 2984.490 1001.910 2985.670 ;
        RECT 999.130 2806.090 1000.310 2807.270 ;
        RECT 1000.730 2806.090 1001.910 2807.270 ;
        RECT 999.130 2804.490 1000.310 2805.670 ;
        RECT 1000.730 2804.490 1001.910 2805.670 ;
        RECT 999.130 2626.090 1000.310 2627.270 ;
        RECT 1000.730 2626.090 1001.910 2627.270 ;
        RECT 999.130 2624.490 1000.310 2625.670 ;
        RECT 1000.730 2624.490 1001.910 2625.670 ;
        RECT 999.130 2446.090 1000.310 2447.270 ;
        RECT 1000.730 2446.090 1001.910 2447.270 ;
        RECT 999.130 2444.490 1000.310 2445.670 ;
        RECT 1000.730 2444.490 1001.910 2445.670 ;
        RECT 999.130 2266.090 1000.310 2267.270 ;
        RECT 1000.730 2266.090 1001.910 2267.270 ;
        RECT 999.130 2264.490 1000.310 2265.670 ;
        RECT 1000.730 2264.490 1001.910 2265.670 ;
        RECT 999.130 2086.090 1000.310 2087.270 ;
        RECT 1000.730 2086.090 1001.910 2087.270 ;
        RECT 999.130 2084.490 1000.310 2085.670 ;
        RECT 1000.730 2084.490 1001.910 2085.670 ;
        RECT 999.130 1906.090 1000.310 1907.270 ;
        RECT 1000.730 1906.090 1001.910 1907.270 ;
        RECT 999.130 1904.490 1000.310 1905.670 ;
        RECT 1000.730 1904.490 1001.910 1905.670 ;
        RECT 999.130 1726.090 1000.310 1727.270 ;
        RECT 1000.730 1726.090 1001.910 1727.270 ;
        RECT 999.130 1724.490 1000.310 1725.670 ;
        RECT 1000.730 1724.490 1001.910 1725.670 ;
        RECT 999.130 1546.090 1000.310 1547.270 ;
        RECT 1000.730 1546.090 1001.910 1547.270 ;
        RECT 999.130 1544.490 1000.310 1545.670 ;
        RECT 1000.730 1544.490 1001.910 1545.670 ;
        RECT 999.130 1366.090 1000.310 1367.270 ;
        RECT 1000.730 1366.090 1001.910 1367.270 ;
        RECT 999.130 1364.490 1000.310 1365.670 ;
        RECT 1000.730 1364.490 1001.910 1365.670 ;
        RECT 999.130 1186.090 1000.310 1187.270 ;
        RECT 1000.730 1186.090 1001.910 1187.270 ;
        RECT 999.130 1184.490 1000.310 1185.670 ;
        RECT 1000.730 1184.490 1001.910 1185.670 ;
        RECT 1179.130 3527.810 1180.310 3528.990 ;
        RECT 1180.730 3527.810 1181.910 3528.990 ;
        RECT 1179.130 3526.210 1180.310 3527.390 ;
        RECT 1180.730 3526.210 1181.910 3527.390 ;
        RECT 1179.130 3346.090 1180.310 3347.270 ;
        RECT 1180.730 3346.090 1181.910 3347.270 ;
        RECT 1179.130 3344.490 1180.310 3345.670 ;
        RECT 1180.730 3344.490 1181.910 3345.670 ;
        RECT 1179.130 3166.090 1180.310 3167.270 ;
        RECT 1180.730 3166.090 1181.910 3167.270 ;
        RECT 1179.130 3164.490 1180.310 3165.670 ;
        RECT 1180.730 3164.490 1181.910 3165.670 ;
        RECT 1179.130 2986.090 1180.310 2987.270 ;
        RECT 1180.730 2986.090 1181.910 2987.270 ;
        RECT 1179.130 2984.490 1180.310 2985.670 ;
        RECT 1180.730 2984.490 1181.910 2985.670 ;
        RECT 1179.130 2806.090 1180.310 2807.270 ;
        RECT 1180.730 2806.090 1181.910 2807.270 ;
        RECT 1179.130 2804.490 1180.310 2805.670 ;
        RECT 1180.730 2804.490 1181.910 2805.670 ;
        RECT 1179.130 2626.090 1180.310 2627.270 ;
        RECT 1180.730 2626.090 1181.910 2627.270 ;
        RECT 1179.130 2624.490 1180.310 2625.670 ;
        RECT 1180.730 2624.490 1181.910 2625.670 ;
        RECT 1179.130 2446.090 1180.310 2447.270 ;
        RECT 1180.730 2446.090 1181.910 2447.270 ;
        RECT 1179.130 2444.490 1180.310 2445.670 ;
        RECT 1180.730 2444.490 1181.910 2445.670 ;
        RECT 1179.130 2266.090 1180.310 2267.270 ;
        RECT 1180.730 2266.090 1181.910 2267.270 ;
        RECT 1179.130 2264.490 1180.310 2265.670 ;
        RECT 1180.730 2264.490 1181.910 2265.670 ;
        RECT 1179.130 2086.090 1180.310 2087.270 ;
        RECT 1180.730 2086.090 1181.910 2087.270 ;
        RECT 1179.130 2084.490 1180.310 2085.670 ;
        RECT 1180.730 2084.490 1181.910 2085.670 ;
        RECT 1179.130 1906.090 1180.310 1907.270 ;
        RECT 1180.730 1906.090 1181.910 1907.270 ;
        RECT 1179.130 1904.490 1180.310 1905.670 ;
        RECT 1180.730 1904.490 1181.910 1905.670 ;
        RECT 1179.130 1726.090 1180.310 1727.270 ;
        RECT 1180.730 1726.090 1181.910 1727.270 ;
        RECT 1179.130 1724.490 1180.310 1725.670 ;
        RECT 1180.730 1724.490 1181.910 1725.670 ;
        RECT 1179.130 1546.090 1180.310 1547.270 ;
        RECT 1180.730 1546.090 1181.910 1547.270 ;
        RECT 1179.130 1544.490 1180.310 1545.670 ;
        RECT 1180.730 1544.490 1181.910 1545.670 ;
        RECT 1179.130 1366.090 1180.310 1367.270 ;
        RECT 1180.730 1366.090 1181.910 1367.270 ;
        RECT 1179.130 1364.490 1180.310 1365.670 ;
        RECT 1180.730 1364.490 1181.910 1365.670 ;
        RECT 1179.130 1186.090 1180.310 1187.270 ;
        RECT 1180.730 1186.090 1181.910 1187.270 ;
        RECT 1179.130 1184.490 1180.310 1185.670 ;
        RECT 1180.730 1184.490 1181.910 1185.670 ;
        RECT 99.130 1006.090 100.310 1007.270 ;
        RECT 100.730 1006.090 101.910 1007.270 ;
        RECT 99.130 1004.490 100.310 1005.670 ;
        RECT 100.730 1004.490 101.910 1005.670 ;
        RECT 1179.130 1006.090 1180.310 1007.270 ;
        RECT 1180.730 1006.090 1181.910 1007.270 ;
        RECT 1179.130 1004.490 1180.310 1005.670 ;
        RECT 1180.730 1004.490 1181.910 1005.670 ;
        RECT 99.130 826.090 100.310 827.270 ;
        RECT 100.730 826.090 101.910 827.270 ;
        RECT 99.130 824.490 100.310 825.670 ;
        RECT 100.730 824.490 101.910 825.670 ;
        RECT 99.130 646.090 100.310 647.270 ;
        RECT 100.730 646.090 101.910 647.270 ;
        RECT 99.130 644.490 100.310 645.670 ;
        RECT 100.730 644.490 101.910 645.670 ;
        RECT 99.130 466.090 100.310 467.270 ;
        RECT 100.730 466.090 101.910 467.270 ;
        RECT 99.130 464.490 100.310 465.670 ;
        RECT 100.730 464.490 101.910 465.670 ;
        RECT 298.050 826.090 299.230 827.270 ;
        RECT 298.050 824.490 299.230 825.670 ;
        RECT 298.050 646.090 299.230 647.270 ;
        RECT 298.050 644.490 299.230 645.670 ;
        RECT 298.050 466.090 299.230 467.270 ;
        RECT 298.050 464.490 299.230 465.670 ;
        RECT 451.650 826.090 452.830 827.270 ;
        RECT 451.650 824.490 452.830 825.670 ;
        RECT 451.650 646.090 452.830 647.270 ;
        RECT 451.650 644.490 452.830 645.670 ;
        RECT 451.650 466.090 452.830 467.270 ;
        RECT 451.650 464.490 452.830 465.670 ;
        RECT 605.250 826.090 606.430 827.270 ;
        RECT 605.250 824.490 606.430 825.670 ;
        RECT 605.250 646.090 606.430 647.270 ;
        RECT 605.250 644.490 606.430 645.670 ;
        RECT 605.250 466.090 606.430 467.270 ;
        RECT 605.250 464.490 606.430 465.670 ;
        RECT 758.850 826.090 760.030 827.270 ;
        RECT 758.850 824.490 760.030 825.670 ;
        RECT 758.850 646.090 760.030 647.270 ;
        RECT 758.850 644.490 760.030 645.670 ;
        RECT 758.850 466.090 760.030 467.270 ;
        RECT 758.850 464.490 760.030 465.670 ;
        RECT 912.450 826.090 913.630 827.270 ;
        RECT 912.450 824.490 913.630 825.670 ;
        RECT 912.450 646.090 913.630 647.270 ;
        RECT 912.450 644.490 913.630 645.670 ;
        RECT 912.450 466.090 913.630 467.270 ;
        RECT 912.450 464.490 913.630 465.670 ;
        RECT 1066.050 826.090 1067.230 827.270 ;
        RECT 1066.050 824.490 1067.230 825.670 ;
        RECT 1066.050 646.090 1067.230 647.270 ;
        RECT 1066.050 644.490 1067.230 645.670 ;
        RECT 1066.050 466.090 1067.230 467.270 ;
        RECT 1066.050 464.490 1067.230 465.670 ;
        RECT 1179.130 826.090 1180.310 827.270 ;
        RECT 1180.730 826.090 1181.910 827.270 ;
        RECT 1179.130 824.490 1180.310 825.670 ;
        RECT 1180.730 824.490 1181.910 825.670 ;
        RECT 1179.130 646.090 1180.310 647.270 ;
        RECT 1180.730 646.090 1181.910 647.270 ;
        RECT 1179.130 644.490 1180.310 645.670 ;
        RECT 1180.730 644.490 1181.910 645.670 ;
        RECT 1179.130 466.090 1180.310 467.270 ;
        RECT 1180.730 466.090 1181.910 467.270 ;
        RECT 1179.130 464.490 1180.310 465.670 ;
        RECT 1180.730 464.490 1181.910 465.670 ;
        RECT 99.130 286.090 100.310 287.270 ;
        RECT 100.730 286.090 101.910 287.270 ;
        RECT 99.130 284.490 100.310 285.670 ;
        RECT 100.730 284.490 101.910 285.670 ;
        RECT 99.130 106.090 100.310 107.270 ;
        RECT 100.730 106.090 101.910 107.270 ;
        RECT 99.130 104.490 100.310 105.670 ;
        RECT 100.730 104.490 101.910 105.670 ;
        RECT 99.130 -7.710 100.310 -6.530 ;
        RECT 100.730 -7.710 101.910 -6.530 ;
        RECT 99.130 -9.310 100.310 -8.130 ;
        RECT 100.730 -9.310 101.910 -8.130 ;
        RECT 279.130 286.090 280.310 287.270 ;
        RECT 280.730 286.090 281.910 287.270 ;
        RECT 279.130 284.490 280.310 285.670 ;
        RECT 280.730 284.490 281.910 285.670 ;
        RECT 279.130 106.090 280.310 107.270 ;
        RECT 280.730 106.090 281.910 107.270 ;
        RECT 279.130 104.490 280.310 105.670 ;
        RECT 280.730 104.490 281.910 105.670 ;
        RECT 279.130 -7.710 280.310 -6.530 ;
        RECT 280.730 -7.710 281.910 -6.530 ;
        RECT 279.130 -9.310 280.310 -8.130 ;
        RECT 280.730 -9.310 281.910 -8.130 ;
        RECT 459.130 286.090 460.310 287.270 ;
        RECT 460.730 286.090 461.910 287.270 ;
        RECT 459.130 284.490 460.310 285.670 ;
        RECT 460.730 284.490 461.910 285.670 ;
        RECT 459.130 106.090 460.310 107.270 ;
        RECT 460.730 106.090 461.910 107.270 ;
        RECT 459.130 104.490 460.310 105.670 ;
        RECT 460.730 104.490 461.910 105.670 ;
        RECT 459.130 -7.710 460.310 -6.530 ;
        RECT 460.730 -7.710 461.910 -6.530 ;
        RECT 459.130 -9.310 460.310 -8.130 ;
        RECT 460.730 -9.310 461.910 -8.130 ;
        RECT 639.130 286.090 640.310 287.270 ;
        RECT 640.730 286.090 641.910 287.270 ;
        RECT 639.130 284.490 640.310 285.670 ;
        RECT 640.730 284.490 641.910 285.670 ;
        RECT 639.130 106.090 640.310 107.270 ;
        RECT 640.730 106.090 641.910 107.270 ;
        RECT 639.130 104.490 640.310 105.670 ;
        RECT 640.730 104.490 641.910 105.670 ;
        RECT 639.130 -7.710 640.310 -6.530 ;
        RECT 640.730 -7.710 641.910 -6.530 ;
        RECT 639.130 -9.310 640.310 -8.130 ;
        RECT 640.730 -9.310 641.910 -8.130 ;
        RECT 819.130 286.090 820.310 287.270 ;
        RECT 820.730 286.090 821.910 287.270 ;
        RECT 819.130 284.490 820.310 285.670 ;
        RECT 820.730 284.490 821.910 285.670 ;
        RECT 819.130 106.090 820.310 107.270 ;
        RECT 820.730 106.090 821.910 107.270 ;
        RECT 819.130 104.490 820.310 105.670 ;
        RECT 820.730 104.490 821.910 105.670 ;
        RECT 819.130 -7.710 820.310 -6.530 ;
        RECT 820.730 -7.710 821.910 -6.530 ;
        RECT 819.130 -9.310 820.310 -8.130 ;
        RECT 820.730 -9.310 821.910 -8.130 ;
        RECT 999.130 286.090 1000.310 287.270 ;
        RECT 1000.730 286.090 1001.910 287.270 ;
        RECT 999.130 284.490 1000.310 285.670 ;
        RECT 1000.730 284.490 1001.910 285.670 ;
        RECT 999.130 106.090 1000.310 107.270 ;
        RECT 1000.730 106.090 1001.910 107.270 ;
        RECT 999.130 104.490 1000.310 105.670 ;
        RECT 1000.730 104.490 1001.910 105.670 ;
        RECT 999.130 -7.710 1000.310 -6.530 ;
        RECT 1000.730 -7.710 1001.910 -6.530 ;
        RECT 999.130 -9.310 1000.310 -8.130 ;
        RECT 1000.730 -9.310 1001.910 -8.130 ;
        RECT 1179.130 286.090 1180.310 287.270 ;
        RECT 1180.730 286.090 1181.910 287.270 ;
        RECT 1179.130 284.490 1180.310 285.670 ;
        RECT 1180.730 284.490 1181.910 285.670 ;
        RECT 1179.130 106.090 1180.310 107.270 ;
        RECT 1180.730 106.090 1181.910 107.270 ;
        RECT 1179.130 104.490 1180.310 105.670 ;
        RECT 1180.730 104.490 1181.910 105.670 ;
        RECT 1179.130 -7.710 1180.310 -6.530 ;
        RECT 1180.730 -7.710 1181.910 -6.530 ;
        RECT 1179.130 -9.310 1180.310 -8.130 ;
        RECT 1180.730 -9.310 1181.910 -8.130 ;
        RECT 1359.130 3527.810 1360.310 3528.990 ;
        RECT 1360.730 3527.810 1361.910 3528.990 ;
        RECT 1359.130 3526.210 1360.310 3527.390 ;
        RECT 1360.730 3526.210 1361.910 3527.390 ;
        RECT 1359.130 3346.090 1360.310 3347.270 ;
        RECT 1360.730 3346.090 1361.910 3347.270 ;
        RECT 1359.130 3344.490 1360.310 3345.670 ;
        RECT 1360.730 3344.490 1361.910 3345.670 ;
        RECT 1359.130 3166.090 1360.310 3167.270 ;
        RECT 1360.730 3166.090 1361.910 3167.270 ;
        RECT 1359.130 3164.490 1360.310 3165.670 ;
        RECT 1360.730 3164.490 1361.910 3165.670 ;
        RECT 1359.130 2986.090 1360.310 2987.270 ;
        RECT 1360.730 2986.090 1361.910 2987.270 ;
        RECT 1359.130 2984.490 1360.310 2985.670 ;
        RECT 1360.730 2984.490 1361.910 2985.670 ;
        RECT 1359.130 2806.090 1360.310 2807.270 ;
        RECT 1360.730 2806.090 1361.910 2807.270 ;
        RECT 1359.130 2804.490 1360.310 2805.670 ;
        RECT 1360.730 2804.490 1361.910 2805.670 ;
        RECT 1359.130 2626.090 1360.310 2627.270 ;
        RECT 1360.730 2626.090 1361.910 2627.270 ;
        RECT 1359.130 2624.490 1360.310 2625.670 ;
        RECT 1360.730 2624.490 1361.910 2625.670 ;
        RECT 1359.130 2446.090 1360.310 2447.270 ;
        RECT 1360.730 2446.090 1361.910 2447.270 ;
        RECT 1359.130 2444.490 1360.310 2445.670 ;
        RECT 1360.730 2444.490 1361.910 2445.670 ;
        RECT 1359.130 2266.090 1360.310 2267.270 ;
        RECT 1360.730 2266.090 1361.910 2267.270 ;
        RECT 1359.130 2264.490 1360.310 2265.670 ;
        RECT 1360.730 2264.490 1361.910 2265.670 ;
        RECT 1359.130 2086.090 1360.310 2087.270 ;
        RECT 1360.730 2086.090 1361.910 2087.270 ;
        RECT 1359.130 2084.490 1360.310 2085.670 ;
        RECT 1360.730 2084.490 1361.910 2085.670 ;
        RECT 1359.130 1906.090 1360.310 1907.270 ;
        RECT 1360.730 1906.090 1361.910 1907.270 ;
        RECT 1359.130 1904.490 1360.310 1905.670 ;
        RECT 1360.730 1904.490 1361.910 1905.670 ;
        RECT 1359.130 1726.090 1360.310 1727.270 ;
        RECT 1360.730 1726.090 1361.910 1727.270 ;
        RECT 1359.130 1724.490 1360.310 1725.670 ;
        RECT 1360.730 1724.490 1361.910 1725.670 ;
        RECT 1359.130 1546.090 1360.310 1547.270 ;
        RECT 1360.730 1546.090 1361.910 1547.270 ;
        RECT 1359.130 1544.490 1360.310 1545.670 ;
        RECT 1360.730 1544.490 1361.910 1545.670 ;
        RECT 1359.130 1366.090 1360.310 1367.270 ;
        RECT 1360.730 1366.090 1361.910 1367.270 ;
        RECT 1359.130 1364.490 1360.310 1365.670 ;
        RECT 1360.730 1364.490 1361.910 1365.670 ;
        RECT 1359.130 1186.090 1360.310 1187.270 ;
        RECT 1360.730 1186.090 1361.910 1187.270 ;
        RECT 1359.130 1184.490 1360.310 1185.670 ;
        RECT 1360.730 1184.490 1361.910 1185.670 ;
        RECT 1359.130 1006.090 1360.310 1007.270 ;
        RECT 1360.730 1006.090 1361.910 1007.270 ;
        RECT 1359.130 1004.490 1360.310 1005.670 ;
        RECT 1360.730 1004.490 1361.910 1005.670 ;
        RECT 1359.130 826.090 1360.310 827.270 ;
        RECT 1360.730 826.090 1361.910 827.270 ;
        RECT 1359.130 824.490 1360.310 825.670 ;
        RECT 1360.730 824.490 1361.910 825.670 ;
        RECT 1359.130 646.090 1360.310 647.270 ;
        RECT 1360.730 646.090 1361.910 647.270 ;
        RECT 1359.130 644.490 1360.310 645.670 ;
        RECT 1360.730 644.490 1361.910 645.670 ;
        RECT 1359.130 466.090 1360.310 467.270 ;
        RECT 1360.730 466.090 1361.910 467.270 ;
        RECT 1359.130 464.490 1360.310 465.670 ;
        RECT 1360.730 464.490 1361.910 465.670 ;
        RECT 1359.130 286.090 1360.310 287.270 ;
        RECT 1360.730 286.090 1361.910 287.270 ;
        RECT 1359.130 284.490 1360.310 285.670 ;
        RECT 1360.730 284.490 1361.910 285.670 ;
        RECT 1359.130 106.090 1360.310 107.270 ;
        RECT 1360.730 106.090 1361.910 107.270 ;
        RECT 1359.130 104.490 1360.310 105.670 ;
        RECT 1360.730 104.490 1361.910 105.670 ;
        RECT 1359.130 -7.710 1360.310 -6.530 ;
        RECT 1360.730 -7.710 1361.910 -6.530 ;
        RECT 1359.130 -9.310 1360.310 -8.130 ;
        RECT 1360.730 -9.310 1361.910 -8.130 ;
        RECT 1539.130 3527.810 1540.310 3528.990 ;
        RECT 1540.730 3527.810 1541.910 3528.990 ;
        RECT 1539.130 3526.210 1540.310 3527.390 ;
        RECT 1540.730 3526.210 1541.910 3527.390 ;
        RECT 1539.130 3346.090 1540.310 3347.270 ;
        RECT 1540.730 3346.090 1541.910 3347.270 ;
        RECT 1539.130 3344.490 1540.310 3345.670 ;
        RECT 1540.730 3344.490 1541.910 3345.670 ;
        RECT 1539.130 3166.090 1540.310 3167.270 ;
        RECT 1540.730 3166.090 1541.910 3167.270 ;
        RECT 1539.130 3164.490 1540.310 3165.670 ;
        RECT 1540.730 3164.490 1541.910 3165.670 ;
        RECT 1539.130 2986.090 1540.310 2987.270 ;
        RECT 1540.730 2986.090 1541.910 2987.270 ;
        RECT 1539.130 2984.490 1540.310 2985.670 ;
        RECT 1540.730 2984.490 1541.910 2985.670 ;
        RECT 1539.130 2806.090 1540.310 2807.270 ;
        RECT 1540.730 2806.090 1541.910 2807.270 ;
        RECT 1539.130 2804.490 1540.310 2805.670 ;
        RECT 1540.730 2804.490 1541.910 2805.670 ;
        RECT 1539.130 2626.090 1540.310 2627.270 ;
        RECT 1540.730 2626.090 1541.910 2627.270 ;
        RECT 1539.130 2624.490 1540.310 2625.670 ;
        RECT 1540.730 2624.490 1541.910 2625.670 ;
        RECT 1539.130 2446.090 1540.310 2447.270 ;
        RECT 1540.730 2446.090 1541.910 2447.270 ;
        RECT 1539.130 2444.490 1540.310 2445.670 ;
        RECT 1540.730 2444.490 1541.910 2445.670 ;
        RECT 1539.130 2266.090 1540.310 2267.270 ;
        RECT 1540.730 2266.090 1541.910 2267.270 ;
        RECT 1539.130 2264.490 1540.310 2265.670 ;
        RECT 1540.730 2264.490 1541.910 2265.670 ;
        RECT 1539.130 2086.090 1540.310 2087.270 ;
        RECT 1540.730 2086.090 1541.910 2087.270 ;
        RECT 1539.130 2084.490 1540.310 2085.670 ;
        RECT 1540.730 2084.490 1541.910 2085.670 ;
        RECT 1539.130 1906.090 1540.310 1907.270 ;
        RECT 1540.730 1906.090 1541.910 1907.270 ;
        RECT 1539.130 1904.490 1540.310 1905.670 ;
        RECT 1540.730 1904.490 1541.910 1905.670 ;
        RECT 1539.130 1726.090 1540.310 1727.270 ;
        RECT 1540.730 1726.090 1541.910 1727.270 ;
        RECT 1539.130 1724.490 1540.310 1725.670 ;
        RECT 1540.730 1724.490 1541.910 1725.670 ;
        RECT 1539.130 1546.090 1540.310 1547.270 ;
        RECT 1540.730 1546.090 1541.910 1547.270 ;
        RECT 1539.130 1544.490 1540.310 1545.670 ;
        RECT 1540.730 1544.490 1541.910 1545.670 ;
        RECT 1539.130 1366.090 1540.310 1367.270 ;
        RECT 1540.730 1366.090 1541.910 1367.270 ;
        RECT 1539.130 1364.490 1540.310 1365.670 ;
        RECT 1540.730 1364.490 1541.910 1365.670 ;
        RECT 1539.130 1186.090 1540.310 1187.270 ;
        RECT 1540.730 1186.090 1541.910 1187.270 ;
        RECT 1539.130 1184.490 1540.310 1185.670 ;
        RECT 1540.730 1184.490 1541.910 1185.670 ;
        RECT 1539.130 1006.090 1540.310 1007.270 ;
        RECT 1540.730 1006.090 1541.910 1007.270 ;
        RECT 1539.130 1004.490 1540.310 1005.670 ;
        RECT 1540.730 1004.490 1541.910 1005.670 ;
        RECT 1539.130 826.090 1540.310 827.270 ;
        RECT 1540.730 826.090 1541.910 827.270 ;
        RECT 1539.130 824.490 1540.310 825.670 ;
        RECT 1540.730 824.490 1541.910 825.670 ;
        RECT 1539.130 646.090 1540.310 647.270 ;
        RECT 1540.730 646.090 1541.910 647.270 ;
        RECT 1539.130 644.490 1540.310 645.670 ;
        RECT 1540.730 644.490 1541.910 645.670 ;
        RECT 1539.130 466.090 1540.310 467.270 ;
        RECT 1540.730 466.090 1541.910 467.270 ;
        RECT 1539.130 464.490 1540.310 465.670 ;
        RECT 1540.730 464.490 1541.910 465.670 ;
        RECT 1539.130 286.090 1540.310 287.270 ;
        RECT 1540.730 286.090 1541.910 287.270 ;
        RECT 1539.130 284.490 1540.310 285.670 ;
        RECT 1540.730 284.490 1541.910 285.670 ;
        RECT 1539.130 106.090 1540.310 107.270 ;
        RECT 1540.730 106.090 1541.910 107.270 ;
        RECT 1539.130 104.490 1540.310 105.670 ;
        RECT 1540.730 104.490 1541.910 105.670 ;
        RECT 1539.130 -7.710 1540.310 -6.530 ;
        RECT 1540.730 -7.710 1541.910 -6.530 ;
        RECT 1539.130 -9.310 1540.310 -8.130 ;
        RECT 1540.730 -9.310 1541.910 -8.130 ;
        RECT 1719.130 3527.810 1720.310 3528.990 ;
        RECT 1720.730 3527.810 1721.910 3528.990 ;
        RECT 1719.130 3526.210 1720.310 3527.390 ;
        RECT 1720.730 3526.210 1721.910 3527.390 ;
        RECT 1719.130 3346.090 1720.310 3347.270 ;
        RECT 1720.730 3346.090 1721.910 3347.270 ;
        RECT 1719.130 3344.490 1720.310 3345.670 ;
        RECT 1720.730 3344.490 1721.910 3345.670 ;
        RECT 1719.130 3166.090 1720.310 3167.270 ;
        RECT 1720.730 3166.090 1721.910 3167.270 ;
        RECT 1719.130 3164.490 1720.310 3165.670 ;
        RECT 1720.730 3164.490 1721.910 3165.670 ;
        RECT 1719.130 2986.090 1720.310 2987.270 ;
        RECT 1720.730 2986.090 1721.910 2987.270 ;
        RECT 1719.130 2984.490 1720.310 2985.670 ;
        RECT 1720.730 2984.490 1721.910 2985.670 ;
        RECT 1719.130 2806.090 1720.310 2807.270 ;
        RECT 1720.730 2806.090 1721.910 2807.270 ;
        RECT 1719.130 2804.490 1720.310 2805.670 ;
        RECT 1720.730 2804.490 1721.910 2805.670 ;
        RECT 1719.130 2626.090 1720.310 2627.270 ;
        RECT 1720.730 2626.090 1721.910 2627.270 ;
        RECT 1719.130 2624.490 1720.310 2625.670 ;
        RECT 1720.730 2624.490 1721.910 2625.670 ;
        RECT 1719.130 2446.090 1720.310 2447.270 ;
        RECT 1720.730 2446.090 1721.910 2447.270 ;
        RECT 1719.130 2444.490 1720.310 2445.670 ;
        RECT 1720.730 2444.490 1721.910 2445.670 ;
        RECT 1719.130 2266.090 1720.310 2267.270 ;
        RECT 1720.730 2266.090 1721.910 2267.270 ;
        RECT 1719.130 2264.490 1720.310 2265.670 ;
        RECT 1720.730 2264.490 1721.910 2265.670 ;
        RECT 1719.130 2086.090 1720.310 2087.270 ;
        RECT 1720.730 2086.090 1721.910 2087.270 ;
        RECT 1719.130 2084.490 1720.310 2085.670 ;
        RECT 1720.730 2084.490 1721.910 2085.670 ;
        RECT 1719.130 1906.090 1720.310 1907.270 ;
        RECT 1720.730 1906.090 1721.910 1907.270 ;
        RECT 1719.130 1904.490 1720.310 1905.670 ;
        RECT 1720.730 1904.490 1721.910 1905.670 ;
        RECT 1719.130 1726.090 1720.310 1727.270 ;
        RECT 1720.730 1726.090 1721.910 1727.270 ;
        RECT 1719.130 1724.490 1720.310 1725.670 ;
        RECT 1720.730 1724.490 1721.910 1725.670 ;
        RECT 1719.130 1546.090 1720.310 1547.270 ;
        RECT 1720.730 1546.090 1721.910 1547.270 ;
        RECT 1719.130 1544.490 1720.310 1545.670 ;
        RECT 1720.730 1544.490 1721.910 1545.670 ;
        RECT 1719.130 1366.090 1720.310 1367.270 ;
        RECT 1720.730 1366.090 1721.910 1367.270 ;
        RECT 1719.130 1364.490 1720.310 1365.670 ;
        RECT 1720.730 1364.490 1721.910 1365.670 ;
        RECT 1719.130 1186.090 1720.310 1187.270 ;
        RECT 1720.730 1186.090 1721.910 1187.270 ;
        RECT 1719.130 1184.490 1720.310 1185.670 ;
        RECT 1720.730 1184.490 1721.910 1185.670 ;
        RECT 1719.130 1006.090 1720.310 1007.270 ;
        RECT 1720.730 1006.090 1721.910 1007.270 ;
        RECT 1719.130 1004.490 1720.310 1005.670 ;
        RECT 1720.730 1004.490 1721.910 1005.670 ;
        RECT 1719.130 826.090 1720.310 827.270 ;
        RECT 1720.730 826.090 1721.910 827.270 ;
        RECT 1719.130 824.490 1720.310 825.670 ;
        RECT 1720.730 824.490 1721.910 825.670 ;
        RECT 1719.130 646.090 1720.310 647.270 ;
        RECT 1720.730 646.090 1721.910 647.270 ;
        RECT 1719.130 644.490 1720.310 645.670 ;
        RECT 1720.730 644.490 1721.910 645.670 ;
        RECT 1719.130 466.090 1720.310 467.270 ;
        RECT 1720.730 466.090 1721.910 467.270 ;
        RECT 1719.130 464.490 1720.310 465.670 ;
        RECT 1720.730 464.490 1721.910 465.670 ;
        RECT 1719.130 286.090 1720.310 287.270 ;
        RECT 1720.730 286.090 1721.910 287.270 ;
        RECT 1719.130 284.490 1720.310 285.670 ;
        RECT 1720.730 284.490 1721.910 285.670 ;
        RECT 1719.130 106.090 1720.310 107.270 ;
        RECT 1720.730 106.090 1721.910 107.270 ;
        RECT 1719.130 104.490 1720.310 105.670 ;
        RECT 1720.730 104.490 1721.910 105.670 ;
        RECT 1719.130 -7.710 1720.310 -6.530 ;
        RECT 1720.730 -7.710 1721.910 -6.530 ;
        RECT 1719.130 -9.310 1720.310 -8.130 ;
        RECT 1720.730 -9.310 1721.910 -8.130 ;
        RECT 1899.130 3527.810 1900.310 3528.990 ;
        RECT 1900.730 3527.810 1901.910 3528.990 ;
        RECT 1899.130 3526.210 1900.310 3527.390 ;
        RECT 1900.730 3526.210 1901.910 3527.390 ;
        RECT 1899.130 3346.090 1900.310 3347.270 ;
        RECT 1900.730 3346.090 1901.910 3347.270 ;
        RECT 1899.130 3344.490 1900.310 3345.670 ;
        RECT 1900.730 3344.490 1901.910 3345.670 ;
        RECT 1899.130 3166.090 1900.310 3167.270 ;
        RECT 1900.730 3166.090 1901.910 3167.270 ;
        RECT 1899.130 3164.490 1900.310 3165.670 ;
        RECT 1900.730 3164.490 1901.910 3165.670 ;
        RECT 1899.130 2986.090 1900.310 2987.270 ;
        RECT 1900.730 2986.090 1901.910 2987.270 ;
        RECT 1899.130 2984.490 1900.310 2985.670 ;
        RECT 1900.730 2984.490 1901.910 2985.670 ;
        RECT 1899.130 2806.090 1900.310 2807.270 ;
        RECT 1900.730 2806.090 1901.910 2807.270 ;
        RECT 1899.130 2804.490 1900.310 2805.670 ;
        RECT 1900.730 2804.490 1901.910 2805.670 ;
        RECT 1899.130 2626.090 1900.310 2627.270 ;
        RECT 1900.730 2626.090 1901.910 2627.270 ;
        RECT 1899.130 2624.490 1900.310 2625.670 ;
        RECT 1900.730 2624.490 1901.910 2625.670 ;
        RECT 1899.130 2446.090 1900.310 2447.270 ;
        RECT 1900.730 2446.090 1901.910 2447.270 ;
        RECT 1899.130 2444.490 1900.310 2445.670 ;
        RECT 1900.730 2444.490 1901.910 2445.670 ;
        RECT 1899.130 2266.090 1900.310 2267.270 ;
        RECT 1900.730 2266.090 1901.910 2267.270 ;
        RECT 1899.130 2264.490 1900.310 2265.670 ;
        RECT 1900.730 2264.490 1901.910 2265.670 ;
        RECT 1899.130 2086.090 1900.310 2087.270 ;
        RECT 1900.730 2086.090 1901.910 2087.270 ;
        RECT 1899.130 2084.490 1900.310 2085.670 ;
        RECT 1900.730 2084.490 1901.910 2085.670 ;
        RECT 1899.130 1906.090 1900.310 1907.270 ;
        RECT 1900.730 1906.090 1901.910 1907.270 ;
        RECT 1899.130 1904.490 1900.310 1905.670 ;
        RECT 1900.730 1904.490 1901.910 1905.670 ;
        RECT 1899.130 1726.090 1900.310 1727.270 ;
        RECT 1900.730 1726.090 1901.910 1727.270 ;
        RECT 1899.130 1724.490 1900.310 1725.670 ;
        RECT 1900.730 1724.490 1901.910 1725.670 ;
        RECT 1899.130 1546.090 1900.310 1547.270 ;
        RECT 1900.730 1546.090 1901.910 1547.270 ;
        RECT 1899.130 1544.490 1900.310 1545.670 ;
        RECT 1900.730 1544.490 1901.910 1545.670 ;
        RECT 1899.130 1366.090 1900.310 1367.270 ;
        RECT 1900.730 1366.090 1901.910 1367.270 ;
        RECT 1899.130 1364.490 1900.310 1365.670 ;
        RECT 1900.730 1364.490 1901.910 1365.670 ;
        RECT 1899.130 1186.090 1900.310 1187.270 ;
        RECT 1900.730 1186.090 1901.910 1187.270 ;
        RECT 1899.130 1184.490 1900.310 1185.670 ;
        RECT 1900.730 1184.490 1901.910 1185.670 ;
        RECT 1899.130 1006.090 1900.310 1007.270 ;
        RECT 1900.730 1006.090 1901.910 1007.270 ;
        RECT 1899.130 1004.490 1900.310 1005.670 ;
        RECT 1900.730 1004.490 1901.910 1005.670 ;
        RECT 1899.130 826.090 1900.310 827.270 ;
        RECT 1900.730 826.090 1901.910 827.270 ;
        RECT 1899.130 824.490 1900.310 825.670 ;
        RECT 1900.730 824.490 1901.910 825.670 ;
        RECT 1899.130 646.090 1900.310 647.270 ;
        RECT 1900.730 646.090 1901.910 647.270 ;
        RECT 1899.130 644.490 1900.310 645.670 ;
        RECT 1900.730 644.490 1901.910 645.670 ;
        RECT 1899.130 466.090 1900.310 467.270 ;
        RECT 1900.730 466.090 1901.910 467.270 ;
        RECT 1899.130 464.490 1900.310 465.670 ;
        RECT 1900.730 464.490 1901.910 465.670 ;
        RECT 1899.130 286.090 1900.310 287.270 ;
        RECT 1900.730 286.090 1901.910 287.270 ;
        RECT 1899.130 284.490 1900.310 285.670 ;
        RECT 1900.730 284.490 1901.910 285.670 ;
        RECT 1899.130 106.090 1900.310 107.270 ;
        RECT 1900.730 106.090 1901.910 107.270 ;
        RECT 1899.130 104.490 1900.310 105.670 ;
        RECT 1900.730 104.490 1901.910 105.670 ;
        RECT 1899.130 -7.710 1900.310 -6.530 ;
        RECT 1900.730 -7.710 1901.910 -6.530 ;
        RECT 1899.130 -9.310 1900.310 -8.130 ;
        RECT 1900.730 -9.310 1901.910 -8.130 ;
        RECT 2079.130 3527.810 2080.310 3528.990 ;
        RECT 2080.730 3527.810 2081.910 3528.990 ;
        RECT 2079.130 3526.210 2080.310 3527.390 ;
        RECT 2080.730 3526.210 2081.910 3527.390 ;
        RECT 2079.130 3346.090 2080.310 3347.270 ;
        RECT 2080.730 3346.090 2081.910 3347.270 ;
        RECT 2079.130 3344.490 2080.310 3345.670 ;
        RECT 2080.730 3344.490 2081.910 3345.670 ;
        RECT 2079.130 3166.090 2080.310 3167.270 ;
        RECT 2080.730 3166.090 2081.910 3167.270 ;
        RECT 2079.130 3164.490 2080.310 3165.670 ;
        RECT 2080.730 3164.490 2081.910 3165.670 ;
        RECT 2079.130 2986.090 2080.310 2987.270 ;
        RECT 2080.730 2986.090 2081.910 2987.270 ;
        RECT 2079.130 2984.490 2080.310 2985.670 ;
        RECT 2080.730 2984.490 2081.910 2985.670 ;
        RECT 2079.130 2806.090 2080.310 2807.270 ;
        RECT 2080.730 2806.090 2081.910 2807.270 ;
        RECT 2079.130 2804.490 2080.310 2805.670 ;
        RECT 2080.730 2804.490 2081.910 2805.670 ;
        RECT 2079.130 2626.090 2080.310 2627.270 ;
        RECT 2080.730 2626.090 2081.910 2627.270 ;
        RECT 2079.130 2624.490 2080.310 2625.670 ;
        RECT 2080.730 2624.490 2081.910 2625.670 ;
        RECT 2079.130 2446.090 2080.310 2447.270 ;
        RECT 2080.730 2446.090 2081.910 2447.270 ;
        RECT 2079.130 2444.490 2080.310 2445.670 ;
        RECT 2080.730 2444.490 2081.910 2445.670 ;
        RECT 2079.130 2266.090 2080.310 2267.270 ;
        RECT 2080.730 2266.090 2081.910 2267.270 ;
        RECT 2079.130 2264.490 2080.310 2265.670 ;
        RECT 2080.730 2264.490 2081.910 2265.670 ;
        RECT 2079.130 2086.090 2080.310 2087.270 ;
        RECT 2080.730 2086.090 2081.910 2087.270 ;
        RECT 2079.130 2084.490 2080.310 2085.670 ;
        RECT 2080.730 2084.490 2081.910 2085.670 ;
        RECT 2079.130 1906.090 2080.310 1907.270 ;
        RECT 2080.730 1906.090 2081.910 1907.270 ;
        RECT 2079.130 1904.490 2080.310 1905.670 ;
        RECT 2080.730 1904.490 2081.910 1905.670 ;
        RECT 2079.130 1726.090 2080.310 1727.270 ;
        RECT 2080.730 1726.090 2081.910 1727.270 ;
        RECT 2079.130 1724.490 2080.310 1725.670 ;
        RECT 2080.730 1724.490 2081.910 1725.670 ;
        RECT 2079.130 1546.090 2080.310 1547.270 ;
        RECT 2080.730 1546.090 2081.910 1547.270 ;
        RECT 2079.130 1544.490 2080.310 1545.670 ;
        RECT 2080.730 1544.490 2081.910 1545.670 ;
        RECT 2079.130 1366.090 2080.310 1367.270 ;
        RECT 2080.730 1366.090 2081.910 1367.270 ;
        RECT 2079.130 1364.490 2080.310 1365.670 ;
        RECT 2080.730 1364.490 2081.910 1365.670 ;
        RECT 2079.130 1186.090 2080.310 1187.270 ;
        RECT 2080.730 1186.090 2081.910 1187.270 ;
        RECT 2079.130 1184.490 2080.310 1185.670 ;
        RECT 2080.730 1184.490 2081.910 1185.670 ;
        RECT 2079.130 1006.090 2080.310 1007.270 ;
        RECT 2080.730 1006.090 2081.910 1007.270 ;
        RECT 2079.130 1004.490 2080.310 1005.670 ;
        RECT 2080.730 1004.490 2081.910 1005.670 ;
        RECT 2079.130 826.090 2080.310 827.270 ;
        RECT 2080.730 826.090 2081.910 827.270 ;
        RECT 2079.130 824.490 2080.310 825.670 ;
        RECT 2080.730 824.490 2081.910 825.670 ;
        RECT 2079.130 646.090 2080.310 647.270 ;
        RECT 2080.730 646.090 2081.910 647.270 ;
        RECT 2079.130 644.490 2080.310 645.670 ;
        RECT 2080.730 644.490 2081.910 645.670 ;
        RECT 2079.130 466.090 2080.310 467.270 ;
        RECT 2080.730 466.090 2081.910 467.270 ;
        RECT 2079.130 464.490 2080.310 465.670 ;
        RECT 2080.730 464.490 2081.910 465.670 ;
        RECT 2079.130 286.090 2080.310 287.270 ;
        RECT 2080.730 286.090 2081.910 287.270 ;
        RECT 2079.130 284.490 2080.310 285.670 ;
        RECT 2080.730 284.490 2081.910 285.670 ;
        RECT 2079.130 106.090 2080.310 107.270 ;
        RECT 2080.730 106.090 2081.910 107.270 ;
        RECT 2079.130 104.490 2080.310 105.670 ;
        RECT 2080.730 104.490 2081.910 105.670 ;
        RECT 2079.130 -7.710 2080.310 -6.530 ;
        RECT 2080.730 -7.710 2081.910 -6.530 ;
        RECT 2079.130 -9.310 2080.310 -8.130 ;
        RECT 2080.730 -9.310 2081.910 -8.130 ;
        RECT 2259.130 3527.810 2260.310 3528.990 ;
        RECT 2260.730 3527.810 2261.910 3528.990 ;
        RECT 2259.130 3526.210 2260.310 3527.390 ;
        RECT 2260.730 3526.210 2261.910 3527.390 ;
        RECT 2259.130 3346.090 2260.310 3347.270 ;
        RECT 2260.730 3346.090 2261.910 3347.270 ;
        RECT 2259.130 3344.490 2260.310 3345.670 ;
        RECT 2260.730 3344.490 2261.910 3345.670 ;
        RECT 2259.130 3166.090 2260.310 3167.270 ;
        RECT 2260.730 3166.090 2261.910 3167.270 ;
        RECT 2259.130 3164.490 2260.310 3165.670 ;
        RECT 2260.730 3164.490 2261.910 3165.670 ;
        RECT 2259.130 2986.090 2260.310 2987.270 ;
        RECT 2260.730 2986.090 2261.910 2987.270 ;
        RECT 2259.130 2984.490 2260.310 2985.670 ;
        RECT 2260.730 2984.490 2261.910 2985.670 ;
        RECT 2259.130 2806.090 2260.310 2807.270 ;
        RECT 2260.730 2806.090 2261.910 2807.270 ;
        RECT 2259.130 2804.490 2260.310 2805.670 ;
        RECT 2260.730 2804.490 2261.910 2805.670 ;
        RECT 2259.130 2626.090 2260.310 2627.270 ;
        RECT 2260.730 2626.090 2261.910 2627.270 ;
        RECT 2259.130 2624.490 2260.310 2625.670 ;
        RECT 2260.730 2624.490 2261.910 2625.670 ;
        RECT 2259.130 2446.090 2260.310 2447.270 ;
        RECT 2260.730 2446.090 2261.910 2447.270 ;
        RECT 2259.130 2444.490 2260.310 2445.670 ;
        RECT 2260.730 2444.490 2261.910 2445.670 ;
        RECT 2259.130 2266.090 2260.310 2267.270 ;
        RECT 2260.730 2266.090 2261.910 2267.270 ;
        RECT 2259.130 2264.490 2260.310 2265.670 ;
        RECT 2260.730 2264.490 2261.910 2265.670 ;
        RECT 2259.130 2086.090 2260.310 2087.270 ;
        RECT 2260.730 2086.090 2261.910 2087.270 ;
        RECT 2259.130 2084.490 2260.310 2085.670 ;
        RECT 2260.730 2084.490 2261.910 2085.670 ;
        RECT 2259.130 1906.090 2260.310 1907.270 ;
        RECT 2260.730 1906.090 2261.910 1907.270 ;
        RECT 2259.130 1904.490 2260.310 1905.670 ;
        RECT 2260.730 1904.490 2261.910 1905.670 ;
        RECT 2259.130 1726.090 2260.310 1727.270 ;
        RECT 2260.730 1726.090 2261.910 1727.270 ;
        RECT 2259.130 1724.490 2260.310 1725.670 ;
        RECT 2260.730 1724.490 2261.910 1725.670 ;
        RECT 2259.130 1546.090 2260.310 1547.270 ;
        RECT 2260.730 1546.090 2261.910 1547.270 ;
        RECT 2259.130 1544.490 2260.310 1545.670 ;
        RECT 2260.730 1544.490 2261.910 1545.670 ;
        RECT 2259.130 1366.090 2260.310 1367.270 ;
        RECT 2260.730 1366.090 2261.910 1367.270 ;
        RECT 2259.130 1364.490 2260.310 1365.670 ;
        RECT 2260.730 1364.490 2261.910 1365.670 ;
        RECT 2259.130 1186.090 2260.310 1187.270 ;
        RECT 2260.730 1186.090 2261.910 1187.270 ;
        RECT 2259.130 1184.490 2260.310 1185.670 ;
        RECT 2260.730 1184.490 2261.910 1185.670 ;
        RECT 2259.130 1006.090 2260.310 1007.270 ;
        RECT 2260.730 1006.090 2261.910 1007.270 ;
        RECT 2259.130 1004.490 2260.310 1005.670 ;
        RECT 2260.730 1004.490 2261.910 1005.670 ;
        RECT 2259.130 826.090 2260.310 827.270 ;
        RECT 2260.730 826.090 2261.910 827.270 ;
        RECT 2259.130 824.490 2260.310 825.670 ;
        RECT 2260.730 824.490 2261.910 825.670 ;
        RECT 2259.130 646.090 2260.310 647.270 ;
        RECT 2260.730 646.090 2261.910 647.270 ;
        RECT 2259.130 644.490 2260.310 645.670 ;
        RECT 2260.730 644.490 2261.910 645.670 ;
        RECT 2259.130 466.090 2260.310 467.270 ;
        RECT 2260.730 466.090 2261.910 467.270 ;
        RECT 2259.130 464.490 2260.310 465.670 ;
        RECT 2260.730 464.490 2261.910 465.670 ;
        RECT 2259.130 286.090 2260.310 287.270 ;
        RECT 2260.730 286.090 2261.910 287.270 ;
        RECT 2259.130 284.490 2260.310 285.670 ;
        RECT 2260.730 284.490 2261.910 285.670 ;
        RECT 2259.130 106.090 2260.310 107.270 ;
        RECT 2260.730 106.090 2261.910 107.270 ;
        RECT 2259.130 104.490 2260.310 105.670 ;
        RECT 2260.730 104.490 2261.910 105.670 ;
        RECT 2259.130 -7.710 2260.310 -6.530 ;
        RECT 2260.730 -7.710 2261.910 -6.530 ;
        RECT 2259.130 -9.310 2260.310 -8.130 ;
        RECT 2260.730 -9.310 2261.910 -8.130 ;
        RECT 2439.130 3527.810 2440.310 3528.990 ;
        RECT 2440.730 3527.810 2441.910 3528.990 ;
        RECT 2439.130 3526.210 2440.310 3527.390 ;
        RECT 2440.730 3526.210 2441.910 3527.390 ;
        RECT 2439.130 3346.090 2440.310 3347.270 ;
        RECT 2440.730 3346.090 2441.910 3347.270 ;
        RECT 2439.130 3344.490 2440.310 3345.670 ;
        RECT 2440.730 3344.490 2441.910 3345.670 ;
        RECT 2439.130 3166.090 2440.310 3167.270 ;
        RECT 2440.730 3166.090 2441.910 3167.270 ;
        RECT 2439.130 3164.490 2440.310 3165.670 ;
        RECT 2440.730 3164.490 2441.910 3165.670 ;
        RECT 2439.130 2986.090 2440.310 2987.270 ;
        RECT 2440.730 2986.090 2441.910 2987.270 ;
        RECT 2439.130 2984.490 2440.310 2985.670 ;
        RECT 2440.730 2984.490 2441.910 2985.670 ;
        RECT 2439.130 2806.090 2440.310 2807.270 ;
        RECT 2440.730 2806.090 2441.910 2807.270 ;
        RECT 2439.130 2804.490 2440.310 2805.670 ;
        RECT 2440.730 2804.490 2441.910 2805.670 ;
        RECT 2439.130 2626.090 2440.310 2627.270 ;
        RECT 2440.730 2626.090 2441.910 2627.270 ;
        RECT 2439.130 2624.490 2440.310 2625.670 ;
        RECT 2440.730 2624.490 2441.910 2625.670 ;
        RECT 2439.130 2446.090 2440.310 2447.270 ;
        RECT 2440.730 2446.090 2441.910 2447.270 ;
        RECT 2439.130 2444.490 2440.310 2445.670 ;
        RECT 2440.730 2444.490 2441.910 2445.670 ;
        RECT 2439.130 2266.090 2440.310 2267.270 ;
        RECT 2440.730 2266.090 2441.910 2267.270 ;
        RECT 2439.130 2264.490 2440.310 2265.670 ;
        RECT 2440.730 2264.490 2441.910 2265.670 ;
        RECT 2439.130 2086.090 2440.310 2087.270 ;
        RECT 2440.730 2086.090 2441.910 2087.270 ;
        RECT 2439.130 2084.490 2440.310 2085.670 ;
        RECT 2440.730 2084.490 2441.910 2085.670 ;
        RECT 2439.130 1906.090 2440.310 1907.270 ;
        RECT 2440.730 1906.090 2441.910 1907.270 ;
        RECT 2439.130 1904.490 2440.310 1905.670 ;
        RECT 2440.730 1904.490 2441.910 1905.670 ;
        RECT 2439.130 1726.090 2440.310 1727.270 ;
        RECT 2440.730 1726.090 2441.910 1727.270 ;
        RECT 2439.130 1724.490 2440.310 1725.670 ;
        RECT 2440.730 1724.490 2441.910 1725.670 ;
        RECT 2439.130 1546.090 2440.310 1547.270 ;
        RECT 2440.730 1546.090 2441.910 1547.270 ;
        RECT 2439.130 1544.490 2440.310 1545.670 ;
        RECT 2440.730 1544.490 2441.910 1545.670 ;
        RECT 2439.130 1366.090 2440.310 1367.270 ;
        RECT 2440.730 1366.090 2441.910 1367.270 ;
        RECT 2439.130 1364.490 2440.310 1365.670 ;
        RECT 2440.730 1364.490 2441.910 1365.670 ;
        RECT 2439.130 1186.090 2440.310 1187.270 ;
        RECT 2440.730 1186.090 2441.910 1187.270 ;
        RECT 2439.130 1184.490 2440.310 1185.670 ;
        RECT 2440.730 1184.490 2441.910 1185.670 ;
        RECT 2439.130 1006.090 2440.310 1007.270 ;
        RECT 2440.730 1006.090 2441.910 1007.270 ;
        RECT 2439.130 1004.490 2440.310 1005.670 ;
        RECT 2440.730 1004.490 2441.910 1005.670 ;
        RECT 2439.130 826.090 2440.310 827.270 ;
        RECT 2440.730 826.090 2441.910 827.270 ;
        RECT 2439.130 824.490 2440.310 825.670 ;
        RECT 2440.730 824.490 2441.910 825.670 ;
        RECT 2439.130 646.090 2440.310 647.270 ;
        RECT 2440.730 646.090 2441.910 647.270 ;
        RECT 2439.130 644.490 2440.310 645.670 ;
        RECT 2440.730 644.490 2441.910 645.670 ;
        RECT 2439.130 466.090 2440.310 467.270 ;
        RECT 2440.730 466.090 2441.910 467.270 ;
        RECT 2439.130 464.490 2440.310 465.670 ;
        RECT 2440.730 464.490 2441.910 465.670 ;
        RECT 2439.130 286.090 2440.310 287.270 ;
        RECT 2440.730 286.090 2441.910 287.270 ;
        RECT 2439.130 284.490 2440.310 285.670 ;
        RECT 2440.730 284.490 2441.910 285.670 ;
        RECT 2439.130 106.090 2440.310 107.270 ;
        RECT 2440.730 106.090 2441.910 107.270 ;
        RECT 2439.130 104.490 2440.310 105.670 ;
        RECT 2440.730 104.490 2441.910 105.670 ;
        RECT 2439.130 -7.710 2440.310 -6.530 ;
        RECT 2440.730 -7.710 2441.910 -6.530 ;
        RECT 2439.130 -9.310 2440.310 -8.130 ;
        RECT 2440.730 -9.310 2441.910 -8.130 ;
        RECT 2619.130 3527.810 2620.310 3528.990 ;
        RECT 2620.730 3527.810 2621.910 3528.990 ;
        RECT 2619.130 3526.210 2620.310 3527.390 ;
        RECT 2620.730 3526.210 2621.910 3527.390 ;
        RECT 2619.130 3346.090 2620.310 3347.270 ;
        RECT 2620.730 3346.090 2621.910 3347.270 ;
        RECT 2619.130 3344.490 2620.310 3345.670 ;
        RECT 2620.730 3344.490 2621.910 3345.670 ;
        RECT 2619.130 3166.090 2620.310 3167.270 ;
        RECT 2620.730 3166.090 2621.910 3167.270 ;
        RECT 2619.130 3164.490 2620.310 3165.670 ;
        RECT 2620.730 3164.490 2621.910 3165.670 ;
        RECT 2619.130 2986.090 2620.310 2987.270 ;
        RECT 2620.730 2986.090 2621.910 2987.270 ;
        RECT 2619.130 2984.490 2620.310 2985.670 ;
        RECT 2620.730 2984.490 2621.910 2985.670 ;
        RECT 2619.130 2806.090 2620.310 2807.270 ;
        RECT 2620.730 2806.090 2621.910 2807.270 ;
        RECT 2619.130 2804.490 2620.310 2805.670 ;
        RECT 2620.730 2804.490 2621.910 2805.670 ;
        RECT 2619.130 2626.090 2620.310 2627.270 ;
        RECT 2620.730 2626.090 2621.910 2627.270 ;
        RECT 2619.130 2624.490 2620.310 2625.670 ;
        RECT 2620.730 2624.490 2621.910 2625.670 ;
        RECT 2619.130 2446.090 2620.310 2447.270 ;
        RECT 2620.730 2446.090 2621.910 2447.270 ;
        RECT 2619.130 2444.490 2620.310 2445.670 ;
        RECT 2620.730 2444.490 2621.910 2445.670 ;
        RECT 2619.130 2266.090 2620.310 2267.270 ;
        RECT 2620.730 2266.090 2621.910 2267.270 ;
        RECT 2619.130 2264.490 2620.310 2265.670 ;
        RECT 2620.730 2264.490 2621.910 2265.670 ;
        RECT 2619.130 2086.090 2620.310 2087.270 ;
        RECT 2620.730 2086.090 2621.910 2087.270 ;
        RECT 2619.130 2084.490 2620.310 2085.670 ;
        RECT 2620.730 2084.490 2621.910 2085.670 ;
        RECT 2619.130 1906.090 2620.310 1907.270 ;
        RECT 2620.730 1906.090 2621.910 1907.270 ;
        RECT 2619.130 1904.490 2620.310 1905.670 ;
        RECT 2620.730 1904.490 2621.910 1905.670 ;
        RECT 2619.130 1726.090 2620.310 1727.270 ;
        RECT 2620.730 1726.090 2621.910 1727.270 ;
        RECT 2619.130 1724.490 2620.310 1725.670 ;
        RECT 2620.730 1724.490 2621.910 1725.670 ;
        RECT 2619.130 1546.090 2620.310 1547.270 ;
        RECT 2620.730 1546.090 2621.910 1547.270 ;
        RECT 2619.130 1544.490 2620.310 1545.670 ;
        RECT 2620.730 1544.490 2621.910 1545.670 ;
        RECT 2619.130 1366.090 2620.310 1367.270 ;
        RECT 2620.730 1366.090 2621.910 1367.270 ;
        RECT 2619.130 1364.490 2620.310 1365.670 ;
        RECT 2620.730 1364.490 2621.910 1365.670 ;
        RECT 2619.130 1186.090 2620.310 1187.270 ;
        RECT 2620.730 1186.090 2621.910 1187.270 ;
        RECT 2619.130 1184.490 2620.310 1185.670 ;
        RECT 2620.730 1184.490 2621.910 1185.670 ;
        RECT 2619.130 1006.090 2620.310 1007.270 ;
        RECT 2620.730 1006.090 2621.910 1007.270 ;
        RECT 2619.130 1004.490 2620.310 1005.670 ;
        RECT 2620.730 1004.490 2621.910 1005.670 ;
        RECT 2619.130 826.090 2620.310 827.270 ;
        RECT 2620.730 826.090 2621.910 827.270 ;
        RECT 2619.130 824.490 2620.310 825.670 ;
        RECT 2620.730 824.490 2621.910 825.670 ;
        RECT 2619.130 646.090 2620.310 647.270 ;
        RECT 2620.730 646.090 2621.910 647.270 ;
        RECT 2619.130 644.490 2620.310 645.670 ;
        RECT 2620.730 644.490 2621.910 645.670 ;
        RECT 2619.130 466.090 2620.310 467.270 ;
        RECT 2620.730 466.090 2621.910 467.270 ;
        RECT 2619.130 464.490 2620.310 465.670 ;
        RECT 2620.730 464.490 2621.910 465.670 ;
        RECT 2619.130 286.090 2620.310 287.270 ;
        RECT 2620.730 286.090 2621.910 287.270 ;
        RECT 2619.130 284.490 2620.310 285.670 ;
        RECT 2620.730 284.490 2621.910 285.670 ;
        RECT 2619.130 106.090 2620.310 107.270 ;
        RECT 2620.730 106.090 2621.910 107.270 ;
        RECT 2619.130 104.490 2620.310 105.670 ;
        RECT 2620.730 104.490 2621.910 105.670 ;
        RECT 2619.130 -7.710 2620.310 -6.530 ;
        RECT 2620.730 -7.710 2621.910 -6.530 ;
        RECT 2619.130 -9.310 2620.310 -8.130 ;
        RECT 2620.730 -9.310 2621.910 -8.130 ;
        RECT 2799.130 3527.810 2800.310 3528.990 ;
        RECT 2800.730 3527.810 2801.910 3528.990 ;
        RECT 2799.130 3526.210 2800.310 3527.390 ;
        RECT 2800.730 3526.210 2801.910 3527.390 ;
        RECT 2799.130 3346.090 2800.310 3347.270 ;
        RECT 2800.730 3346.090 2801.910 3347.270 ;
        RECT 2799.130 3344.490 2800.310 3345.670 ;
        RECT 2800.730 3344.490 2801.910 3345.670 ;
        RECT 2799.130 3166.090 2800.310 3167.270 ;
        RECT 2800.730 3166.090 2801.910 3167.270 ;
        RECT 2799.130 3164.490 2800.310 3165.670 ;
        RECT 2800.730 3164.490 2801.910 3165.670 ;
        RECT 2799.130 2986.090 2800.310 2987.270 ;
        RECT 2800.730 2986.090 2801.910 2987.270 ;
        RECT 2799.130 2984.490 2800.310 2985.670 ;
        RECT 2800.730 2984.490 2801.910 2985.670 ;
        RECT 2799.130 2806.090 2800.310 2807.270 ;
        RECT 2800.730 2806.090 2801.910 2807.270 ;
        RECT 2799.130 2804.490 2800.310 2805.670 ;
        RECT 2800.730 2804.490 2801.910 2805.670 ;
        RECT 2799.130 2626.090 2800.310 2627.270 ;
        RECT 2800.730 2626.090 2801.910 2627.270 ;
        RECT 2799.130 2624.490 2800.310 2625.670 ;
        RECT 2800.730 2624.490 2801.910 2625.670 ;
        RECT 2799.130 2446.090 2800.310 2447.270 ;
        RECT 2800.730 2446.090 2801.910 2447.270 ;
        RECT 2799.130 2444.490 2800.310 2445.670 ;
        RECT 2800.730 2444.490 2801.910 2445.670 ;
        RECT 2799.130 2266.090 2800.310 2267.270 ;
        RECT 2800.730 2266.090 2801.910 2267.270 ;
        RECT 2799.130 2264.490 2800.310 2265.670 ;
        RECT 2800.730 2264.490 2801.910 2265.670 ;
        RECT 2799.130 2086.090 2800.310 2087.270 ;
        RECT 2800.730 2086.090 2801.910 2087.270 ;
        RECT 2799.130 2084.490 2800.310 2085.670 ;
        RECT 2800.730 2084.490 2801.910 2085.670 ;
        RECT 2799.130 1906.090 2800.310 1907.270 ;
        RECT 2800.730 1906.090 2801.910 1907.270 ;
        RECT 2799.130 1904.490 2800.310 1905.670 ;
        RECT 2800.730 1904.490 2801.910 1905.670 ;
        RECT 2799.130 1726.090 2800.310 1727.270 ;
        RECT 2800.730 1726.090 2801.910 1727.270 ;
        RECT 2799.130 1724.490 2800.310 1725.670 ;
        RECT 2800.730 1724.490 2801.910 1725.670 ;
        RECT 2799.130 1546.090 2800.310 1547.270 ;
        RECT 2800.730 1546.090 2801.910 1547.270 ;
        RECT 2799.130 1544.490 2800.310 1545.670 ;
        RECT 2800.730 1544.490 2801.910 1545.670 ;
        RECT 2799.130 1366.090 2800.310 1367.270 ;
        RECT 2800.730 1366.090 2801.910 1367.270 ;
        RECT 2799.130 1364.490 2800.310 1365.670 ;
        RECT 2800.730 1364.490 2801.910 1365.670 ;
        RECT 2799.130 1186.090 2800.310 1187.270 ;
        RECT 2800.730 1186.090 2801.910 1187.270 ;
        RECT 2799.130 1184.490 2800.310 1185.670 ;
        RECT 2800.730 1184.490 2801.910 1185.670 ;
        RECT 2799.130 1006.090 2800.310 1007.270 ;
        RECT 2800.730 1006.090 2801.910 1007.270 ;
        RECT 2799.130 1004.490 2800.310 1005.670 ;
        RECT 2800.730 1004.490 2801.910 1005.670 ;
        RECT 2799.130 826.090 2800.310 827.270 ;
        RECT 2800.730 826.090 2801.910 827.270 ;
        RECT 2799.130 824.490 2800.310 825.670 ;
        RECT 2800.730 824.490 2801.910 825.670 ;
        RECT 2799.130 646.090 2800.310 647.270 ;
        RECT 2800.730 646.090 2801.910 647.270 ;
        RECT 2799.130 644.490 2800.310 645.670 ;
        RECT 2800.730 644.490 2801.910 645.670 ;
        RECT 2799.130 466.090 2800.310 467.270 ;
        RECT 2800.730 466.090 2801.910 467.270 ;
        RECT 2799.130 464.490 2800.310 465.670 ;
        RECT 2800.730 464.490 2801.910 465.670 ;
        RECT 2799.130 286.090 2800.310 287.270 ;
        RECT 2800.730 286.090 2801.910 287.270 ;
        RECT 2799.130 284.490 2800.310 285.670 ;
        RECT 2800.730 284.490 2801.910 285.670 ;
        RECT 2799.130 106.090 2800.310 107.270 ;
        RECT 2800.730 106.090 2801.910 107.270 ;
        RECT 2799.130 104.490 2800.310 105.670 ;
        RECT 2800.730 104.490 2801.910 105.670 ;
        RECT 2799.130 -7.710 2800.310 -6.530 ;
        RECT 2800.730 -7.710 2801.910 -6.530 ;
        RECT 2799.130 -9.310 2800.310 -8.130 ;
        RECT 2800.730 -9.310 2801.910 -8.130 ;
        RECT 2931.510 3527.810 2932.690 3528.990 ;
        RECT 2933.110 3527.810 2934.290 3528.990 ;
        RECT 2931.510 3526.210 2932.690 3527.390 ;
        RECT 2933.110 3526.210 2934.290 3527.390 ;
        RECT 2931.510 3346.090 2932.690 3347.270 ;
        RECT 2933.110 3346.090 2934.290 3347.270 ;
        RECT 2931.510 3344.490 2932.690 3345.670 ;
        RECT 2933.110 3344.490 2934.290 3345.670 ;
        RECT 2931.510 3166.090 2932.690 3167.270 ;
        RECT 2933.110 3166.090 2934.290 3167.270 ;
        RECT 2931.510 3164.490 2932.690 3165.670 ;
        RECT 2933.110 3164.490 2934.290 3165.670 ;
        RECT 2931.510 2986.090 2932.690 2987.270 ;
        RECT 2933.110 2986.090 2934.290 2987.270 ;
        RECT 2931.510 2984.490 2932.690 2985.670 ;
        RECT 2933.110 2984.490 2934.290 2985.670 ;
        RECT 2931.510 2806.090 2932.690 2807.270 ;
        RECT 2933.110 2806.090 2934.290 2807.270 ;
        RECT 2931.510 2804.490 2932.690 2805.670 ;
        RECT 2933.110 2804.490 2934.290 2805.670 ;
        RECT 2931.510 2626.090 2932.690 2627.270 ;
        RECT 2933.110 2626.090 2934.290 2627.270 ;
        RECT 2931.510 2624.490 2932.690 2625.670 ;
        RECT 2933.110 2624.490 2934.290 2625.670 ;
        RECT 2931.510 2446.090 2932.690 2447.270 ;
        RECT 2933.110 2446.090 2934.290 2447.270 ;
        RECT 2931.510 2444.490 2932.690 2445.670 ;
        RECT 2933.110 2444.490 2934.290 2445.670 ;
        RECT 2931.510 2266.090 2932.690 2267.270 ;
        RECT 2933.110 2266.090 2934.290 2267.270 ;
        RECT 2931.510 2264.490 2932.690 2265.670 ;
        RECT 2933.110 2264.490 2934.290 2265.670 ;
        RECT 2931.510 2086.090 2932.690 2087.270 ;
        RECT 2933.110 2086.090 2934.290 2087.270 ;
        RECT 2931.510 2084.490 2932.690 2085.670 ;
        RECT 2933.110 2084.490 2934.290 2085.670 ;
        RECT 2931.510 1906.090 2932.690 1907.270 ;
        RECT 2933.110 1906.090 2934.290 1907.270 ;
        RECT 2931.510 1904.490 2932.690 1905.670 ;
        RECT 2933.110 1904.490 2934.290 1905.670 ;
        RECT 2931.510 1726.090 2932.690 1727.270 ;
        RECT 2933.110 1726.090 2934.290 1727.270 ;
        RECT 2931.510 1724.490 2932.690 1725.670 ;
        RECT 2933.110 1724.490 2934.290 1725.670 ;
        RECT 2931.510 1546.090 2932.690 1547.270 ;
        RECT 2933.110 1546.090 2934.290 1547.270 ;
        RECT 2931.510 1544.490 2932.690 1545.670 ;
        RECT 2933.110 1544.490 2934.290 1545.670 ;
        RECT 2931.510 1366.090 2932.690 1367.270 ;
        RECT 2933.110 1366.090 2934.290 1367.270 ;
        RECT 2931.510 1364.490 2932.690 1365.670 ;
        RECT 2933.110 1364.490 2934.290 1365.670 ;
        RECT 2931.510 1186.090 2932.690 1187.270 ;
        RECT 2933.110 1186.090 2934.290 1187.270 ;
        RECT 2931.510 1184.490 2932.690 1185.670 ;
        RECT 2933.110 1184.490 2934.290 1185.670 ;
        RECT 2931.510 1006.090 2932.690 1007.270 ;
        RECT 2933.110 1006.090 2934.290 1007.270 ;
        RECT 2931.510 1004.490 2932.690 1005.670 ;
        RECT 2933.110 1004.490 2934.290 1005.670 ;
        RECT 2931.510 826.090 2932.690 827.270 ;
        RECT 2933.110 826.090 2934.290 827.270 ;
        RECT 2931.510 824.490 2932.690 825.670 ;
        RECT 2933.110 824.490 2934.290 825.670 ;
        RECT 2931.510 646.090 2932.690 647.270 ;
        RECT 2933.110 646.090 2934.290 647.270 ;
        RECT 2931.510 644.490 2932.690 645.670 ;
        RECT 2933.110 644.490 2934.290 645.670 ;
        RECT 2931.510 466.090 2932.690 467.270 ;
        RECT 2933.110 466.090 2934.290 467.270 ;
        RECT 2931.510 464.490 2932.690 465.670 ;
        RECT 2933.110 464.490 2934.290 465.670 ;
        RECT 2931.510 286.090 2932.690 287.270 ;
        RECT 2933.110 286.090 2934.290 287.270 ;
        RECT 2931.510 284.490 2932.690 285.670 ;
        RECT 2933.110 284.490 2934.290 285.670 ;
        RECT 2931.510 106.090 2932.690 107.270 ;
        RECT 2933.110 106.090 2934.290 107.270 ;
        RECT 2931.510 104.490 2932.690 105.670 ;
        RECT 2933.110 104.490 2934.290 105.670 ;
        RECT 2931.510 -7.710 2932.690 -6.530 ;
        RECT 2933.110 -7.710 2934.290 -6.530 ;
        RECT 2931.510 -9.310 2932.690 -8.130 ;
        RECT 2933.110 -9.310 2934.290 -8.130 ;
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
        RECT -14.830 3344.330 2934.450 3347.430 ;
        RECT -14.830 3164.330 2934.450 3167.430 ;
        RECT -14.830 2984.330 2934.450 2987.430 ;
        RECT -14.830 2804.330 2934.450 2807.430 ;
        RECT -14.830 2624.330 2934.450 2627.430 ;
        RECT -14.830 2444.330 2934.450 2447.430 ;
        RECT -14.830 2264.330 2934.450 2267.430 ;
        RECT -14.830 2084.330 2934.450 2087.430 ;
        RECT -14.830 1904.330 2934.450 1907.430 ;
        RECT -14.830 1724.330 2934.450 1727.430 ;
        RECT -14.830 1544.330 2934.450 1547.430 ;
        RECT -14.830 1364.330 2934.450 1367.430 ;
        RECT -14.830 1184.330 2934.450 1187.430 ;
        RECT -14.830 1004.330 2934.450 1007.430 ;
        RECT -14.830 824.330 2934.450 827.430 ;
        RECT -14.830 644.330 2934.450 647.430 ;
        RECT -14.830 464.330 2934.450 467.430 ;
        RECT -14.830 284.330 2934.450 287.430 ;
        RECT -14.830 104.330 2934.450 107.430 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
        RECT 297.570 1010.000 300.670 3538.750 ;
        RECT 477.570 1010.000 480.670 3538.750 ;
        RECT 657.570 1010.000 660.670 3538.750 ;
        RECT 837.570 1010.000 840.670 3538.750 ;
        RECT 1017.570 1010.000 1020.670 3538.750 ;
        RECT 297.570 -19.070 300.670 390.000 ;
        RECT 477.570 -19.070 480.670 390.000 ;
        RECT 657.570 -19.070 660.670 390.000 ;
        RECT 837.570 -19.070 840.670 390.000 ;
        RECT 1017.570 -19.070 1020.670 390.000 ;
        RECT 1197.570 -19.070 1200.670 3538.750 ;
        RECT 1377.570 -19.070 1380.670 3538.750 ;
        RECT 1557.570 -19.070 1560.670 3538.750 ;
        RECT 1737.570 -19.070 1740.670 3538.750 ;
        RECT 1917.570 -19.070 1920.670 3538.750 ;
        RECT 2097.570 -19.070 2100.670 3538.750 ;
        RECT 2277.570 -19.070 2280.670 3538.750 ;
        RECT 2457.570 -19.070 2460.670 3538.750 ;
        RECT 2637.570 -19.070 2640.670 3538.750 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
      LAYER via4 ;
        RECT -24.270 3537.410 -23.090 3538.590 ;
        RECT -22.670 3537.410 -21.490 3538.590 ;
        RECT -24.270 3535.810 -23.090 3536.990 ;
        RECT -22.670 3535.810 -21.490 3536.990 ;
        RECT -24.270 3364.690 -23.090 3365.870 ;
        RECT -22.670 3364.690 -21.490 3365.870 ;
        RECT -24.270 3363.090 -23.090 3364.270 ;
        RECT -22.670 3363.090 -21.490 3364.270 ;
        RECT -24.270 3184.690 -23.090 3185.870 ;
        RECT -22.670 3184.690 -21.490 3185.870 ;
        RECT -24.270 3183.090 -23.090 3184.270 ;
        RECT -22.670 3183.090 -21.490 3184.270 ;
        RECT -24.270 3004.690 -23.090 3005.870 ;
        RECT -22.670 3004.690 -21.490 3005.870 ;
        RECT -24.270 3003.090 -23.090 3004.270 ;
        RECT -22.670 3003.090 -21.490 3004.270 ;
        RECT -24.270 2824.690 -23.090 2825.870 ;
        RECT -22.670 2824.690 -21.490 2825.870 ;
        RECT -24.270 2823.090 -23.090 2824.270 ;
        RECT -22.670 2823.090 -21.490 2824.270 ;
        RECT -24.270 2644.690 -23.090 2645.870 ;
        RECT -22.670 2644.690 -21.490 2645.870 ;
        RECT -24.270 2643.090 -23.090 2644.270 ;
        RECT -22.670 2643.090 -21.490 2644.270 ;
        RECT -24.270 2464.690 -23.090 2465.870 ;
        RECT -22.670 2464.690 -21.490 2465.870 ;
        RECT -24.270 2463.090 -23.090 2464.270 ;
        RECT -22.670 2463.090 -21.490 2464.270 ;
        RECT -24.270 2284.690 -23.090 2285.870 ;
        RECT -22.670 2284.690 -21.490 2285.870 ;
        RECT -24.270 2283.090 -23.090 2284.270 ;
        RECT -22.670 2283.090 -21.490 2284.270 ;
        RECT -24.270 2104.690 -23.090 2105.870 ;
        RECT -22.670 2104.690 -21.490 2105.870 ;
        RECT -24.270 2103.090 -23.090 2104.270 ;
        RECT -22.670 2103.090 -21.490 2104.270 ;
        RECT -24.270 1924.690 -23.090 1925.870 ;
        RECT -22.670 1924.690 -21.490 1925.870 ;
        RECT -24.270 1923.090 -23.090 1924.270 ;
        RECT -22.670 1923.090 -21.490 1924.270 ;
        RECT -24.270 1744.690 -23.090 1745.870 ;
        RECT -22.670 1744.690 -21.490 1745.870 ;
        RECT -24.270 1743.090 -23.090 1744.270 ;
        RECT -22.670 1743.090 -21.490 1744.270 ;
        RECT -24.270 1564.690 -23.090 1565.870 ;
        RECT -22.670 1564.690 -21.490 1565.870 ;
        RECT -24.270 1563.090 -23.090 1564.270 ;
        RECT -22.670 1563.090 -21.490 1564.270 ;
        RECT -24.270 1384.690 -23.090 1385.870 ;
        RECT -22.670 1384.690 -21.490 1385.870 ;
        RECT -24.270 1383.090 -23.090 1384.270 ;
        RECT -22.670 1383.090 -21.490 1384.270 ;
        RECT -24.270 1204.690 -23.090 1205.870 ;
        RECT -22.670 1204.690 -21.490 1205.870 ;
        RECT -24.270 1203.090 -23.090 1204.270 ;
        RECT -22.670 1203.090 -21.490 1204.270 ;
        RECT -24.270 1024.690 -23.090 1025.870 ;
        RECT -22.670 1024.690 -21.490 1025.870 ;
        RECT -24.270 1023.090 -23.090 1024.270 ;
        RECT -22.670 1023.090 -21.490 1024.270 ;
        RECT -24.270 844.690 -23.090 845.870 ;
        RECT -22.670 844.690 -21.490 845.870 ;
        RECT -24.270 843.090 -23.090 844.270 ;
        RECT -22.670 843.090 -21.490 844.270 ;
        RECT -24.270 664.690 -23.090 665.870 ;
        RECT -22.670 664.690 -21.490 665.870 ;
        RECT -24.270 663.090 -23.090 664.270 ;
        RECT -22.670 663.090 -21.490 664.270 ;
        RECT -24.270 484.690 -23.090 485.870 ;
        RECT -22.670 484.690 -21.490 485.870 ;
        RECT -24.270 483.090 -23.090 484.270 ;
        RECT -22.670 483.090 -21.490 484.270 ;
        RECT -24.270 304.690 -23.090 305.870 ;
        RECT -22.670 304.690 -21.490 305.870 ;
        RECT -24.270 303.090 -23.090 304.270 ;
        RECT -22.670 303.090 -21.490 304.270 ;
        RECT -24.270 124.690 -23.090 125.870 ;
        RECT -22.670 124.690 -21.490 125.870 ;
        RECT -24.270 123.090 -23.090 124.270 ;
        RECT -22.670 123.090 -21.490 124.270 ;
        RECT -24.270 -17.310 -23.090 -16.130 ;
        RECT -22.670 -17.310 -21.490 -16.130 ;
        RECT -24.270 -18.910 -23.090 -17.730 ;
        RECT -22.670 -18.910 -21.490 -17.730 ;
        RECT 117.730 3537.410 118.910 3538.590 ;
        RECT 119.330 3537.410 120.510 3538.590 ;
        RECT 117.730 3535.810 118.910 3536.990 ;
        RECT 119.330 3535.810 120.510 3536.990 ;
        RECT 117.730 3364.690 118.910 3365.870 ;
        RECT 119.330 3364.690 120.510 3365.870 ;
        RECT 117.730 3363.090 118.910 3364.270 ;
        RECT 119.330 3363.090 120.510 3364.270 ;
        RECT 117.730 3184.690 118.910 3185.870 ;
        RECT 119.330 3184.690 120.510 3185.870 ;
        RECT 117.730 3183.090 118.910 3184.270 ;
        RECT 119.330 3183.090 120.510 3184.270 ;
        RECT 117.730 3004.690 118.910 3005.870 ;
        RECT 119.330 3004.690 120.510 3005.870 ;
        RECT 117.730 3003.090 118.910 3004.270 ;
        RECT 119.330 3003.090 120.510 3004.270 ;
        RECT 117.730 2824.690 118.910 2825.870 ;
        RECT 119.330 2824.690 120.510 2825.870 ;
        RECT 117.730 2823.090 118.910 2824.270 ;
        RECT 119.330 2823.090 120.510 2824.270 ;
        RECT 117.730 2644.690 118.910 2645.870 ;
        RECT 119.330 2644.690 120.510 2645.870 ;
        RECT 117.730 2643.090 118.910 2644.270 ;
        RECT 119.330 2643.090 120.510 2644.270 ;
        RECT 117.730 2464.690 118.910 2465.870 ;
        RECT 119.330 2464.690 120.510 2465.870 ;
        RECT 117.730 2463.090 118.910 2464.270 ;
        RECT 119.330 2463.090 120.510 2464.270 ;
        RECT 117.730 2284.690 118.910 2285.870 ;
        RECT 119.330 2284.690 120.510 2285.870 ;
        RECT 117.730 2283.090 118.910 2284.270 ;
        RECT 119.330 2283.090 120.510 2284.270 ;
        RECT 117.730 2104.690 118.910 2105.870 ;
        RECT 119.330 2104.690 120.510 2105.870 ;
        RECT 117.730 2103.090 118.910 2104.270 ;
        RECT 119.330 2103.090 120.510 2104.270 ;
        RECT 117.730 1924.690 118.910 1925.870 ;
        RECT 119.330 1924.690 120.510 1925.870 ;
        RECT 117.730 1923.090 118.910 1924.270 ;
        RECT 119.330 1923.090 120.510 1924.270 ;
        RECT 117.730 1744.690 118.910 1745.870 ;
        RECT 119.330 1744.690 120.510 1745.870 ;
        RECT 117.730 1743.090 118.910 1744.270 ;
        RECT 119.330 1743.090 120.510 1744.270 ;
        RECT 117.730 1564.690 118.910 1565.870 ;
        RECT 119.330 1564.690 120.510 1565.870 ;
        RECT 117.730 1563.090 118.910 1564.270 ;
        RECT 119.330 1563.090 120.510 1564.270 ;
        RECT 117.730 1384.690 118.910 1385.870 ;
        RECT 119.330 1384.690 120.510 1385.870 ;
        RECT 117.730 1383.090 118.910 1384.270 ;
        RECT 119.330 1383.090 120.510 1384.270 ;
        RECT 117.730 1204.690 118.910 1205.870 ;
        RECT 119.330 1204.690 120.510 1205.870 ;
        RECT 117.730 1203.090 118.910 1204.270 ;
        RECT 119.330 1203.090 120.510 1204.270 ;
        RECT 117.730 1024.690 118.910 1025.870 ;
        RECT 119.330 1024.690 120.510 1025.870 ;
        RECT 117.730 1023.090 118.910 1024.270 ;
        RECT 119.330 1023.090 120.510 1024.270 ;
        RECT 297.730 3537.410 298.910 3538.590 ;
        RECT 299.330 3537.410 300.510 3538.590 ;
        RECT 297.730 3535.810 298.910 3536.990 ;
        RECT 299.330 3535.810 300.510 3536.990 ;
        RECT 297.730 3364.690 298.910 3365.870 ;
        RECT 299.330 3364.690 300.510 3365.870 ;
        RECT 297.730 3363.090 298.910 3364.270 ;
        RECT 299.330 3363.090 300.510 3364.270 ;
        RECT 297.730 3184.690 298.910 3185.870 ;
        RECT 299.330 3184.690 300.510 3185.870 ;
        RECT 297.730 3183.090 298.910 3184.270 ;
        RECT 299.330 3183.090 300.510 3184.270 ;
        RECT 297.730 3004.690 298.910 3005.870 ;
        RECT 299.330 3004.690 300.510 3005.870 ;
        RECT 297.730 3003.090 298.910 3004.270 ;
        RECT 299.330 3003.090 300.510 3004.270 ;
        RECT 297.730 2824.690 298.910 2825.870 ;
        RECT 299.330 2824.690 300.510 2825.870 ;
        RECT 297.730 2823.090 298.910 2824.270 ;
        RECT 299.330 2823.090 300.510 2824.270 ;
        RECT 297.730 2644.690 298.910 2645.870 ;
        RECT 299.330 2644.690 300.510 2645.870 ;
        RECT 297.730 2643.090 298.910 2644.270 ;
        RECT 299.330 2643.090 300.510 2644.270 ;
        RECT 297.730 2464.690 298.910 2465.870 ;
        RECT 299.330 2464.690 300.510 2465.870 ;
        RECT 297.730 2463.090 298.910 2464.270 ;
        RECT 299.330 2463.090 300.510 2464.270 ;
        RECT 297.730 2284.690 298.910 2285.870 ;
        RECT 299.330 2284.690 300.510 2285.870 ;
        RECT 297.730 2283.090 298.910 2284.270 ;
        RECT 299.330 2283.090 300.510 2284.270 ;
        RECT 297.730 2104.690 298.910 2105.870 ;
        RECT 299.330 2104.690 300.510 2105.870 ;
        RECT 297.730 2103.090 298.910 2104.270 ;
        RECT 299.330 2103.090 300.510 2104.270 ;
        RECT 297.730 1924.690 298.910 1925.870 ;
        RECT 299.330 1924.690 300.510 1925.870 ;
        RECT 297.730 1923.090 298.910 1924.270 ;
        RECT 299.330 1923.090 300.510 1924.270 ;
        RECT 297.730 1744.690 298.910 1745.870 ;
        RECT 299.330 1744.690 300.510 1745.870 ;
        RECT 297.730 1743.090 298.910 1744.270 ;
        RECT 299.330 1743.090 300.510 1744.270 ;
        RECT 297.730 1564.690 298.910 1565.870 ;
        RECT 299.330 1564.690 300.510 1565.870 ;
        RECT 297.730 1563.090 298.910 1564.270 ;
        RECT 299.330 1563.090 300.510 1564.270 ;
        RECT 297.730 1384.690 298.910 1385.870 ;
        RECT 299.330 1384.690 300.510 1385.870 ;
        RECT 297.730 1383.090 298.910 1384.270 ;
        RECT 299.330 1383.090 300.510 1384.270 ;
        RECT 297.730 1204.690 298.910 1205.870 ;
        RECT 299.330 1204.690 300.510 1205.870 ;
        RECT 297.730 1203.090 298.910 1204.270 ;
        RECT 299.330 1203.090 300.510 1204.270 ;
        RECT 297.730 1024.690 298.910 1025.870 ;
        RECT 299.330 1024.690 300.510 1025.870 ;
        RECT 297.730 1023.090 298.910 1024.270 ;
        RECT 299.330 1023.090 300.510 1024.270 ;
        RECT 477.730 3537.410 478.910 3538.590 ;
        RECT 479.330 3537.410 480.510 3538.590 ;
        RECT 477.730 3535.810 478.910 3536.990 ;
        RECT 479.330 3535.810 480.510 3536.990 ;
        RECT 477.730 3364.690 478.910 3365.870 ;
        RECT 479.330 3364.690 480.510 3365.870 ;
        RECT 477.730 3363.090 478.910 3364.270 ;
        RECT 479.330 3363.090 480.510 3364.270 ;
        RECT 477.730 3184.690 478.910 3185.870 ;
        RECT 479.330 3184.690 480.510 3185.870 ;
        RECT 477.730 3183.090 478.910 3184.270 ;
        RECT 479.330 3183.090 480.510 3184.270 ;
        RECT 477.730 3004.690 478.910 3005.870 ;
        RECT 479.330 3004.690 480.510 3005.870 ;
        RECT 477.730 3003.090 478.910 3004.270 ;
        RECT 479.330 3003.090 480.510 3004.270 ;
        RECT 477.730 2824.690 478.910 2825.870 ;
        RECT 479.330 2824.690 480.510 2825.870 ;
        RECT 477.730 2823.090 478.910 2824.270 ;
        RECT 479.330 2823.090 480.510 2824.270 ;
        RECT 477.730 2644.690 478.910 2645.870 ;
        RECT 479.330 2644.690 480.510 2645.870 ;
        RECT 477.730 2643.090 478.910 2644.270 ;
        RECT 479.330 2643.090 480.510 2644.270 ;
        RECT 477.730 2464.690 478.910 2465.870 ;
        RECT 479.330 2464.690 480.510 2465.870 ;
        RECT 477.730 2463.090 478.910 2464.270 ;
        RECT 479.330 2463.090 480.510 2464.270 ;
        RECT 477.730 2284.690 478.910 2285.870 ;
        RECT 479.330 2284.690 480.510 2285.870 ;
        RECT 477.730 2283.090 478.910 2284.270 ;
        RECT 479.330 2283.090 480.510 2284.270 ;
        RECT 477.730 2104.690 478.910 2105.870 ;
        RECT 479.330 2104.690 480.510 2105.870 ;
        RECT 477.730 2103.090 478.910 2104.270 ;
        RECT 479.330 2103.090 480.510 2104.270 ;
        RECT 477.730 1924.690 478.910 1925.870 ;
        RECT 479.330 1924.690 480.510 1925.870 ;
        RECT 477.730 1923.090 478.910 1924.270 ;
        RECT 479.330 1923.090 480.510 1924.270 ;
        RECT 477.730 1744.690 478.910 1745.870 ;
        RECT 479.330 1744.690 480.510 1745.870 ;
        RECT 477.730 1743.090 478.910 1744.270 ;
        RECT 479.330 1743.090 480.510 1744.270 ;
        RECT 477.730 1564.690 478.910 1565.870 ;
        RECT 479.330 1564.690 480.510 1565.870 ;
        RECT 477.730 1563.090 478.910 1564.270 ;
        RECT 479.330 1563.090 480.510 1564.270 ;
        RECT 477.730 1384.690 478.910 1385.870 ;
        RECT 479.330 1384.690 480.510 1385.870 ;
        RECT 477.730 1383.090 478.910 1384.270 ;
        RECT 479.330 1383.090 480.510 1384.270 ;
        RECT 477.730 1204.690 478.910 1205.870 ;
        RECT 479.330 1204.690 480.510 1205.870 ;
        RECT 477.730 1203.090 478.910 1204.270 ;
        RECT 479.330 1203.090 480.510 1204.270 ;
        RECT 477.730 1024.690 478.910 1025.870 ;
        RECT 479.330 1024.690 480.510 1025.870 ;
        RECT 477.730 1023.090 478.910 1024.270 ;
        RECT 479.330 1023.090 480.510 1024.270 ;
        RECT 657.730 3537.410 658.910 3538.590 ;
        RECT 659.330 3537.410 660.510 3538.590 ;
        RECT 657.730 3535.810 658.910 3536.990 ;
        RECT 659.330 3535.810 660.510 3536.990 ;
        RECT 657.730 3364.690 658.910 3365.870 ;
        RECT 659.330 3364.690 660.510 3365.870 ;
        RECT 657.730 3363.090 658.910 3364.270 ;
        RECT 659.330 3363.090 660.510 3364.270 ;
        RECT 657.730 3184.690 658.910 3185.870 ;
        RECT 659.330 3184.690 660.510 3185.870 ;
        RECT 657.730 3183.090 658.910 3184.270 ;
        RECT 659.330 3183.090 660.510 3184.270 ;
        RECT 657.730 3004.690 658.910 3005.870 ;
        RECT 659.330 3004.690 660.510 3005.870 ;
        RECT 657.730 3003.090 658.910 3004.270 ;
        RECT 659.330 3003.090 660.510 3004.270 ;
        RECT 657.730 2824.690 658.910 2825.870 ;
        RECT 659.330 2824.690 660.510 2825.870 ;
        RECT 657.730 2823.090 658.910 2824.270 ;
        RECT 659.330 2823.090 660.510 2824.270 ;
        RECT 657.730 2644.690 658.910 2645.870 ;
        RECT 659.330 2644.690 660.510 2645.870 ;
        RECT 657.730 2643.090 658.910 2644.270 ;
        RECT 659.330 2643.090 660.510 2644.270 ;
        RECT 657.730 2464.690 658.910 2465.870 ;
        RECT 659.330 2464.690 660.510 2465.870 ;
        RECT 657.730 2463.090 658.910 2464.270 ;
        RECT 659.330 2463.090 660.510 2464.270 ;
        RECT 657.730 2284.690 658.910 2285.870 ;
        RECT 659.330 2284.690 660.510 2285.870 ;
        RECT 657.730 2283.090 658.910 2284.270 ;
        RECT 659.330 2283.090 660.510 2284.270 ;
        RECT 657.730 2104.690 658.910 2105.870 ;
        RECT 659.330 2104.690 660.510 2105.870 ;
        RECT 657.730 2103.090 658.910 2104.270 ;
        RECT 659.330 2103.090 660.510 2104.270 ;
        RECT 657.730 1924.690 658.910 1925.870 ;
        RECT 659.330 1924.690 660.510 1925.870 ;
        RECT 657.730 1923.090 658.910 1924.270 ;
        RECT 659.330 1923.090 660.510 1924.270 ;
        RECT 657.730 1744.690 658.910 1745.870 ;
        RECT 659.330 1744.690 660.510 1745.870 ;
        RECT 657.730 1743.090 658.910 1744.270 ;
        RECT 659.330 1743.090 660.510 1744.270 ;
        RECT 657.730 1564.690 658.910 1565.870 ;
        RECT 659.330 1564.690 660.510 1565.870 ;
        RECT 657.730 1563.090 658.910 1564.270 ;
        RECT 659.330 1563.090 660.510 1564.270 ;
        RECT 657.730 1384.690 658.910 1385.870 ;
        RECT 659.330 1384.690 660.510 1385.870 ;
        RECT 657.730 1383.090 658.910 1384.270 ;
        RECT 659.330 1383.090 660.510 1384.270 ;
        RECT 657.730 1204.690 658.910 1205.870 ;
        RECT 659.330 1204.690 660.510 1205.870 ;
        RECT 657.730 1203.090 658.910 1204.270 ;
        RECT 659.330 1203.090 660.510 1204.270 ;
        RECT 657.730 1024.690 658.910 1025.870 ;
        RECT 659.330 1024.690 660.510 1025.870 ;
        RECT 657.730 1023.090 658.910 1024.270 ;
        RECT 659.330 1023.090 660.510 1024.270 ;
        RECT 837.730 3537.410 838.910 3538.590 ;
        RECT 839.330 3537.410 840.510 3538.590 ;
        RECT 837.730 3535.810 838.910 3536.990 ;
        RECT 839.330 3535.810 840.510 3536.990 ;
        RECT 837.730 3364.690 838.910 3365.870 ;
        RECT 839.330 3364.690 840.510 3365.870 ;
        RECT 837.730 3363.090 838.910 3364.270 ;
        RECT 839.330 3363.090 840.510 3364.270 ;
        RECT 837.730 3184.690 838.910 3185.870 ;
        RECT 839.330 3184.690 840.510 3185.870 ;
        RECT 837.730 3183.090 838.910 3184.270 ;
        RECT 839.330 3183.090 840.510 3184.270 ;
        RECT 837.730 3004.690 838.910 3005.870 ;
        RECT 839.330 3004.690 840.510 3005.870 ;
        RECT 837.730 3003.090 838.910 3004.270 ;
        RECT 839.330 3003.090 840.510 3004.270 ;
        RECT 837.730 2824.690 838.910 2825.870 ;
        RECT 839.330 2824.690 840.510 2825.870 ;
        RECT 837.730 2823.090 838.910 2824.270 ;
        RECT 839.330 2823.090 840.510 2824.270 ;
        RECT 837.730 2644.690 838.910 2645.870 ;
        RECT 839.330 2644.690 840.510 2645.870 ;
        RECT 837.730 2643.090 838.910 2644.270 ;
        RECT 839.330 2643.090 840.510 2644.270 ;
        RECT 837.730 2464.690 838.910 2465.870 ;
        RECT 839.330 2464.690 840.510 2465.870 ;
        RECT 837.730 2463.090 838.910 2464.270 ;
        RECT 839.330 2463.090 840.510 2464.270 ;
        RECT 837.730 2284.690 838.910 2285.870 ;
        RECT 839.330 2284.690 840.510 2285.870 ;
        RECT 837.730 2283.090 838.910 2284.270 ;
        RECT 839.330 2283.090 840.510 2284.270 ;
        RECT 837.730 2104.690 838.910 2105.870 ;
        RECT 839.330 2104.690 840.510 2105.870 ;
        RECT 837.730 2103.090 838.910 2104.270 ;
        RECT 839.330 2103.090 840.510 2104.270 ;
        RECT 837.730 1924.690 838.910 1925.870 ;
        RECT 839.330 1924.690 840.510 1925.870 ;
        RECT 837.730 1923.090 838.910 1924.270 ;
        RECT 839.330 1923.090 840.510 1924.270 ;
        RECT 837.730 1744.690 838.910 1745.870 ;
        RECT 839.330 1744.690 840.510 1745.870 ;
        RECT 837.730 1743.090 838.910 1744.270 ;
        RECT 839.330 1743.090 840.510 1744.270 ;
        RECT 837.730 1564.690 838.910 1565.870 ;
        RECT 839.330 1564.690 840.510 1565.870 ;
        RECT 837.730 1563.090 838.910 1564.270 ;
        RECT 839.330 1563.090 840.510 1564.270 ;
        RECT 837.730 1384.690 838.910 1385.870 ;
        RECT 839.330 1384.690 840.510 1385.870 ;
        RECT 837.730 1383.090 838.910 1384.270 ;
        RECT 839.330 1383.090 840.510 1384.270 ;
        RECT 837.730 1204.690 838.910 1205.870 ;
        RECT 839.330 1204.690 840.510 1205.870 ;
        RECT 837.730 1203.090 838.910 1204.270 ;
        RECT 839.330 1203.090 840.510 1204.270 ;
        RECT 837.730 1024.690 838.910 1025.870 ;
        RECT 839.330 1024.690 840.510 1025.870 ;
        RECT 837.730 1023.090 838.910 1024.270 ;
        RECT 839.330 1023.090 840.510 1024.270 ;
        RECT 1017.730 3537.410 1018.910 3538.590 ;
        RECT 1019.330 3537.410 1020.510 3538.590 ;
        RECT 1017.730 3535.810 1018.910 3536.990 ;
        RECT 1019.330 3535.810 1020.510 3536.990 ;
        RECT 1017.730 3364.690 1018.910 3365.870 ;
        RECT 1019.330 3364.690 1020.510 3365.870 ;
        RECT 1017.730 3363.090 1018.910 3364.270 ;
        RECT 1019.330 3363.090 1020.510 3364.270 ;
        RECT 1017.730 3184.690 1018.910 3185.870 ;
        RECT 1019.330 3184.690 1020.510 3185.870 ;
        RECT 1017.730 3183.090 1018.910 3184.270 ;
        RECT 1019.330 3183.090 1020.510 3184.270 ;
        RECT 1017.730 3004.690 1018.910 3005.870 ;
        RECT 1019.330 3004.690 1020.510 3005.870 ;
        RECT 1017.730 3003.090 1018.910 3004.270 ;
        RECT 1019.330 3003.090 1020.510 3004.270 ;
        RECT 1017.730 2824.690 1018.910 2825.870 ;
        RECT 1019.330 2824.690 1020.510 2825.870 ;
        RECT 1017.730 2823.090 1018.910 2824.270 ;
        RECT 1019.330 2823.090 1020.510 2824.270 ;
        RECT 1017.730 2644.690 1018.910 2645.870 ;
        RECT 1019.330 2644.690 1020.510 2645.870 ;
        RECT 1017.730 2643.090 1018.910 2644.270 ;
        RECT 1019.330 2643.090 1020.510 2644.270 ;
        RECT 1017.730 2464.690 1018.910 2465.870 ;
        RECT 1019.330 2464.690 1020.510 2465.870 ;
        RECT 1017.730 2463.090 1018.910 2464.270 ;
        RECT 1019.330 2463.090 1020.510 2464.270 ;
        RECT 1017.730 2284.690 1018.910 2285.870 ;
        RECT 1019.330 2284.690 1020.510 2285.870 ;
        RECT 1017.730 2283.090 1018.910 2284.270 ;
        RECT 1019.330 2283.090 1020.510 2284.270 ;
        RECT 1017.730 2104.690 1018.910 2105.870 ;
        RECT 1019.330 2104.690 1020.510 2105.870 ;
        RECT 1017.730 2103.090 1018.910 2104.270 ;
        RECT 1019.330 2103.090 1020.510 2104.270 ;
        RECT 1017.730 1924.690 1018.910 1925.870 ;
        RECT 1019.330 1924.690 1020.510 1925.870 ;
        RECT 1017.730 1923.090 1018.910 1924.270 ;
        RECT 1019.330 1923.090 1020.510 1924.270 ;
        RECT 1017.730 1744.690 1018.910 1745.870 ;
        RECT 1019.330 1744.690 1020.510 1745.870 ;
        RECT 1017.730 1743.090 1018.910 1744.270 ;
        RECT 1019.330 1743.090 1020.510 1744.270 ;
        RECT 1017.730 1564.690 1018.910 1565.870 ;
        RECT 1019.330 1564.690 1020.510 1565.870 ;
        RECT 1017.730 1563.090 1018.910 1564.270 ;
        RECT 1019.330 1563.090 1020.510 1564.270 ;
        RECT 1017.730 1384.690 1018.910 1385.870 ;
        RECT 1019.330 1384.690 1020.510 1385.870 ;
        RECT 1017.730 1383.090 1018.910 1384.270 ;
        RECT 1019.330 1383.090 1020.510 1384.270 ;
        RECT 1017.730 1204.690 1018.910 1205.870 ;
        RECT 1019.330 1204.690 1020.510 1205.870 ;
        RECT 1017.730 1203.090 1018.910 1204.270 ;
        RECT 1019.330 1203.090 1020.510 1204.270 ;
        RECT 1017.730 1024.690 1018.910 1025.870 ;
        RECT 1019.330 1024.690 1020.510 1025.870 ;
        RECT 1017.730 1023.090 1018.910 1024.270 ;
        RECT 1019.330 1023.090 1020.510 1024.270 ;
        RECT 1197.730 3537.410 1198.910 3538.590 ;
        RECT 1199.330 3537.410 1200.510 3538.590 ;
        RECT 1197.730 3535.810 1198.910 3536.990 ;
        RECT 1199.330 3535.810 1200.510 3536.990 ;
        RECT 1197.730 3364.690 1198.910 3365.870 ;
        RECT 1199.330 3364.690 1200.510 3365.870 ;
        RECT 1197.730 3363.090 1198.910 3364.270 ;
        RECT 1199.330 3363.090 1200.510 3364.270 ;
        RECT 1197.730 3184.690 1198.910 3185.870 ;
        RECT 1199.330 3184.690 1200.510 3185.870 ;
        RECT 1197.730 3183.090 1198.910 3184.270 ;
        RECT 1199.330 3183.090 1200.510 3184.270 ;
        RECT 1197.730 3004.690 1198.910 3005.870 ;
        RECT 1199.330 3004.690 1200.510 3005.870 ;
        RECT 1197.730 3003.090 1198.910 3004.270 ;
        RECT 1199.330 3003.090 1200.510 3004.270 ;
        RECT 1197.730 2824.690 1198.910 2825.870 ;
        RECT 1199.330 2824.690 1200.510 2825.870 ;
        RECT 1197.730 2823.090 1198.910 2824.270 ;
        RECT 1199.330 2823.090 1200.510 2824.270 ;
        RECT 1197.730 2644.690 1198.910 2645.870 ;
        RECT 1199.330 2644.690 1200.510 2645.870 ;
        RECT 1197.730 2643.090 1198.910 2644.270 ;
        RECT 1199.330 2643.090 1200.510 2644.270 ;
        RECT 1197.730 2464.690 1198.910 2465.870 ;
        RECT 1199.330 2464.690 1200.510 2465.870 ;
        RECT 1197.730 2463.090 1198.910 2464.270 ;
        RECT 1199.330 2463.090 1200.510 2464.270 ;
        RECT 1197.730 2284.690 1198.910 2285.870 ;
        RECT 1199.330 2284.690 1200.510 2285.870 ;
        RECT 1197.730 2283.090 1198.910 2284.270 ;
        RECT 1199.330 2283.090 1200.510 2284.270 ;
        RECT 1197.730 2104.690 1198.910 2105.870 ;
        RECT 1199.330 2104.690 1200.510 2105.870 ;
        RECT 1197.730 2103.090 1198.910 2104.270 ;
        RECT 1199.330 2103.090 1200.510 2104.270 ;
        RECT 1197.730 1924.690 1198.910 1925.870 ;
        RECT 1199.330 1924.690 1200.510 1925.870 ;
        RECT 1197.730 1923.090 1198.910 1924.270 ;
        RECT 1199.330 1923.090 1200.510 1924.270 ;
        RECT 1197.730 1744.690 1198.910 1745.870 ;
        RECT 1199.330 1744.690 1200.510 1745.870 ;
        RECT 1197.730 1743.090 1198.910 1744.270 ;
        RECT 1199.330 1743.090 1200.510 1744.270 ;
        RECT 1197.730 1564.690 1198.910 1565.870 ;
        RECT 1199.330 1564.690 1200.510 1565.870 ;
        RECT 1197.730 1563.090 1198.910 1564.270 ;
        RECT 1199.330 1563.090 1200.510 1564.270 ;
        RECT 1197.730 1384.690 1198.910 1385.870 ;
        RECT 1199.330 1384.690 1200.510 1385.870 ;
        RECT 1197.730 1383.090 1198.910 1384.270 ;
        RECT 1199.330 1383.090 1200.510 1384.270 ;
        RECT 1197.730 1204.690 1198.910 1205.870 ;
        RECT 1199.330 1204.690 1200.510 1205.870 ;
        RECT 1197.730 1203.090 1198.910 1204.270 ;
        RECT 1199.330 1203.090 1200.510 1204.270 ;
        RECT 1197.730 1024.690 1198.910 1025.870 ;
        RECT 1199.330 1024.690 1200.510 1025.870 ;
        RECT 1197.730 1023.090 1198.910 1024.270 ;
        RECT 1199.330 1023.090 1200.510 1024.270 ;
        RECT 117.730 844.690 118.910 845.870 ;
        RECT 119.330 844.690 120.510 845.870 ;
        RECT 117.730 843.090 118.910 844.270 ;
        RECT 119.330 843.090 120.510 844.270 ;
        RECT 117.730 664.690 118.910 665.870 ;
        RECT 119.330 664.690 120.510 665.870 ;
        RECT 117.730 663.090 118.910 664.270 ;
        RECT 119.330 663.090 120.510 664.270 ;
        RECT 117.730 484.690 118.910 485.870 ;
        RECT 119.330 484.690 120.510 485.870 ;
        RECT 117.730 483.090 118.910 484.270 ;
        RECT 119.330 483.090 120.510 484.270 ;
        RECT 1197.730 844.690 1198.910 845.870 ;
        RECT 1199.330 844.690 1200.510 845.870 ;
        RECT 1197.730 843.090 1198.910 844.270 ;
        RECT 1199.330 843.090 1200.510 844.270 ;
        RECT 1197.730 664.690 1198.910 665.870 ;
        RECT 1199.330 664.690 1200.510 665.870 ;
        RECT 1197.730 663.090 1198.910 664.270 ;
        RECT 1199.330 663.090 1200.510 664.270 ;
        RECT 1197.730 484.690 1198.910 485.870 ;
        RECT 1199.330 484.690 1200.510 485.870 ;
        RECT 1197.730 483.090 1198.910 484.270 ;
        RECT 1199.330 483.090 1200.510 484.270 ;
        RECT 117.730 304.690 118.910 305.870 ;
        RECT 119.330 304.690 120.510 305.870 ;
        RECT 117.730 303.090 118.910 304.270 ;
        RECT 119.330 303.090 120.510 304.270 ;
        RECT 117.730 124.690 118.910 125.870 ;
        RECT 119.330 124.690 120.510 125.870 ;
        RECT 117.730 123.090 118.910 124.270 ;
        RECT 119.330 123.090 120.510 124.270 ;
        RECT 117.730 -17.310 118.910 -16.130 ;
        RECT 119.330 -17.310 120.510 -16.130 ;
        RECT 117.730 -18.910 118.910 -17.730 ;
        RECT 119.330 -18.910 120.510 -17.730 ;
        RECT 297.730 304.690 298.910 305.870 ;
        RECT 299.330 304.690 300.510 305.870 ;
        RECT 297.730 303.090 298.910 304.270 ;
        RECT 299.330 303.090 300.510 304.270 ;
        RECT 297.730 124.690 298.910 125.870 ;
        RECT 299.330 124.690 300.510 125.870 ;
        RECT 297.730 123.090 298.910 124.270 ;
        RECT 299.330 123.090 300.510 124.270 ;
        RECT 297.730 -17.310 298.910 -16.130 ;
        RECT 299.330 -17.310 300.510 -16.130 ;
        RECT 297.730 -18.910 298.910 -17.730 ;
        RECT 299.330 -18.910 300.510 -17.730 ;
        RECT 477.730 304.690 478.910 305.870 ;
        RECT 479.330 304.690 480.510 305.870 ;
        RECT 477.730 303.090 478.910 304.270 ;
        RECT 479.330 303.090 480.510 304.270 ;
        RECT 477.730 124.690 478.910 125.870 ;
        RECT 479.330 124.690 480.510 125.870 ;
        RECT 477.730 123.090 478.910 124.270 ;
        RECT 479.330 123.090 480.510 124.270 ;
        RECT 477.730 -17.310 478.910 -16.130 ;
        RECT 479.330 -17.310 480.510 -16.130 ;
        RECT 477.730 -18.910 478.910 -17.730 ;
        RECT 479.330 -18.910 480.510 -17.730 ;
        RECT 657.730 304.690 658.910 305.870 ;
        RECT 659.330 304.690 660.510 305.870 ;
        RECT 657.730 303.090 658.910 304.270 ;
        RECT 659.330 303.090 660.510 304.270 ;
        RECT 657.730 124.690 658.910 125.870 ;
        RECT 659.330 124.690 660.510 125.870 ;
        RECT 657.730 123.090 658.910 124.270 ;
        RECT 659.330 123.090 660.510 124.270 ;
        RECT 657.730 -17.310 658.910 -16.130 ;
        RECT 659.330 -17.310 660.510 -16.130 ;
        RECT 657.730 -18.910 658.910 -17.730 ;
        RECT 659.330 -18.910 660.510 -17.730 ;
        RECT 837.730 304.690 838.910 305.870 ;
        RECT 839.330 304.690 840.510 305.870 ;
        RECT 837.730 303.090 838.910 304.270 ;
        RECT 839.330 303.090 840.510 304.270 ;
        RECT 837.730 124.690 838.910 125.870 ;
        RECT 839.330 124.690 840.510 125.870 ;
        RECT 837.730 123.090 838.910 124.270 ;
        RECT 839.330 123.090 840.510 124.270 ;
        RECT 837.730 -17.310 838.910 -16.130 ;
        RECT 839.330 -17.310 840.510 -16.130 ;
        RECT 837.730 -18.910 838.910 -17.730 ;
        RECT 839.330 -18.910 840.510 -17.730 ;
        RECT 1017.730 304.690 1018.910 305.870 ;
        RECT 1019.330 304.690 1020.510 305.870 ;
        RECT 1017.730 303.090 1018.910 304.270 ;
        RECT 1019.330 303.090 1020.510 304.270 ;
        RECT 1017.730 124.690 1018.910 125.870 ;
        RECT 1019.330 124.690 1020.510 125.870 ;
        RECT 1017.730 123.090 1018.910 124.270 ;
        RECT 1019.330 123.090 1020.510 124.270 ;
        RECT 1017.730 -17.310 1018.910 -16.130 ;
        RECT 1019.330 -17.310 1020.510 -16.130 ;
        RECT 1017.730 -18.910 1018.910 -17.730 ;
        RECT 1019.330 -18.910 1020.510 -17.730 ;
        RECT 1197.730 304.690 1198.910 305.870 ;
        RECT 1199.330 304.690 1200.510 305.870 ;
        RECT 1197.730 303.090 1198.910 304.270 ;
        RECT 1199.330 303.090 1200.510 304.270 ;
        RECT 1197.730 124.690 1198.910 125.870 ;
        RECT 1199.330 124.690 1200.510 125.870 ;
        RECT 1197.730 123.090 1198.910 124.270 ;
        RECT 1199.330 123.090 1200.510 124.270 ;
        RECT 1197.730 -17.310 1198.910 -16.130 ;
        RECT 1199.330 -17.310 1200.510 -16.130 ;
        RECT 1197.730 -18.910 1198.910 -17.730 ;
        RECT 1199.330 -18.910 1200.510 -17.730 ;
        RECT 1377.730 3537.410 1378.910 3538.590 ;
        RECT 1379.330 3537.410 1380.510 3538.590 ;
        RECT 1377.730 3535.810 1378.910 3536.990 ;
        RECT 1379.330 3535.810 1380.510 3536.990 ;
        RECT 1377.730 3364.690 1378.910 3365.870 ;
        RECT 1379.330 3364.690 1380.510 3365.870 ;
        RECT 1377.730 3363.090 1378.910 3364.270 ;
        RECT 1379.330 3363.090 1380.510 3364.270 ;
        RECT 1377.730 3184.690 1378.910 3185.870 ;
        RECT 1379.330 3184.690 1380.510 3185.870 ;
        RECT 1377.730 3183.090 1378.910 3184.270 ;
        RECT 1379.330 3183.090 1380.510 3184.270 ;
        RECT 1377.730 3004.690 1378.910 3005.870 ;
        RECT 1379.330 3004.690 1380.510 3005.870 ;
        RECT 1377.730 3003.090 1378.910 3004.270 ;
        RECT 1379.330 3003.090 1380.510 3004.270 ;
        RECT 1377.730 2824.690 1378.910 2825.870 ;
        RECT 1379.330 2824.690 1380.510 2825.870 ;
        RECT 1377.730 2823.090 1378.910 2824.270 ;
        RECT 1379.330 2823.090 1380.510 2824.270 ;
        RECT 1377.730 2644.690 1378.910 2645.870 ;
        RECT 1379.330 2644.690 1380.510 2645.870 ;
        RECT 1377.730 2643.090 1378.910 2644.270 ;
        RECT 1379.330 2643.090 1380.510 2644.270 ;
        RECT 1377.730 2464.690 1378.910 2465.870 ;
        RECT 1379.330 2464.690 1380.510 2465.870 ;
        RECT 1377.730 2463.090 1378.910 2464.270 ;
        RECT 1379.330 2463.090 1380.510 2464.270 ;
        RECT 1377.730 2284.690 1378.910 2285.870 ;
        RECT 1379.330 2284.690 1380.510 2285.870 ;
        RECT 1377.730 2283.090 1378.910 2284.270 ;
        RECT 1379.330 2283.090 1380.510 2284.270 ;
        RECT 1377.730 2104.690 1378.910 2105.870 ;
        RECT 1379.330 2104.690 1380.510 2105.870 ;
        RECT 1377.730 2103.090 1378.910 2104.270 ;
        RECT 1379.330 2103.090 1380.510 2104.270 ;
        RECT 1377.730 1924.690 1378.910 1925.870 ;
        RECT 1379.330 1924.690 1380.510 1925.870 ;
        RECT 1377.730 1923.090 1378.910 1924.270 ;
        RECT 1379.330 1923.090 1380.510 1924.270 ;
        RECT 1377.730 1744.690 1378.910 1745.870 ;
        RECT 1379.330 1744.690 1380.510 1745.870 ;
        RECT 1377.730 1743.090 1378.910 1744.270 ;
        RECT 1379.330 1743.090 1380.510 1744.270 ;
        RECT 1377.730 1564.690 1378.910 1565.870 ;
        RECT 1379.330 1564.690 1380.510 1565.870 ;
        RECT 1377.730 1563.090 1378.910 1564.270 ;
        RECT 1379.330 1563.090 1380.510 1564.270 ;
        RECT 1377.730 1384.690 1378.910 1385.870 ;
        RECT 1379.330 1384.690 1380.510 1385.870 ;
        RECT 1377.730 1383.090 1378.910 1384.270 ;
        RECT 1379.330 1383.090 1380.510 1384.270 ;
        RECT 1377.730 1204.690 1378.910 1205.870 ;
        RECT 1379.330 1204.690 1380.510 1205.870 ;
        RECT 1377.730 1203.090 1378.910 1204.270 ;
        RECT 1379.330 1203.090 1380.510 1204.270 ;
        RECT 1377.730 1024.690 1378.910 1025.870 ;
        RECT 1379.330 1024.690 1380.510 1025.870 ;
        RECT 1377.730 1023.090 1378.910 1024.270 ;
        RECT 1379.330 1023.090 1380.510 1024.270 ;
        RECT 1377.730 844.690 1378.910 845.870 ;
        RECT 1379.330 844.690 1380.510 845.870 ;
        RECT 1377.730 843.090 1378.910 844.270 ;
        RECT 1379.330 843.090 1380.510 844.270 ;
        RECT 1377.730 664.690 1378.910 665.870 ;
        RECT 1379.330 664.690 1380.510 665.870 ;
        RECT 1377.730 663.090 1378.910 664.270 ;
        RECT 1379.330 663.090 1380.510 664.270 ;
        RECT 1377.730 484.690 1378.910 485.870 ;
        RECT 1379.330 484.690 1380.510 485.870 ;
        RECT 1377.730 483.090 1378.910 484.270 ;
        RECT 1379.330 483.090 1380.510 484.270 ;
        RECT 1377.730 304.690 1378.910 305.870 ;
        RECT 1379.330 304.690 1380.510 305.870 ;
        RECT 1377.730 303.090 1378.910 304.270 ;
        RECT 1379.330 303.090 1380.510 304.270 ;
        RECT 1377.730 124.690 1378.910 125.870 ;
        RECT 1379.330 124.690 1380.510 125.870 ;
        RECT 1377.730 123.090 1378.910 124.270 ;
        RECT 1379.330 123.090 1380.510 124.270 ;
        RECT 1377.730 -17.310 1378.910 -16.130 ;
        RECT 1379.330 -17.310 1380.510 -16.130 ;
        RECT 1377.730 -18.910 1378.910 -17.730 ;
        RECT 1379.330 -18.910 1380.510 -17.730 ;
        RECT 1557.730 3537.410 1558.910 3538.590 ;
        RECT 1559.330 3537.410 1560.510 3538.590 ;
        RECT 1557.730 3535.810 1558.910 3536.990 ;
        RECT 1559.330 3535.810 1560.510 3536.990 ;
        RECT 1557.730 3364.690 1558.910 3365.870 ;
        RECT 1559.330 3364.690 1560.510 3365.870 ;
        RECT 1557.730 3363.090 1558.910 3364.270 ;
        RECT 1559.330 3363.090 1560.510 3364.270 ;
        RECT 1557.730 3184.690 1558.910 3185.870 ;
        RECT 1559.330 3184.690 1560.510 3185.870 ;
        RECT 1557.730 3183.090 1558.910 3184.270 ;
        RECT 1559.330 3183.090 1560.510 3184.270 ;
        RECT 1557.730 3004.690 1558.910 3005.870 ;
        RECT 1559.330 3004.690 1560.510 3005.870 ;
        RECT 1557.730 3003.090 1558.910 3004.270 ;
        RECT 1559.330 3003.090 1560.510 3004.270 ;
        RECT 1557.730 2824.690 1558.910 2825.870 ;
        RECT 1559.330 2824.690 1560.510 2825.870 ;
        RECT 1557.730 2823.090 1558.910 2824.270 ;
        RECT 1559.330 2823.090 1560.510 2824.270 ;
        RECT 1557.730 2644.690 1558.910 2645.870 ;
        RECT 1559.330 2644.690 1560.510 2645.870 ;
        RECT 1557.730 2643.090 1558.910 2644.270 ;
        RECT 1559.330 2643.090 1560.510 2644.270 ;
        RECT 1557.730 2464.690 1558.910 2465.870 ;
        RECT 1559.330 2464.690 1560.510 2465.870 ;
        RECT 1557.730 2463.090 1558.910 2464.270 ;
        RECT 1559.330 2463.090 1560.510 2464.270 ;
        RECT 1557.730 2284.690 1558.910 2285.870 ;
        RECT 1559.330 2284.690 1560.510 2285.870 ;
        RECT 1557.730 2283.090 1558.910 2284.270 ;
        RECT 1559.330 2283.090 1560.510 2284.270 ;
        RECT 1557.730 2104.690 1558.910 2105.870 ;
        RECT 1559.330 2104.690 1560.510 2105.870 ;
        RECT 1557.730 2103.090 1558.910 2104.270 ;
        RECT 1559.330 2103.090 1560.510 2104.270 ;
        RECT 1557.730 1924.690 1558.910 1925.870 ;
        RECT 1559.330 1924.690 1560.510 1925.870 ;
        RECT 1557.730 1923.090 1558.910 1924.270 ;
        RECT 1559.330 1923.090 1560.510 1924.270 ;
        RECT 1557.730 1744.690 1558.910 1745.870 ;
        RECT 1559.330 1744.690 1560.510 1745.870 ;
        RECT 1557.730 1743.090 1558.910 1744.270 ;
        RECT 1559.330 1743.090 1560.510 1744.270 ;
        RECT 1557.730 1564.690 1558.910 1565.870 ;
        RECT 1559.330 1564.690 1560.510 1565.870 ;
        RECT 1557.730 1563.090 1558.910 1564.270 ;
        RECT 1559.330 1563.090 1560.510 1564.270 ;
        RECT 1557.730 1384.690 1558.910 1385.870 ;
        RECT 1559.330 1384.690 1560.510 1385.870 ;
        RECT 1557.730 1383.090 1558.910 1384.270 ;
        RECT 1559.330 1383.090 1560.510 1384.270 ;
        RECT 1557.730 1204.690 1558.910 1205.870 ;
        RECT 1559.330 1204.690 1560.510 1205.870 ;
        RECT 1557.730 1203.090 1558.910 1204.270 ;
        RECT 1559.330 1203.090 1560.510 1204.270 ;
        RECT 1557.730 1024.690 1558.910 1025.870 ;
        RECT 1559.330 1024.690 1560.510 1025.870 ;
        RECT 1557.730 1023.090 1558.910 1024.270 ;
        RECT 1559.330 1023.090 1560.510 1024.270 ;
        RECT 1557.730 844.690 1558.910 845.870 ;
        RECT 1559.330 844.690 1560.510 845.870 ;
        RECT 1557.730 843.090 1558.910 844.270 ;
        RECT 1559.330 843.090 1560.510 844.270 ;
        RECT 1557.730 664.690 1558.910 665.870 ;
        RECT 1559.330 664.690 1560.510 665.870 ;
        RECT 1557.730 663.090 1558.910 664.270 ;
        RECT 1559.330 663.090 1560.510 664.270 ;
        RECT 1557.730 484.690 1558.910 485.870 ;
        RECT 1559.330 484.690 1560.510 485.870 ;
        RECT 1557.730 483.090 1558.910 484.270 ;
        RECT 1559.330 483.090 1560.510 484.270 ;
        RECT 1557.730 304.690 1558.910 305.870 ;
        RECT 1559.330 304.690 1560.510 305.870 ;
        RECT 1557.730 303.090 1558.910 304.270 ;
        RECT 1559.330 303.090 1560.510 304.270 ;
        RECT 1557.730 124.690 1558.910 125.870 ;
        RECT 1559.330 124.690 1560.510 125.870 ;
        RECT 1557.730 123.090 1558.910 124.270 ;
        RECT 1559.330 123.090 1560.510 124.270 ;
        RECT 1557.730 -17.310 1558.910 -16.130 ;
        RECT 1559.330 -17.310 1560.510 -16.130 ;
        RECT 1557.730 -18.910 1558.910 -17.730 ;
        RECT 1559.330 -18.910 1560.510 -17.730 ;
        RECT 1737.730 3537.410 1738.910 3538.590 ;
        RECT 1739.330 3537.410 1740.510 3538.590 ;
        RECT 1737.730 3535.810 1738.910 3536.990 ;
        RECT 1739.330 3535.810 1740.510 3536.990 ;
        RECT 1737.730 3364.690 1738.910 3365.870 ;
        RECT 1739.330 3364.690 1740.510 3365.870 ;
        RECT 1737.730 3363.090 1738.910 3364.270 ;
        RECT 1739.330 3363.090 1740.510 3364.270 ;
        RECT 1737.730 3184.690 1738.910 3185.870 ;
        RECT 1739.330 3184.690 1740.510 3185.870 ;
        RECT 1737.730 3183.090 1738.910 3184.270 ;
        RECT 1739.330 3183.090 1740.510 3184.270 ;
        RECT 1737.730 3004.690 1738.910 3005.870 ;
        RECT 1739.330 3004.690 1740.510 3005.870 ;
        RECT 1737.730 3003.090 1738.910 3004.270 ;
        RECT 1739.330 3003.090 1740.510 3004.270 ;
        RECT 1737.730 2824.690 1738.910 2825.870 ;
        RECT 1739.330 2824.690 1740.510 2825.870 ;
        RECT 1737.730 2823.090 1738.910 2824.270 ;
        RECT 1739.330 2823.090 1740.510 2824.270 ;
        RECT 1737.730 2644.690 1738.910 2645.870 ;
        RECT 1739.330 2644.690 1740.510 2645.870 ;
        RECT 1737.730 2643.090 1738.910 2644.270 ;
        RECT 1739.330 2643.090 1740.510 2644.270 ;
        RECT 1737.730 2464.690 1738.910 2465.870 ;
        RECT 1739.330 2464.690 1740.510 2465.870 ;
        RECT 1737.730 2463.090 1738.910 2464.270 ;
        RECT 1739.330 2463.090 1740.510 2464.270 ;
        RECT 1737.730 2284.690 1738.910 2285.870 ;
        RECT 1739.330 2284.690 1740.510 2285.870 ;
        RECT 1737.730 2283.090 1738.910 2284.270 ;
        RECT 1739.330 2283.090 1740.510 2284.270 ;
        RECT 1737.730 2104.690 1738.910 2105.870 ;
        RECT 1739.330 2104.690 1740.510 2105.870 ;
        RECT 1737.730 2103.090 1738.910 2104.270 ;
        RECT 1739.330 2103.090 1740.510 2104.270 ;
        RECT 1737.730 1924.690 1738.910 1925.870 ;
        RECT 1739.330 1924.690 1740.510 1925.870 ;
        RECT 1737.730 1923.090 1738.910 1924.270 ;
        RECT 1739.330 1923.090 1740.510 1924.270 ;
        RECT 1737.730 1744.690 1738.910 1745.870 ;
        RECT 1739.330 1744.690 1740.510 1745.870 ;
        RECT 1737.730 1743.090 1738.910 1744.270 ;
        RECT 1739.330 1743.090 1740.510 1744.270 ;
        RECT 1737.730 1564.690 1738.910 1565.870 ;
        RECT 1739.330 1564.690 1740.510 1565.870 ;
        RECT 1737.730 1563.090 1738.910 1564.270 ;
        RECT 1739.330 1563.090 1740.510 1564.270 ;
        RECT 1737.730 1384.690 1738.910 1385.870 ;
        RECT 1739.330 1384.690 1740.510 1385.870 ;
        RECT 1737.730 1383.090 1738.910 1384.270 ;
        RECT 1739.330 1383.090 1740.510 1384.270 ;
        RECT 1737.730 1204.690 1738.910 1205.870 ;
        RECT 1739.330 1204.690 1740.510 1205.870 ;
        RECT 1737.730 1203.090 1738.910 1204.270 ;
        RECT 1739.330 1203.090 1740.510 1204.270 ;
        RECT 1737.730 1024.690 1738.910 1025.870 ;
        RECT 1739.330 1024.690 1740.510 1025.870 ;
        RECT 1737.730 1023.090 1738.910 1024.270 ;
        RECT 1739.330 1023.090 1740.510 1024.270 ;
        RECT 1737.730 844.690 1738.910 845.870 ;
        RECT 1739.330 844.690 1740.510 845.870 ;
        RECT 1737.730 843.090 1738.910 844.270 ;
        RECT 1739.330 843.090 1740.510 844.270 ;
        RECT 1737.730 664.690 1738.910 665.870 ;
        RECT 1739.330 664.690 1740.510 665.870 ;
        RECT 1737.730 663.090 1738.910 664.270 ;
        RECT 1739.330 663.090 1740.510 664.270 ;
        RECT 1737.730 484.690 1738.910 485.870 ;
        RECT 1739.330 484.690 1740.510 485.870 ;
        RECT 1737.730 483.090 1738.910 484.270 ;
        RECT 1739.330 483.090 1740.510 484.270 ;
        RECT 1737.730 304.690 1738.910 305.870 ;
        RECT 1739.330 304.690 1740.510 305.870 ;
        RECT 1737.730 303.090 1738.910 304.270 ;
        RECT 1739.330 303.090 1740.510 304.270 ;
        RECT 1737.730 124.690 1738.910 125.870 ;
        RECT 1739.330 124.690 1740.510 125.870 ;
        RECT 1737.730 123.090 1738.910 124.270 ;
        RECT 1739.330 123.090 1740.510 124.270 ;
        RECT 1737.730 -17.310 1738.910 -16.130 ;
        RECT 1739.330 -17.310 1740.510 -16.130 ;
        RECT 1737.730 -18.910 1738.910 -17.730 ;
        RECT 1739.330 -18.910 1740.510 -17.730 ;
        RECT 1917.730 3537.410 1918.910 3538.590 ;
        RECT 1919.330 3537.410 1920.510 3538.590 ;
        RECT 1917.730 3535.810 1918.910 3536.990 ;
        RECT 1919.330 3535.810 1920.510 3536.990 ;
        RECT 1917.730 3364.690 1918.910 3365.870 ;
        RECT 1919.330 3364.690 1920.510 3365.870 ;
        RECT 1917.730 3363.090 1918.910 3364.270 ;
        RECT 1919.330 3363.090 1920.510 3364.270 ;
        RECT 1917.730 3184.690 1918.910 3185.870 ;
        RECT 1919.330 3184.690 1920.510 3185.870 ;
        RECT 1917.730 3183.090 1918.910 3184.270 ;
        RECT 1919.330 3183.090 1920.510 3184.270 ;
        RECT 1917.730 3004.690 1918.910 3005.870 ;
        RECT 1919.330 3004.690 1920.510 3005.870 ;
        RECT 1917.730 3003.090 1918.910 3004.270 ;
        RECT 1919.330 3003.090 1920.510 3004.270 ;
        RECT 1917.730 2824.690 1918.910 2825.870 ;
        RECT 1919.330 2824.690 1920.510 2825.870 ;
        RECT 1917.730 2823.090 1918.910 2824.270 ;
        RECT 1919.330 2823.090 1920.510 2824.270 ;
        RECT 1917.730 2644.690 1918.910 2645.870 ;
        RECT 1919.330 2644.690 1920.510 2645.870 ;
        RECT 1917.730 2643.090 1918.910 2644.270 ;
        RECT 1919.330 2643.090 1920.510 2644.270 ;
        RECT 1917.730 2464.690 1918.910 2465.870 ;
        RECT 1919.330 2464.690 1920.510 2465.870 ;
        RECT 1917.730 2463.090 1918.910 2464.270 ;
        RECT 1919.330 2463.090 1920.510 2464.270 ;
        RECT 1917.730 2284.690 1918.910 2285.870 ;
        RECT 1919.330 2284.690 1920.510 2285.870 ;
        RECT 1917.730 2283.090 1918.910 2284.270 ;
        RECT 1919.330 2283.090 1920.510 2284.270 ;
        RECT 1917.730 2104.690 1918.910 2105.870 ;
        RECT 1919.330 2104.690 1920.510 2105.870 ;
        RECT 1917.730 2103.090 1918.910 2104.270 ;
        RECT 1919.330 2103.090 1920.510 2104.270 ;
        RECT 1917.730 1924.690 1918.910 1925.870 ;
        RECT 1919.330 1924.690 1920.510 1925.870 ;
        RECT 1917.730 1923.090 1918.910 1924.270 ;
        RECT 1919.330 1923.090 1920.510 1924.270 ;
        RECT 1917.730 1744.690 1918.910 1745.870 ;
        RECT 1919.330 1744.690 1920.510 1745.870 ;
        RECT 1917.730 1743.090 1918.910 1744.270 ;
        RECT 1919.330 1743.090 1920.510 1744.270 ;
        RECT 1917.730 1564.690 1918.910 1565.870 ;
        RECT 1919.330 1564.690 1920.510 1565.870 ;
        RECT 1917.730 1563.090 1918.910 1564.270 ;
        RECT 1919.330 1563.090 1920.510 1564.270 ;
        RECT 1917.730 1384.690 1918.910 1385.870 ;
        RECT 1919.330 1384.690 1920.510 1385.870 ;
        RECT 1917.730 1383.090 1918.910 1384.270 ;
        RECT 1919.330 1383.090 1920.510 1384.270 ;
        RECT 1917.730 1204.690 1918.910 1205.870 ;
        RECT 1919.330 1204.690 1920.510 1205.870 ;
        RECT 1917.730 1203.090 1918.910 1204.270 ;
        RECT 1919.330 1203.090 1920.510 1204.270 ;
        RECT 1917.730 1024.690 1918.910 1025.870 ;
        RECT 1919.330 1024.690 1920.510 1025.870 ;
        RECT 1917.730 1023.090 1918.910 1024.270 ;
        RECT 1919.330 1023.090 1920.510 1024.270 ;
        RECT 1917.730 844.690 1918.910 845.870 ;
        RECT 1919.330 844.690 1920.510 845.870 ;
        RECT 1917.730 843.090 1918.910 844.270 ;
        RECT 1919.330 843.090 1920.510 844.270 ;
        RECT 1917.730 664.690 1918.910 665.870 ;
        RECT 1919.330 664.690 1920.510 665.870 ;
        RECT 1917.730 663.090 1918.910 664.270 ;
        RECT 1919.330 663.090 1920.510 664.270 ;
        RECT 1917.730 484.690 1918.910 485.870 ;
        RECT 1919.330 484.690 1920.510 485.870 ;
        RECT 1917.730 483.090 1918.910 484.270 ;
        RECT 1919.330 483.090 1920.510 484.270 ;
        RECT 1917.730 304.690 1918.910 305.870 ;
        RECT 1919.330 304.690 1920.510 305.870 ;
        RECT 1917.730 303.090 1918.910 304.270 ;
        RECT 1919.330 303.090 1920.510 304.270 ;
        RECT 1917.730 124.690 1918.910 125.870 ;
        RECT 1919.330 124.690 1920.510 125.870 ;
        RECT 1917.730 123.090 1918.910 124.270 ;
        RECT 1919.330 123.090 1920.510 124.270 ;
        RECT 1917.730 -17.310 1918.910 -16.130 ;
        RECT 1919.330 -17.310 1920.510 -16.130 ;
        RECT 1917.730 -18.910 1918.910 -17.730 ;
        RECT 1919.330 -18.910 1920.510 -17.730 ;
        RECT 2097.730 3537.410 2098.910 3538.590 ;
        RECT 2099.330 3537.410 2100.510 3538.590 ;
        RECT 2097.730 3535.810 2098.910 3536.990 ;
        RECT 2099.330 3535.810 2100.510 3536.990 ;
        RECT 2097.730 3364.690 2098.910 3365.870 ;
        RECT 2099.330 3364.690 2100.510 3365.870 ;
        RECT 2097.730 3363.090 2098.910 3364.270 ;
        RECT 2099.330 3363.090 2100.510 3364.270 ;
        RECT 2097.730 3184.690 2098.910 3185.870 ;
        RECT 2099.330 3184.690 2100.510 3185.870 ;
        RECT 2097.730 3183.090 2098.910 3184.270 ;
        RECT 2099.330 3183.090 2100.510 3184.270 ;
        RECT 2097.730 3004.690 2098.910 3005.870 ;
        RECT 2099.330 3004.690 2100.510 3005.870 ;
        RECT 2097.730 3003.090 2098.910 3004.270 ;
        RECT 2099.330 3003.090 2100.510 3004.270 ;
        RECT 2097.730 2824.690 2098.910 2825.870 ;
        RECT 2099.330 2824.690 2100.510 2825.870 ;
        RECT 2097.730 2823.090 2098.910 2824.270 ;
        RECT 2099.330 2823.090 2100.510 2824.270 ;
        RECT 2097.730 2644.690 2098.910 2645.870 ;
        RECT 2099.330 2644.690 2100.510 2645.870 ;
        RECT 2097.730 2643.090 2098.910 2644.270 ;
        RECT 2099.330 2643.090 2100.510 2644.270 ;
        RECT 2097.730 2464.690 2098.910 2465.870 ;
        RECT 2099.330 2464.690 2100.510 2465.870 ;
        RECT 2097.730 2463.090 2098.910 2464.270 ;
        RECT 2099.330 2463.090 2100.510 2464.270 ;
        RECT 2097.730 2284.690 2098.910 2285.870 ;
        RECT 2099.330 2284.690 2100.510 2285.870 ;
        RECT 2097.730 2283.090 2098.910 2284.270 ;
        RECT 2099.330 2283.090 2100.510 2284.270 ;
        RECT 2097.730 2104.690 2098.910 2105.870 ;
        RECT 2099.330 2104.690 2100.510 2105.870 ;
        RECT 2097.730 2103.090 2098.910 2104.270 ;
        RECT 2099.330 2103.090 2100.510 2104.270 ;
        RECT 2097.730 1924.690 2098.910 1925.870 ;
        RECT 2099.330 1924.690 2100.510 1925.870 ;
        RECT 2097.730 1923.090 2098.910 1924.270 ;
        RECT 2099.330 1923.090 2100.510 1924.270 ;
        RECT 2097.730 1744.690 2098.910 1745.870 ;
        RECT 2099.330 1744.690 2100.510 1745.870 ;
        RECT 2097.730 1743.090 2098.910 1744.270 ;
        RECT 2099.330 1743.090 2100.510 1744.270 ;
        RECT 2097.730 1564.690 2098.910 1565.870 ;
        RECT 2099.330 1564.690 2100.510 1565.870 ;
        RECT 2097.730 1563.090 2098.910 1564.270 ;
        RECT 2099.330 1563.090 2100.510 1564.270 ;
        RECT 2097.730 1384.690 2098.910 1385.870 ;
        RECT 2099.330 1384.690 2100.510 1385.870 ;
        RECT 2097.730 1383.090 2098.910 1384.270 ;
        RECT 2099.330 1383.090 2100.510 1384.270 ;
        RECT 2097.730 1204.690 2098.910 1205.870 ;
        RECT 2099.330 1204.690 2100.510 1205.870 ;
        RECT 2097.730 1203.090 2098.910 1204.270 ;
        RECT 2099.330 1203.090 2100.510 1204.270 ;
        RECT 2097.730 1024.690 2098.910 1025.870 ;
        RECT 2099.330 1024.690 2100.510 1025.870 ;
        RECT 2097.730 1023.090 2098.910 1024.270 ;
        RECT 2099.330 1023.090 2100.510 1024.270 ;
        RECT 2097.730 844.690 2098.910 845.870 ;
        RECT 2099.330 844.690 2100.510 845.870 ;
        RECT 2097.730 843.090 2098.910 844.270 ;
        RECT 2099.330 843.090 2100.510 844.270 ;
        RECT 2097.730 664.690 2098.910 665.870 ;
        RECT 2099.330 664.690 2100.510 665.870 ;
        RECT 2097.730 663.090 2098.910 664.270 ;
        RECT 2099.330 663.090 2100.510 664.270 ;
        RECT 2097.730 484.690 2098.910 485.870 ;
        RECT 2099.330 484.690 2100.510 485.870 ;
        RECT 2097.730 483.090 2098.910 484.270 ;
        RECT 2099.330 483.090 2100.510 484.270 ;
        RECT 2097.730 304.690 2098.910 305.870 ;
        RECT 2099.330 304.690 2100.510 305.870 ;
        RECT 2097.730 303.090 2098.910 304.270 ;
        RECT 2099.330 303.090 2100.510 304.270 ;
        RECT 2097.730 124.690 2098.910 125.870 ;
        RECT 2099.330 124.690 2100.510 125.870 ;
        RECT 2097.730 123.090 2098.910 124.270 ;
        RECT 2099.330 123.090 2100.510 124.270 ;
        RECT 2097.730 -17.310 2098.910 -16.130 ;
        RECT 2099.330 -17.310 2100.510 -16.130 ;
        RECT 2097.730 -18.910 2098.910 -17.730 ;
        RECT 2099.330 -18.910 2100.510 -17.730 ;
        RECT 2277.730 3537.410 2278.910 3538.590 ;
        RECT 2279.330 3537.410 2280.510 3538.590 ;
        RECT 2277.730 3535.810 2278.910 3536.990 ;
        RECT 2279.330 3535.810 2280.510 3536.990 ;
        RECT 2277.730 3364.690 2278.910 3365.870 ;
        RECT 2279.330 3364.690 2280.510 3365.870 ;
        RECT 2277.730 3363.090 2278.910 3364.270 ;
        RECT 2279.330 3363.090 2280.510 3364.270 ;
        RECT 2277.730 3184.690 2278.910 3185.870 ;
        RECT 2279.330 3184.690 2280.510 3185.870 ;
        RECT 2277.730 3183.090 2278.910 3184.270 ;
        RECT 2279.330 3183.090 2280.510 3184.270 ;
        RECT 2277.730 3004.690 2278.910 3005.870 ;
        RECT 2279.330 3004.690 2280.510 3005.870 ;
        RECT 2277.730 3003.090 2278.910 3004.270 ;
        RECT 2279.330 3003.090 2280.510 3004.270 ;
        RECT 2277.730 2824.690 2278.910 2825.870 ;
        RECT 2279.330 2824.690 2280.510 2825.870 ;
        RECT 2277.730 2823.090 2278.910 2824.270 ;
        RECT 2279.330 2823.090 2280.510 2824.270 ;
        RECT 2277.730 2644.690 2278.910 2645.870 ;
        RECT 2279.330 2644.690 2280.510 2645.870 ;
        RECT 2277.730 2643.090 2278.910 2644.270 ;
        RECT 2279.330 2643.090 2280.510 2644.270 ;
        RECT 2277.730 2464.690 2278.910 2465.870 ;
        RECT 2279.330 2464.690 2280.510 2465.870 ;
        RECT 2277.730 2463.090 2278.910 2464.270 ;
        RECT 2279.330 2463.090 2280.510 2464.270 ;
        RECT 2277.730 2284.690 2278.910 2285.870 ;
        RECT 2279.330 2284.690 2280.510 2285.870 ;
        RECT 2277.730 2283.090 2278.910 2284.270 ;
        RECT 2279.330 2283.090 2280.510 2284.270 ;
        RECT 2277.730 2104.690 2278.910 2105.870 ;
        RECT 2279.330 2104.690 2280.510 2105.870 ;
        RECT 2277.730 2103.090 2278.910 2104.270 ;
        RECT 2279.330 2103.090 2280.510 2104.270 ;
        RECT 2277.730 1924.690 2278.910 1925.870 ;
        RECT 2279.330 1924.690 2280.510 1925.870 ;
        RECT 2277.730 1923.090 2278.910 1924.270 ;
        RECT 2279.330 1923.090 2280.510 1924.270 ;
        RECT 2277.730 1744.690 2278.910 1745.870 ;
        RECT 2279.330 1744.690 2280.510 1745.870 ;
        RECT 2277.730 1743.090 2278.910 1744.270 ;
        RECT 2279.330 1743.090 2280.510 1744.270 ;
        RECT 2277.730 1564.690 2278.910 1565.870 ;
        RECT 2279.330 1564.690 2280.510 1565.870 ;
        RECT 2277.730 1563.090 2278.910 1564.270 ;
        RECT 2279.330 1563.090 2280.510 1564.270 ;
        RECT 2277.730 1384.690 2278.910 1385.870 ;
        RECT 2279.330 1384.690 2280.510 1385.870 ;
        RECT 2277.730 1383.090 2278.910 1384.270 ;
        RECT 2279.330 1383.090 2280.510 1384.270 ;
        RECT 2277.730 1204.690 2278.910 1205.870 ;
        RECT 2279.330 1204.690 2280.510 1205.870 ;
        RECT 2277.730 1203.090 2278.910 1204.270 ;
        RECT 2279.330 1203.090 2280.510 1204.270 ;
        RECT 2277.730 1024.690 2278.910 1025.870 ;
        RECT 2279.330 1024.690 2280.510 1025.870 ;
        RECT 2277.730 1023.090 2278.910 1024.270 ;
        RECT 2279.330 1023.090 2280.510 1024.270 ;
        RECT 2277.730 844.690 2278.910 845.870 ;
        RECT 2279.330 844.690 2280.510 845.870 ;
        RECT 2277.730 843.090 2278.910 844.270 ;
        RECT 2279.330 843.090 2280.510 844.270 ;
        RECT 2277.730 664.690 2278.910 665.870 ;
        RECT 2279.330 664.690 2280.510 665.870 ;
        RECT 2277.730 663.090 2278.910 664.270 ;
        RECT 2279.330 663.090 2280.510 664.270 ;
        RECT 2277.730 484.690 2278.910 485.870 ;
        RECT 2279.330 484.690 2280.510 485.870 ;
        RECT 2277.730 483.090 2278.910 484.270 ;
        RECT 2279.330 483.090 2280.510 484.270 ;
        RECT 2277.730 304.690 2278.910 305.870 ;
        RECT 2279.330 304.690 2280.510 305.870 ;
        RECT 2277.730 303.090 2278.910 304.270 ;
        RECT 2279.330 303.090 2280.510 304.270 ;
        RECT 2277.730 124.690 2278.910 125.870 ;
        RECT 2279.330 124.690 2280.510 125.870 ;
        RECT 2277.730 123.090 2278.910 124.270 ;
        RECT 2279.330 123.090 2280.510 124.270 ;
        RECT 2277.730 -17.310 2278.910 -16.130 ;
        RECT 2279.330 -17.310 2280.510 -16.130 ;
        RECT 2277.730 -18.910 2278.910 -17.730 ;
        RECT 2279.330 -18.910 2280.510 -17.730 ;
        RECT 2457.730 3537.410 2458.910 3538.590 ;
        RECT 2459.330 3537.410 2460.510 3538.590 ;
        RECT 2457.730 3535.810 2458.910 3536.990 ;
        RECT 2459.330 3535.810 2460.510 3536.990 ;
        RECT 2457.730 3364.690 2458.910 3365.870 ;
        RECT 2459.330 3364.690 2460.510 3365.870 ;
        RECT 2457.730 3363.090 2458.910 3364.270 ;
        RECT 2459.330 3363.090 2460.510 3364.270 ;
        RECT 2457.730 3184.690 2458.910 3185.870 ;
        RECT 2459.330 3184.690 2460.510 3185.870 ;
        RECT 2457.730 3183.090 2458.910 3184.270 ;
        RECT 2459.330 3183.090 2460.510 3184.270 ;
        RECT 2457.730 3004.690 2458.910 3005.870 ;
        RECT 2459.330 3004.690 2460.510 3005.870 ;
        RECT 2457.730 3003.090 2458.910 3004.270 ;
        RECT 2459.330 3003.090 2460.510 3004.270 ;
        RECT 2457.730 2824.690 2458.910 2825.870 ;
        RECT 2459.330 2824.690 2460.510 2825.870 ;
        RECT 2457.730 2823.090 2458.910 2824.270 ;
        RECT 2459.330 2823.090 2460.510 2824.270 ;
        RECT 2457.730 2644.690 2458.910 2645.870 ;
        RECT 2459.330 2644.690 2460.510 2645.870 ;
        RECT 2457.730 2643.090 2458.910 2644.270 ;
        RECT 2459.330 2643.090 2460.510 2644.270 ;
        RECT 2457.730 2464.690 2458.910 2465.870 ;
        RECT 2459.330 2464.690 2460.510 2465.870 ;
        RECT 2457.730 2463.090 2458.910 2464.270 ;
        RECT 2459.330 2463.090 2460.510 2464.270 ;
        RECT 2457.730 2284.690 2458.910 2285.870 ;
        RECT 2459.330 2284.690 2460.510 2285.870 ;
        RECT 2457.730 2283.090 2458.910 2284.270 ;
        RECT 2459.330 2283.090 2460.510 2284.270 ;
        RECT 2457.730 2104.690 2458.910 2105.870 ;
        RECT 2459.330 2104.690 2460.510 2105.870 ;
        RECT 2457.730 2103.090 2458.910 2104.270 ;
        RECT 2459.330 2103.090 2460.510 2104.270 ;
        RECT 2457.730 1924.690 2458.910 1925.870 ;
        RECT 2459.330 1924.690 2460.510 1925.870 ;
        RECT 2457.730 1923.090 2458.910 1924.270 ;
        RECT 2459.330 1923.090 2460.510 1924.270 ;
        RECT 2457.730 1744.690 2458.910 1745.870 ;
        RECT 2459.330 1744.690 2460.510 1745.870 ;
        RECT 2457.730 1743.090 2458.910 1744.270 ;
        RECT 2459.330 1743.090 2460.510 1744.270 ;
        RECT 2457.730 1564.690 2458.910 1565.870 ;
        RECT 2459.330 1564.690 2460.510 1565.870 ;
        RECT 2457.730 1563.090 2458.910 1564.270 ;
        RECT 2459.330 1563.090 2460.510 1564.270 ;
        RECT 2457.730 1384.690 2458.910 1385.870 ;
        RECT 2459.330 1384.690 2460.510 1385.870 ;
        RECT 2457.730 1383.090 2458.910 1384.270 ;
        RECT 2459.330 1383.090 2460.510 1384.270 ;
        RECT 2457.730 1204.690 2458.910 1205.870 ;
        RECT 2459.330 1204.690 2460.510 1205.870 ;
        RECT 2457.730 1203.090 2458.910 1204.270 ;
        RECT 2459.330 1203.090 2460.510 1204.270 ;
        RECT 2457.730 1024.690 2458.910 1025.870 ;
        RECT 2459.330 1024.690 2460.510 1025.870 ;
        RECT 2457.730 1023.090 2458.910 1024.270 ;
        RECT 2459.330 1023.090 2460.510 1024.270 ;
        RECT 2457.730 844.690 2458.910 845.870 ;
        RECT 2459.330 844.690 2460.510 845.870 ;
        RECT 2457.730 843.090 2458.910 844.270 ;
        RECT 2459.330 843.090 2460.510 844.270 ;
        RECT 2457.730 664.690 2458.910 665.870 ;
        RECT 2459.330 664.690 2460.510 665.870 ;
        RECT 2457.730 663.090 2458.910 664.270 ;
        RECT 2459.330 663.090 2460.510 664.270 ;
        RECT 2457.730 484.690 2458.910 485.870 ;
        RECT 2459.330 484.690 2460.510 485.870 ;
        RECT 2457.730 483.090 2458.910 484.270 ;
        RECT 2459.330 483.090 2460.510 484.270 ;
        RECT 2457.730 304.690 2458.910 305.870 ;
        RECT 2459.330 304.690 2460.510 305.870 ;
        RECT 2457.730 303.090 2458.910 304.270 ;
        RECT 2459.330 303.090 2460.510 304.270 ;
        RECT 2457.730 124.690 2458.910 125.870 ;
        RECT 2459.330 124.690 2460.510 125.870 ;
        RECT 2457.730 123.090 2458.910 124.270 ;
        RECT 2459.330 123.090 2460.510 124.270 ;
        RECT 2457.730 -17.310 2458.910 -16.130 ;
        RECT 2459.330 -17.310 2460.510 -16.130 ;
        RECT 2457.730 -18.910 2458.910 -17.730 ;
        RECT 2459.330 -18.910 2460.510 -17.730 ;
        RECT 2637.730 3537.410 2638.910 3538.590 ;
        RECT 2639.330 3537.410 2640.510 3538.590 ;
        RECT 2637.730 3535.810 2638.910 3536.990 ;
        RECT 2639.330 3535.810 2640.510 3536.990 ;
        RECT 2637.730 3364.690 2638.910 3365.870 ;
        RECT 2639.330 3364.690 2640.510 3365.870 ;
        RECT 2637.730 3363.090 2638.910 3364.270 ;
        RECT 2639.330 3363.090 2640.510 3364.270 ;
        RECT 2637.730 3184.690 2638.910 3185.870 ;
        RECT 2639.330 3184.690 2640.510 3185.870 ;
        RECT 2637.730 3183.090 2638.910 3184.270 ;
        RECT 2639.330 3183.090 2640.510 3184.270 ;
        RECT 2637.730 3004.690 2638.910 3005.870 ;
        RECT 2639.330 3004.690 2640.510 3005.870 ;
        RECT 2637.730 3003.090 2638.910 3004.270 ;
        RECT 2639.330 3003.090 2640.510 3004.270 ;
        RECT 2637.730 2824.690 2638.910 2825.870 ;
        RECT 2639.330 2824.690 2640.510 2825.870 ;
        RECT 2637.730 2823.090 2638.910 2824.270 ;
        RECT 2639.330 2823.090 2640.510 2824.270 ;
        RECT 2637.730 2644.690 2638.910 2645.870 ;
        RECT 2639.330 2644.690 2640.510 2645.870 ;
        RECT 2637.730 2643.090 2638.910 2644.270 ;
        RECT 2639.330 2643.090 2640.510 2644.270 ;
        RECT 2637.730 2464.690 2638.910 2465.870 ;
        RECT 2639.330 2464.690 2640.510 2465.870 ;
        RECT 2637.730 2463.090 2638.910 2464.270 ;
        RECT 2639.330 2463.090 2640.510 2464.270 ;
        RECT 2637.730 2284.690 2638.910 2285.870 ;
        RECT 2639.330 2284.690 2640.510 2285.870 ;
        RECT 2637.730 2283.090 2638.910 2284.270 ;
        RECT 2639.330 2283.090 2640.510 2284.270 ;
        RECT 2637.730 2104.690 2638.910 2105.870 ;
        RECT 2639.330 2104.690 2640.510 2105.870 ;
        RECT 2637.730 2103.090 2638.910 2104.270 ;
        RECT 2639.330 2103.090 2640.510 2104.270 ;
        RECT 2637.730 1924.690 2638.910 1925.870 ;
        RECT 2639.330 1924.690 2640.510 1925.870 ;
        RECT 2637.730 1923.090 2638.910 1924.270 ;
        RECT 2639.330 1923.090 2640.510 1924.270 ;
        RECT 2637.730 1744.690 2638.910 1745.870 ;
        RECT 2639.330 1744.690 2640.510 1745.870 ;
        RECT 2637.730 1743.090 2638.910 1744.270 ;
        RECT 2639.330 1743.090 2640.510 1744.270 ;
        RECT 2637.730 1564.690 2638.910 1565.870 ;
        RECT 2639.330 1564.690 2640.510 1565.870 ;
        RECT 2637.730 1563.090 2638.910 1564.270 ;
        RECT 2639.330 1563.090 2640.510 1564.270 ;
        RECT 2637.730 1384.690 2638.910 1385.870 ;
        RECT 2639.330 1384.690 2640.510 1385.870 ;
        RECT 2637.730 1383.090 2638.910 1384.270 ;
        RECT 2639.330 1383.090 2640.510 1384.270 ;
        RECT 2637.730 1204.690 2638.910 1205.870 ;
        RECT 2639.330 1204.690 2640.510 1205.870 ;
        RECT 2637.730 1203.090 2638.910 1204.270 ;
        RECT 2639.330 1203.090 2640.510 1204.270 ;
        RECT 2637.730 1024.690 2638.910 1025.870 ;
        RECT 2639.330 1024.690 2640.510 1025.870 ;
        RECT 2637.730 1023.090 2638.910 1024.270 ;
        RECT 2639.330 1023.090 2640.510 1024.270 ;
        RECT 2637.730 844.690 2638.910 845.870 ;
        RECT 2639.330 844.690 2640.510 845.870 ;
        RECT 2637.730 843.090 2638.910 844.270 ;
        RECT 2639.330 843.090 2640.510 844.270 ;
        RECT 2637.730 664.690 2638.910 665.870 ;
        RECT 2639.330 664.690 2640.510 665.870 ;
        RECT 2637.730 663.090 2638.910 664.270 ;
        RECT 2639.330 663.090 2640.510 664.270 ;
        RECT 2637.730 484.690 2638.910 485.870 ;
        RECT 2639.330 484.690 2640.510 485.870 ;
        RECT 2637.730 483.090 2638.910 484.270 ;
        RECT 2639.330 483.090 2640.510 484.270 ;
        RECT 2637.730 304.690 2638.910 305.870 ;
        RECT 2639.330 304.690 2640.510 305.870 ;
        RECT 2637.730 303.090 2638.910 304.270 ;
        RECT 2639.330 303.090 2640.510 304.270 ;
        RECT 2637.730 124.690 2638.910 125.870 ;
        RECT 2639.330 124.690 2640.510 125.870 ;
        RECT 2637.730 123.090 2638.910 124.270 ;
        RECT 2639.330 123.090 2640.510 124.270 ;
        RECT 2637.730 -17.310 2638.910 -16.130 ;
        RECT 2639.330 -17.310 2640.510 -16.130 ;
        RECT 2637.730 -18.910 2638.910 -17.730 ;
        RECT 2639.330 -18.910 2640.510 -17.730 ;
        RECT 2817.730 3537.410 2818.910 3538.590 ;
        RECT 2819.330 3537.410 2820.510 3538.590 ;
        RECT 2817.730 3535.810 2818.910 3536.990 ;
        RECT 2819.330 3535.810 2820.510 3536.990 ;
        RECT 2817.730 3364.690 2818.910 3365.870 ;
        RECT 2819.330 3364.690 2820.510 3365.870 ;
        RECT 2817.730 3363.090 2818.910 3364.270 ;
        RECT 2819.330 3363.090 2820.510 3364.270 ;
        RECT 2817.730 3184.690 2818.910 3185.870 ;
        RECT 2819.330 3184.690 2820.510 3185.870 ;
        RECT 2817.730 3183.090 2818.910 3184.270 ;
        RECT 2819.330 3183.090 2820.510 3184.270 ;
        RECT 2817.730 3004.690 2818.910 3005.870 ;
        RECT 2819.330 3004.690 2820.510 3005.870 ;
        RECT 2817.730 3003.090 2818.910 3004.270 ;
        RECT 2819.330 3003.090 2820.510 3004.270 ;
        RECT 2817.730 2824.690 2818.910 2825.870 ;
        RECT 2819.330 2824.690 2820.510 2825.870 ;
        RECT 2817.730 2823.090 2818.910 2824.270 ;
        RECT 2819.330 2823.090 2820.510 2824.270 ;
        RECT 2817.730 2644.690 2818.910 2645.870 ;
        RECT 2819.330 2644.690 2820.510 2645.870 ;
        RECT 2817.730 2643.090 2818.910 2644.270 ;
        RECT 2819.330 2643.090 2820.510 2644.270 ;
        RECT 2817.730 2464.690 2818.910 2465.870 ;
        RECT 2819.330 2464.690 2820.510 2465.870 ;
        RECT 2817.730 2463.090 2818.910 2464.270 ;
        RECT 2819.330 2463.090 2820.510 2464.270 ;
        RECT 2817.730 2284.690 2818.910 2285.870 ;
        RECT 2819.330 2284.690 2820.510 2285.870 ;
        RECT 2817.730 2283.090 2818.910 2284.270 ;
        RECT 2819.330 2283.090 2820.510 2284.270 ;
        RECT 2817.730 2104.690 2818.910 2105.870 ;
        RECT 2819.330 2104.690 2820.510 2105.870 ;
        RECT 2817.730 2103.090 2818.910 2104.270 ;
        RECT 2819.330 2103.090 2820.510 2104.270 ;
        RECT 2817.730 1924.690 2818.910 1925.870 ;
        RECT 2819.330 1924.690 2820.510 1925.870 ;
        RECT 2817.730 1923.090 2818.910 1924.270 ;
        RECT 2819.330 1923.090 2820.510 1924.270 ;
        RECT 2817.730 1744.690 2818.910 1745.870 ;
        RECT 2819.330 1744.690 2820.510 1745.870 ;
        RECT 2817.730 1743.090 2818.910 1744.270 ;
        RECT 2819.330 1743.090 2820.510 1744.270 ;
        RECT 2817.730 1564.690 2818.910 1565.870 ;
        RECT 2819.330 1564.690 2820.510 1565.870 ;
        RECT 2817.730 1563.090 2818.910 1564.270 ;
        RECT 2819.330 1563.090 2820.510 1564.270 ;
        RECT 2817.730 1384.690 2818.910 1385.870 ;
        RECT 2819.330 1384.690 2820.510 1385.870 ;
        RECT 2817.730 1383.090 2818.910 1384.270 ;
        RECT 2819.330 1383.090 2820.510 1384.270 ;
        RECT 2817.730 1204.690 2818.910 1205.870 ;
        RECT 2819.330 1204.690 2820.510 1205.870 ;
        RECT 2817.730 1203.090 2818.910 1204.270 ;
        RECT 2819.330 1203.090 2820.510 1204.270 ;
        RECT 2817.730 1024.690 2818.910 1025.870 ;
        RECT 2819.330 1024.690 2820.510 1025.870 ;
        RECT 2817.730 1023.090 2818.910 1024.270 ;
        RECT 2819.330 1023.090 2820.510 1024.270 ;
        RECT 2817.730 844.690 2818.910 845.870 ;
        RECT 2819.330 844.690 2820.510 845.870 ;
        RECT 2817.730 843.090 2818.910 844.270 ;
        RECT 2819.330 843.090 2820.510 844.270 ;
        RECT 2817.730 664.690 2818.910 665.870 ;
        RECT 2819.330 664.690 2820.510 665.870 ;
        RECT 2817.730 663.090 2818.910 664.270 ;
        RECT 2819.330 663.090 2820.510 664.270 ;
        RECT 2817.730 484.690 2818.910 485.870 ;
        RECT 2819.330 484.690 2820.510 485.870 ;
        RECT 2817.730 483.090 2818.910 484.270 ;
        RECT 2819.330 483.090 2820.510 484.270 ;
        RECT 2817.730 304.690 2818.910 305.870 ;
        RECT 2819.330 304.690 2820.510 305.870 ;
        RECT 2817.730 303.090 2818.910 304.270 ;
        RECT 2819.330 303.090 2820.510 304.270 ;
        RECT 2817.730 124.690 2818.910 125.870 ;
        RECT 2819.330 124.690 2820.510 125.870 ;
        RECT 2817.730 123.090 2818.910 124.270 ;
        RECT 2819.330 123.090 2820.510 124.270 ;
        RECT 2817.730 -17.310 2818.910 -16.130 ;
        RECT 2819.330 -17.310 2820.510 -16.130 ;
        RECT 2817.730 -18.910 2818.910 -17.730 ;
        RECT 2819.330 -18.910 2820.510 -17.730 ;
        RECT 2941.110 3537.410 2942.290 3538.590 ;
        RECT 2942.710 3537.410 2943.890 3538.590 ;
        RECT 2941.110 3535.810 2942.290 3536.990 ;
        RECT 2942.710 3535.810 2943.890 3536.990 ;
        RECT 2941.110 3364.690 2942.290 3365.870 ;
        RECT 2942.710 3364.690 2943.890 3365.870 ;
        RECT 2941.110 3363.090 2942.290 3364.270 ;
        RECT 2942.710 3363.090 2943.890 3364.270 ;
        RECT 2941.110 3184.690 2942.290 3185.870 ;
        RECT 2942.710 3184.690 2943.890 3185.870 ;
        RECT 2941.110 3183.090 2942.290 3184.270 ;
        RECT 2942.710 3183.090 2943.890 3184.270 ;
        RECT 2941.110 3004.690 2942.290 3005.870 ;
        RECT 2942.710 3004.690 2943.890 3005.870 ;
        RECT 2941.110 3003.090 2942.290 3004.270 ;
        RECT 2942.710 3003.090 2943.890 3004.270 ;
        RECT 2941.110 2824.690 2942.290 2825.870 ;
        RECT 2942.710 2824.690 2943.890 2825.870 ;
        RECT 2941.110 2823.090 2942.290 2824.270 ;
        RECT 2942.710 2823.090 2943.890 2824.270 ;
        RECT 2941.110 2644.690 2942.290 2645.870 ;
        RECT 2942.710 2644.690 2943.890 2645.870 ;
        RECT 2941.110 2643.090 2942.290 2644.270 ;
        RECT 2942.710 2643.090 2943.890 2644.270 ;
        RECT 2941.110 2464.690 2942.290 2465.870 ;
        RECT 2942.710 2464.690 2943.890 2465.870 ;
        RECT 2941.110 2463.090 2942.290 2464.270 ;
        RECT 2942.710 2463.090 2943.890 2464.270 ;
        RECT 2941.110 2284.690 2942.290 2285.870 ;
        RECT 2942.710 2284.690 2943.890 2285.870 ;
        RECT 2941.110 2283.090 2942.290 2284.270 ;
        RECT 2942.710 2283.090 2943.890 2284.270 ;
        RECT 2941.110 2104.690 2942.290 2105.870 ;
        RECT 2942.710 2104.690 2943.890 2105.870 ;
        RECT 2941.110 2103.090 2942.290 2104.270 ;
        RECT 2942.710 2103.090 2943.890 2104.270 ;
        RECT 2941.110 1924.690 2942.290 1925.870 ;
        RECT 2942.710 1924.690 2943.890 1925.870 ;
        RECT 2941.110 1923.090 2942.290 1924.270 ;
        RECT 2942.710 1923.090 2943.890 1924.270 ;
        RECT 2941.110 1744.690 2942.290 1745.870 ;
        RECT 2942.710 1744.690 2943.890 1745.870 ;
        RECT 2941.110 1743.090 2942.290 1744.270 ;
        RECT 2942.710 1743.090 2943.890 1744.270 ;
        RECT 2941.110 1564.690 2942.290 1565.870 ;
        RECT 2942.710 1564.690 2943.890 1565.870 ;
        RECT 2941.110 1563.090 2942.290 1564.270 ;
        RECT 2942.710 1563.090 2943.890 1564.270 ;
        RECT 2941.110 1384.690 2942.290 1385.870 ;
        RECT 2942.710 1384.690 2943.890 1385.870 ;
        RECT 2941.110 1383.090 2942.290 1384.270 ;
        RECT 2942.710 1383.090 2943.890 1384.270 ;
        RECT 2941.110 1204.690 2942.290 1205.870 ;
        RECT 2942.710 1204.690 2943.890 1205.870 ;
        RECT 2941.110 1203.090 2942.290 1204.270 ;
        RECT 2942.710 1203.090 2943.890 1204.270 ;
        RECT 2941.110 1024.690 2942.290 1025.870 ;
        RECT 2942.710 1024.690 2943.890 1025.870 ;
        RECT 2941.110 1023.090 2942.290 1024.270 ;
        RECT 2942.710 1023.090 2943.890 1024.270 ;
        RECT 2941.110 844.690 2942.290 845.870 ;
        RECT 2942.710 844.690 2943.890 845.870 ;
        RECT 2941.110 843.090 2942.290 844.270 ;
        RECT 2942.710 843.090 2943.890 844.270 ;
        RECT 2941.110 664.690 2942.290 665.870 ;
        RECT 2942.710 664.690 2943.890 665.870 ;
        RECT 2941.110 663.090 2942.290 664.270 ;
        RECT 2942.710 663.090 2943.890 664.270 ;
        RECT 2941.110 484.690 2942.290 485.870 ;
        RECT 2942.710 484.690 2943.890 485.870 ;
        RECT 2941.110 483.090 2942.290 484.270 ;
        RECT 2942.710 483.090 2943.890 484.270 ;
        RECT 2941.110 304.690 2942.290 305.870 ;
        RECT 2942.710 304.690 2943.890 305.870 ;
        RECT 2941.110 303.090 2942.290 304.270 ;
        RECT 2942.710 303.090 2943.890 304.270 ;
        RECT 2941.110 124.690 2942.290 125.870 ;
        RECT 2942.710 124.690 2943.890 125.870 ;
        RECT 2941.110 123.090 2942.290 124.270 ;
        RECT 2942.710 123.090 2943.890 124.270 ;
        RECT 2941.110 -17.310 2942.290 -16.130 ;
        RECT 2942.710 -17.310 2943.890 -16.130 ;
        RECT 2941.110 -18.910 2942.290 -17.730 ;
        RECT 2942.710 -18.910 2943.890 -17.730 ;
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
        RECT -24.430 842.930 2944.050 846.030 ;
        RECT -24.430 662.930 2944.050 666.030 ;
        RECT -24.430 482.930 2944.050 486.030 ;
        RECT -24.430 302.930 2944.050 306.030 ;
        RECT -24.430 122.930 2944.050 126.030 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 201.090 303.520 201.410 303.580 ;
        RECT 202.010 303.520 202.330 303.580 ;
        RECT 201.090 303.380 202.330 303.520 ;
        RECT 201.090 303.320 201.410 303.380 ;
        RECT 202.010 303.320 202.330 303.380 ;
      LAYER via ;
        RECT 201.120 303.320 201.380 303.580 ;
        RECT 202.040 303.320 202.300 303.580 ;
      LAYER met2 ;
        RECT 201.930 400.180 202.210 404.000 ;
        RECT 201.930 400.000 202.240 400.180 ;
        RECT 202.100 303.610 202.240 400.000 ;
        RECT 201.120 303.290 201.380 303.610 ;
        RECT 202.040 303.290 202.300 303.610 ;
        RECT 201.180 16.845 201.320 303.290 ;
        RECT 8.370 16.475 8.650 16.845 ;
        RECT 201.110 16.475 201.390 16.845 ;
        RECT 8.440 2.400 8.580 16.475 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 8.370 16.520 8.650 16.800 ;
        RECT 201.110 16.520 201.390 16.800 ;
      LAYER met3 ;
        RECT 8.345 16.810 8.675 16.825 ;
        RECT 201.085 16.810 201.415 16.825 ;
        RECT 8.345 16.510 201.415 16.810 ;
        RECT 8.345 16.495 8.675 16.510 ;
        RECT 201.085 16.495 201.415 16.510 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 200.630 386.480 200.950 386.540 ;
        RECT 202.470 386.480 202.790 386.540 ;
        RECT 200.630 386.340 202.790 386.480 ;
        RECT 200.630 386.280 200.950 386.340 ;
        RECT 202.470 386.280 202.790 386.340 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 200.630 17.580 200.950 17.640 ;
        RECT 14.330 17.440 200.950 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 200.630 17.380 200.950 17.440 ;
      LAYER via ;
        RECT 200.660 386.280 200.920 386.540 ;
        RECT 202.500 386.280 202.760 386.540 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 200.660 17.380 200.920 17.640 ;
      LAYER met2 ;
        RECT 203.770 400.250 204.050 404.000 ;
        RECT 202.560 400.110 204.050 400.250 ;
        RECT 202.560 386.570 202.700 400.110 ;
        RECT 203.770 400.000 204.050 400.110 ;
        RECT 200.660 386.250 200.920 386.570 ;
        RECT 202.500 386.250 202.760 386.570 ;
        RECT 200.720 17.670 200.860 386.250 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 200.660 17.350 200.920 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 208.910 17.920 209.230 17.980 ;
        RECT 38.250 17.780 209.230 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 208.910 17.720 209.230 17.780 ;
      LAYER via ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 208.940 17.720 209.200 17.980 ;
      LAYER met2 ;
        RECT 211.130 400.250 211.410 404.000 ;
        RECT 209.920 400.110 211.410 400.250 ;
        RECT 209.920 324.370 210.060 400.110 ;
        RECT 211.130 400.000 211.410 400.110 ;
        RECT 209.000 324.230 210.060 324.370 ;
        RECT 209.000 18.010 209.140 324.230 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 208.940 17.690 209.200 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 239.270 15.200 239.590 15.260 ;
        RECT 270.090 15.200 270.410 15.260 ;
        RECT 239.270 15.060 270.410 15.200 ;
        RECT 239.270 15.000 239.590 15.060 ;
        RECT 270.090 15.000 270.410 15.060 ;
      LAYER via ;
        RECT 239.300 15.000 239.560 15.260 ;
        RECT 270.120 15.000 270.380 15.260 ;
      LAYER met2 ;
        RECT 272.770 400.250 273.050 404.000 ;
        RECT 271.560 400.110 273.050 400.250 ;
        RECT 271.560 324.370 271.700 400.110 ;
        RECT 272.770 400.000 273.050 400.110 ;
        RECT 270.180 324.230 271.700 324.370 ;
        RECT 270.180 15.290 270.320 324.230 ;
        RECT 239.300 14.970 239.560 15.290 ;
        RECT 270.120 14.970 270.380 15.290 ;
        RECT 239.360 2.400 239.500 14.970 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 255.370 386.820 255.690 386.880 ;
        RECT 278.370 386.820 278.690 386.880 ;
        RECT 255.370 386.680 278.690 386.820 ;
        RECT 255.370 386.620 255.690 386.680 ;
        RECT 278.370 386.620 278.690 386.680 ;
      LAYER via ;
        RECT 255.400 386.620 255.660 386.880 ;
        RECT 278.400 386.620 278.660 386.880 ;
      LAYER met2 ;
        RECT 278.290 400.180 278.570 404.000 ;
        RECT 278.290 400.000 278.600 400.180 ;
        RECT 278.460 386.910 278.600 400.000 ;
        RECT 255.400 386.590 255.660 386.910 ;
        RECT 278.400 386.590 278.660 386.910 ;
        RECT 255.460 1.770 255.600 386.590 ;
        RECT 256.630 1.770 257.190 2.400 ;
        RECT 255.460 1.630 257.190 1.770 ;
        RECT 256.630 -4.800 257.190 1.630 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 274.690 20.300 275.010 20.360 ;
        RECT 283.430 20.300 283.750 20.360 ;
        RECT 274.690 20.160 283.750 20.300 ;
        RECT 274.690 20.100 275.010 20.160 ;
        RECT 283.430 20.100 283.750 20.160 ;
      LAYER via ;
        RECT 274.720 20.100 274.980 20.360 ;
        RECT 283.460 20.100 283.720 20.360 ;
      LAYER met2 ;
        RECT 283.810 400.250 284.090 404.000 ;
        RECT 283.520 400.110 284.090 400.250 ;
        RECT 283.520 20.390 283.660 400.110 ;
        RECT 283.810 400.000 284.090 400.110 ;
        RECT 274.720 20.070 274.980 20.390 ;
        RECT 283.460 20.070 283.720 20.390 ;
        RECT 274.780 2.400 274.920 20.070 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.330 400.180 289.610 404.000 ;
        RECT 289.330 400.000 289.640 400.180 ;
        RECT 289.500 386.470 289.640 400.000 ;
        RECT 289.500 386.330 290.100 386.470 ;
        RECT 289.960 17.410 290.100 386.330 ;
        RECT 289.960 17.270 292.400 17.410 ;
        RECT 292.260 2.400 292.400 17.270 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.330 386.140 290.650 386.200 ;
        RECT 293.550 386.140 293.870 386.200 ;
        RECT 290.330 386.000 293.870 386.140 ;
        RECT 290.330 385.940 290.650 386.000 ;
        RECT 293.550 385.940 293.870 386.000 ;
        RECT 290.330 18.600 290.650 18.660 ;
        RECT 310.110 18.600 310.430 18.660 ;
        RECT 290.330 18.460 310.430 18.600 ;
        RECT 290.330 18.400 290.650 18.460 ;
        RECT 310.110 18.400 310.430 18.460 ;
      LAYER via ;
        RECT 290.360 385.940 290.620 386.200 ;
        RECT 293.580 385.940 293.840 386.200 ;
        RECT 290.360 18.400 290.620 18.660 ;
        RECT 310.140 18.400 310.400 18.660 ;
      LAYER met2 ;
        RECT 294.850 400.250 295.130 404.000 ;
        RECT 293.640 400.110 295.130 400.250 ;
        RECT 293.640 386.230 293.780 400.110 ;
        RECT 294.850 400.000 295.130 400.110 ;
        RECT 290.360 385.910 290.620 386.230 ;
        RECT 293.580 385.910 293.840 386.230 ;
        RECT 290.420 18.690 290.560 385.910 ;
        RECT 290.360 18.370 290.620 18.690 ;
        RECT 310.140 18.370 310.400 18.690 ;
        RECT 310.200 2.400 310.340 18.370 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 300.450 386.480 300.770 386.540 ;
        RECT 306.890 386.480 307.210 386.540 ;
        RECT 300.450 386.340 307.210 386.480 ;
        RECT 300.450 386.280 300.770 386.340 ;
        RECT 306.890 386.280 307.210 386.340 ;
        RECT 306.890 20.640 307.210 20.700 ;
        RECT 325.750 20.640 326.070 20.700 ;
        RECT 306.890 20.500 326.070 20.640 ;
        RECT 306.890 20.440 307.210 20.500 ;
        RECT 325.750 20.440 326.070 20.500 ;
      LAYER via ;
        RECT 300.480 386.280 300.740 386.540 ;
        RECT 306.920 386.280 307.180 386.540 ;
        RECT 306.920 20.440 307.180 20.700 ;
        RECT 325.780 20.440 326.040 20.700 ;
      LAYER met2 ;
        RECT 300.370 400.180 300.650 404.000 ;
        RECT 300.370 400.000 300.680 400.180 ;
        RECT 300.540 386.570 300.680 400.000 ;
        RECT 300.480 386.250 300.740 386.570 ;
        RECT 306.920 386.250 307.180 386.570 ;
        RECT 306.980 20.730 307.120 386.250 ;
        RECT 306.920 20.410 307.180 20.730 ;
        RECT 325.780 20.410 326.040 20.730 ;
        RECT 325.840 1.770 325.980 20.410 ;
        RECT 327.470 1.770 328.030 2.400 ;
        RECT 325.840 1.630 328.030 1.770 ;
        RECT 327.470 -4.800 328.030 1.630 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 303.670 376.280 303.990 376.340 ;
        RECT 305.050 376.280 305.370 376.340 ;
        RECT 303.670 376.140 305.370 376.280 ;
        RECT 303.670 376.080 303.990 376.140 ;
        RECT 305.050 376.080 305.370 376.140 ;
        RECT 303.670 19.620 303.990 19.680 ;
        RECT 345.530 19.620 345.850 19.680 ;
        RECT 303.670 19.480 345.850 19.620 ;
        RECT 303.670 19.420 303.990 19.480 ;
        RECT 345.530 19.420 345.850 19.480 ;
      LAYER via ;
        RECT 303.700 376.080 303.960 376.340 ;
        RECT 305.080 376.080 305.340 376.340 ;
        RECT 303.700 19.420 303.960 19.680 ;
        RECT 345.560 19.420 345.820 19.680 ;
      LAYER met2 ;
        RECT 305.430 400.250 305.710 404.000 ;
        RECT 305.140 400.110 305.710 400.250 ;
        RECT 305.140 376.370 305.280 400.110 ;
        RECT 305.430 400.000 305.710 400.110 ;
        RECT 303.700 376.050 303.960 376.370 ;
        RECT 305.080 376.050 305.340 376.370 ;
        RECT 303.760 19.710 303.900 376.050 ;
        RECT 303.700 19.390 303.960 19.710 ;
        RECT 345.560 19.390 345.820 19.710 ;
        RECT 345.620 2.400 345.760 19.390 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.030 17.240 311.350 17.300 ;
        RECT 363.010 17.240 363.330 17.300 ;
        RECT 311.030 17.100 363.330 17.240 ;
        RECT 311.030 17.040 311.350 17.100 ;
        RECT 363.010 17.040 363.330 17.100 ;
      LAYER via ;
        RECT 311.060 17.040 311.320 17.300 ;
        RECT 363.040 17.040 363.300 17.300 ;
      LAYER met2 ;
        RECT 310.950 400.180 311.230 404.000 ;
        RECT 310.950 400.000 311.260 400.180 ;
        RECT 311.120 17.330 311.260 400.000 ;
        RECT 311.060 17.010 311.320 17.330 ;
        RECT 363.040 17.010 363.300 17.330 ;
        RECT 363.100 2.400 363.240 17.010 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 316.550 392.260 316.870 392.320 ;
        RECT 379.570 392.260 379.890 392.320 ;
        RECT 316.550 392.120 379.890 392.260 ;
        RECT 316.550 392.060 316.870 392.120 ;
        RECT 379.570 392.060 379.890 392.120 ;
      LAYER via ;
        RECT 316.580 392.060 316.840 392.320 ;
        RECT 379.600 392.060 379.860 392.320 ;
      LAYER met2 ;
        RECT 316.470 400.180 316.750 404.000 ;
        RECT 316.470 400.000 316.780 400.180 ;
        RECT 316.640 392.350 316.780 400.000 ;
        RECT 316.580 392.030 316.840 392.350 ;
        RECT 379.600 392.030 379.860 392.350 ;
        RECT 379.660 1.770 379.800 392.030 ;
        RECT 380.830 1.770 381.390 2.400 ;
        RECT 379.660 1.630 381.390 1.770 ;
        RECT 380.830 -4.800 381.390 1.630 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 322.070 391.240 322.390 391.300 ;
        RECT 393.370 391.240 393.690 391.300 ;
        RECT 322.070 391.100 393.690 391.240 ;
        RECT 322.070 391.040 322.390 391.100 ;
        RECT 393.370 391.040 393.690 391.100 ;
      LAYER via ;
        RECT 322.100 391.040 322.360 391.300 ;
        RECT 393.400 391.040 393.660 391.300 ;
      LAYER met2 ;
        RECT 321.990 400.180 322.270 404.000 ;
        RECT 321.990 400.000 322.300 400.180 ;
        RECT 322.160 391.330 322.300 400.000 ;
        RECT 322.100 391.010 322.360 391.330 ;
        RECT 393.400 391.010 393.660 391.330 ;
        RECT 393.460 3.130 393.600 391.010 ;
        RECT 393.460 2.990 396.360 3.130 ;
        RECT 396.220 1.770 396.360 2.990 ;
        RECT 398.310 1.770 398.870 2.400 ;
        RECT 396.220 1.630 398.870 1.770 ;
        RECT 398.310 -4.800 398.870 1.630 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 61.710 19.280 62.030 19.340 ;
        RECT 215.350 19.280 215.670 19.340 ;
        RECT 61.710 19.140 215.670 19.280 ;
        RECT 61.710 19.080 62.030 19.140 ;
        RECT 215.350 19.080 215.670 19.140 ;
      LAYER via ;
        RECT 61.740 19.080 62.000 19.340 ;
        RECT 215.380 19.080 215.640 19.340 ;
      LAYER met2 ;
        RECT 218.490 400.250 218.770 404.000 ;
        RECT 217.280 400.110 218.770 400.250 ;
        RECT 217.280 324.370 217.420 400.110 ;
        RECT 218.490 400.000 218.770 400.110 ;
        RECT 215.440 324.230 217.420 324.370 ;
        RECT 215.440 19.370 215.580 324.230 ;
        RECT 61.740 19.050 62.000 19.370 ;
        RECT 215.380 19.050 215.640 19.370 ;
        RECT 61.800 2.400 61.940 19.050 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 325.290 25.400 325.610 25.460 ;
        RECT 416.370 25.400 416.690 25.460 ;
        RECT 325.290 25.260 416.690 25.400 ;
        RECT 325.290 25.200 325.610 25.260 ;
        RECT 416.370 25.200 416.690 25.260 ;
      LAYER via ;
        RECT 325.320 25.200 325.580 25.460 ;
        RECT 416.400 25.200 416.660 25.460 ;
      LAYER met2 ;
        RECT 327.510 400.250 327.790 404.000 ;
        RECT 326.300 400.110 327.790 400.250 ;
        RECT 326.300 303.670 326.440 400.110 ;
        RECT 327.510 400.000 327.790 400.110 ;
        RECT 325.380 303.530 326.440 303.670 ;
        RECT 325.380 25.490 325.520 303.530 ;
        RECT 325.320 25.170 325.580 25.490 ;
        RECT 416.400 25.170 416.660 25.490 ;
        RECT 416.460 2.400 416.600 25.170 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.730 25.060 332.050 25.120 ;
        RECT 434.310 25.060 434.630 25.120 ;
        RECT 331.730 24.920 434.630 25.060 ;
        RECT 331.730 24.860 332.050 24.920 ;
        RECT 434.310 24.860 434.630 24.920 ;
      LAYER via ;
        RECT 331.760 24.860 332.020 25.120 ;
        RECT 434.340 24.860 434.600 25.120 ;
      LAYER met2 ;
        RECT 333.030 400.250 333.310 404.000 ;
        RECT 331.820 400.110 333.310 400.250 ;
        RECT 331.820 25.150 331.960 400.110 ;
        RECT 333.030 400.000 333.310 400.110 ;
        RECT 331.760 24.830 332.020 25.150 ;
        RECT 434.340 24.830 434.600 25.150 ;
        RECT 434.400 2.400 434.540 24.830 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 338.630 24.720 338.950 24.780 ;
        RECT 451.790 24.720 452.110 24.780 ;
        RECT 338.630 24.580 452.110 24.720 ;
        RECT 338.630 24.520 338.950 24.580 ;
        RECT 451.790 24.520 452.110 24.580 ;
      LAYER via ;
        RECT 338.660 24.520 338.920 24.780 ;
        RECT 451.820 24.520 452.080 24.780 ;
      LAYER met2 ;
        RECT 338.090 400.250 338.370 404.000 ;
        RECT 338.090 400.110 338.860 400.250 ;
        RECT 338.090 400.000 338.370 400.110 ;
        RECT 338.720 24.810 338.860 400.110 ;
        RECT 338.660 24.490 338.920 24.810 ;
        RECT 451.820 24.490 452.080 24.810 ;
        RECT 451.880 2.400 452.020 24.490 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 339.090 375.600 339.410 375.660 ;
        RECT 342.310 375.600 342.630 375.660 ;
        RECT 339.090 375.460 342.630 375.600 ;
        RECT 339.090 375.400 339.410 375.460 ;
        RECT 342.310 375.400 342.630 375.460 ;
        RECT 339.090 24.380 339.410 24.440 ;
        RECT 469.730 24.380 470.050 24.440 ;
        RECT 339.090 24.240 470.050 24.380 ;
        RECT 339.090 24.180 339.410 24.240 ;
        RECT 469.730 24.180 470.050 24.240 ;
      LAYER via ;
        RECT 339.120 375.400 339.380 375.660 ;
        RECT 342.340 375.400 342.600 375.660 ;
        RECT 339.120 24.180 339.380 24.440 ;
        RECT 469.760 24.180 470.020 24.440 ;
      LAYER met2 ;
        RECT 343.610 400.250 343.890 404.000 ;
        RECT 342.400 400.110 343.890 400.250 ;
        RECT 342.400 375.690 342.540 400.110 ;
        RECT 343.610 400.000 343.890 400.110 ;
        RECT 339.120 375.370 339.380 375.690 ;
        RECT 342.340 375.370 342.600 375.690 ;
        RECT 339.180 24.470 339.320 375.370 ;
        RECT 339.120 24.150 339.380 24.470 ;
        RECT 469.760 24.150 470.020 24.470 ;
        RECT 469.820 2.400 469.960 24.150 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 349.210 388.180 349.530 388.240 ;
        RECT 410.390 388.180 410.710 388.240 ;
        RECT 349.210 388.040 410.710 388.180 ;
        RECT 349.210 387.980 349.530 388.040 ;
        RECT 410.390 387.980 410.710 388.040 ;
        RECT 487.210 15.880 487.530 15.940 ;
        RECT 469.130 15.740 487.530 15.880 ;
        RECT 410.850 15.540 411.170 15.600 ;
        RECT 469.130 15.540 469.270 15.740 ;
        RECT 487.210 15.680 487.530 15.740 ;
        RECT 410.850 15.400 469.270 15.540 ;
        RECT 410.850 15.340 411.170 15.400 ;
      LAYER via ;
        RECT 349.240 387.980 349.500 388.240 ;
        RECT 410.420 387.980 410.680 388.240 ;
        RECT 410.880 15.340 411.140 15.600 ;
        RECT 487.240 15.680 487.500 15.940 ;
      LAYER met2 ;
        RECT 349.130 400.180 349.410 404.000 ;
        RECT 349.130 400.000 349.440 400.180 ;
        RECT 349.300 388.270 349.440 400.000 ;
        RECT 349.240 387.950 349.500 388.270 ;
        RECT 410.420 387.950 410.680 388.270 ;
        RECT 410.480 82.870 410.620 387.950 ;
        RECT 410.480 82.730 411.080 82.870 ;
        RECT 410.940 15.630 411.080 82.730 ;
        RECT 487.240 15.650 487.500 15.970 ;
        RECT 410.880 15.310 411.140 15.630 ;
        RECT 487.300 2.400 487.440 15.650 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.430 18.260 352.750 18.320 ;
        RECT 503.310 18.260 503.630 18.320 ;
        RECT 352.430 18.120 503.630 18.260 ;
        RECT 352.430 18.060 352.750 18.120 ;
        RECT 503.310 18.060 503.630 18.120 ;
      LAYER via ;
        RECT 352.460 18.060 352.720 18.320 ;
        RECT 503.340 18.060 503.600 18.320 ;
      LAYER met2 ;
        RECT 354.650 400.250 354.930 404.000 ;
        RECT 353.440 400.110 354.930 400.250 ;
        RECT 353.440 386.480 353.580 400.110 ;
        RECT 354.650 400.000 354.930 400.110 ;
        RECT 352.520 386.340 353.580 386.480 ;
        RECT 352.520 18.350 352.660 386.340 ;
        RECT 352.460 18.030 352.720 18.350 ;
        RECT 503.340 18.030 503.600 18.350 ;
        RECT 503.400 17.410 503.540 18.030 ;
        RECT 503.400 17.270 504.000 17.410 ;
        RECT 503.860 1.770 504.000 17.270 ;
        RECT 505.030 1.770 505.590 2.400 ;
        RECT 503.860 1.630 505.590 1.770 ;
        RECT 505.030 -4.800 505.590 1.630 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 360.250 389.540 360.570 389.600 ;
        RECT 432.010 389.540 432.330 389.600 ;
        RECT 360.250 389.400 432.330 389.540 ;
        RECT 360.250 389.340 360.570 389.400 ;
        RECT 432.010 389.340 432.330 389.400 ;
        RECT 431.090 16.900 431.410 16.960 ;
        RECT 431.090 16.760 469.270 16.900 ;
        RECT 431.090 16.700 431.410 16.760 ;
        RECT 469.130 16.560 469.270 16.760 ;
        RECT 522.630 16.560 522.950 16.620 ;
        RECT 469.130 16.420 522.950 16.560 ;
        RECT 522.630 16.360 522.950 16.420 ;
      LAYER via ;
        RECT 360.280 389.340 360.540 389.600 ;
        RECT 432.040 389.340 432.300 389.600 ;
        RECT 431.120 16.700 431.380 16.960 ;
        RECT 522.660 16.360 522.920 16.620 ;
      LAYER met2 ;
        RECT 360.170 400.180 360.450 404.000 ;
        RECT 360.170 400.000 360.480 400.180 ;
        RECT 360.340 389.630 360.480 400.000 ;
        RECT 360.280 389.310 360.540 389.630 ;
        RECT 432.040 389.310 432.300 389.630 ;
        RECT 432.100 324.370 432.240 389.310 ;
        RECT 431.180 324.230 432.240 324.370 ;
        RECT 431.180 16.990 431.320 324.230 ;
        RECT 431.120 16.670 431.380 16.990 ;
        RECT 522.660 16.330 522.920 16.650 ;
        RECT 522.720 2.400 522.860 16.330 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 388.520 366.090 388.580 ;
        RECT 404.410 388.520 404.730 388.580 ;
        RECT 365.770 388.380 404.730 388.520 ;
        RECT 365.770 388.320 366.090 388.380 ;
        RECT 404.410 388.320 404.730 388.380 ;
        RECT 404.870 19.960 405.190 20.020 ;
        RECT 540.570 19.960 540.890 20.020 ;
        RECT 404.870 19.820 540.890 19.960 ;
        RECT 404.870 19.760 405.190 19.820 ;
        RECT 540.570 19.760 540.890 19.820 ;
      LAYER via ;
        RECT 365.800 388.320 366.060 388.580 ;
        RECT 404.440 388.320 404.700 388.580 ;
        RECT 404.900 19.760 405.160 20.020 ;
        RECT 540.600 19.760 540.860 20.020 ;
      LAYER met2 ;
        RECT 365.690 400.180 365.970 404.000 ;
        RECT 365.690 400.000 366.000 400.180 ;
        RECT 365.860 388.610 366.000 400.000 ;
        RECT 365.800 388.290 366.060 388.610 ;
        RECT 404.440 388.290 404.700 388.610 ;
        RECT 404.500 324.370 404.640 388.290 ;
        RECT 403.580 324.230 404.640 324.370 ;
        RECT 403.580 82.870 403.720 324.230 ;
        RECT 403.580 82.730 405.100 82.870 ;
        RECT 404.960 20.050 405.100 82.730 ;
        RECT 404.900 19.730 405.160 20.050 ;
        RECT 540.600 19.730 540.860 20.050 ;
        RECT 540.660 2.400 540.800 19.730 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 370.830 392.600 371.150 392.660 ;
        RECT 466.510 392.600 466.830 392.660 ;
        RECT 370.830 392.460 466.830 392.600 ;
        RECT 370.830 392.400 371.150 392.460 ;
        RECT 466.510 392.400 466.830 392.460 ;
        RECT 465.590 20.640 465.910 20.700 ;
        RECT 558.050 20.640 558.370 20.700 ;
        RECT 465.590 20.500 558.370 20.640 ;
        RECT 465.590 20.440 465.910 20.500 ;
        RECT 558.050 20.440 558.370 20.500 ;
      LAYER via ;
        RECT 370.860 392.400 371.120 392.660 ;
        RECT 466.540 392.400 466.800 392.660 ;
        RECT 465.620 20.440 465.880 20.700 ;
        RECT 558.080 20.440 558.340 20.700 ;
      LAYER met2 ;
        RECT 370.750 400.180 371.030 404.000 ;
        RECT 370.750 400.000 371.060 400.180 ;
        RECT 370.920 392.690 371.060 400.000 ;
        RECT 370.860 392.370 371.120 392.690 ;
        RECT 466.540 392.370 466.800 392.690 ;
        RECT 466.600 324.370 466.740 392.370 ;
        RECT 465.680 324.230 466.740 324.370 ;
        RECT 465.680 20.730 465.820 324.230 ;
        RECT 465.620 20.410 465.880 20.730 ;
        RECT 558.080 20.410 558.340 20.730 ;
        RECT 558.140 2.400 558.280 20.410 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 373.130 17.580 373.450 17.640 ;
        RECT 575.990 17.580 576.310 17.640 ;
        RECT 373.130 17.440 576.310 17.580 ;
        RECT 373.130 17.380 373.450 17.440 ;
        RECT 575.990 17.380 576.310 17.440 ;
      LAYER via ;
        RECT 373.160 17.380 373.420 17.640 ;
        RECT 576.020 17.380 576.280 17.640 ;
      LAYER met2 ;
        RECT 376.270 400.250 376.550 404.000 ;
        RECT 375.060 400.110 376.550 400.250 ;
        RECT 375.060 324.370 375.200 400.110 ;
        RECT 376.270 400.000 376.550 400.110 ;
        RECT 373.220 324.230 375.200 324.370 ;
        RECT 373.220 17.670 373.360 324.230 ;
        RECT 373.160 17.350 373.420 17.670 ;
        RECT 576.020 17.350 576.280 17.670 ;
        RECT 576.080 2.400 576.220 17.350 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 85.170 19.620 85.490 19.680 ;
        RECT 221.330 19.620 221.650 19.680 ;
        RECT 85.170 19.480 221.650 19.620 ;
        RECT 85.170 19.420 85.490 19.480 ;
        RECT 221.330 19.420 221.650 19.480 ;
      LAYER via ;
        RECT 85.200 19.420 85.460 19.680 ;
        RECT 221.360 19.420 221.620 19.680 ;
      LAYER met2 ;
        RECT 225.850 400.250 226.130 404.000 ;
        RECT 224.640 400.110 226.130 400.250 ;
        RECT 224.640 390.730 224.780 400.110 ;
        RECT 225.850 400.000 226.130 400.110 ;
        RECT 221.420 390.590 224.780 390.730 ;
        RECT 221.420 19.710 221.560 390.590 ;
        RECT 85.200 19.390 85.460 19.710 ;
        RECT 221.360 19.390 221.620 19.710 ;
        RECT 85.260 2.400 85.400 19.390 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 381.870 392.940 382.190 393.000 ;
        RECT 444.890 392.940 445.210 393.000 ;
        RECT 381.870 392.800 445.210 392.940 ;
        RECT 381.870 392.740 382.190 392.800 ;
        RECT 444.890 392.740 445.210 392.800 ;
        RECT 444.890 387.500 445.210 387.560 ;
        RECT 444.890 387.360 448.570 387.500 ;
        RECT 444.890 387.300 445.210 387.360 ;
        RECT 448.430 386.820 448.570 387.360 ;
        RECT 479.390 386.820 479.710 386.880 ;
        RECT 448.430 386.680 479.710 386.820 ;
        RECT 479.390 386.620 479.710 386.680 ;
        RECT 479.390 20.300 479.710 20.360 ;
        RECT 499.630 20.300 499.950 20.360 ;
        RECT 479.390 20.160 499.950 20.300 ;
        RECT 479.390 20.100 479.710 20.160 ;
        RECT 499.630 20.100 499.950 20.160 ;
        RECT 499.630 16.900 499.950 16.960 ;
        RECT 593.930 16.900 594.250 16.960 ;
        RECT 499.630 16.760 594.250 16.900 ;
        RECT 499.630 16.700 499.950 16.760 ;
        RECT 593.930 16.700 594.250 16.760 ;
      LAYER via ;
        RECT 381.900 392.740 382.160 393.000 ;
        RECT 444.920 392.740 445.180 393.000 ;
        RECT 444.920 387.300 445.180 387.560 ;
        RECT 479.420 386.620 479.680 386.880 ;
        RECT 479.420 20.100 479.680 20.360 ;
        RECT 499.660 20.100 499.920 20.360 ;
        RECT 499.660 16.700 499.920 16.960 ;
        RECT 593.960 16.700 594.220 16.960 ;
      LAYER met2 ;
        RECT 381.790 400.180 382.070 404.000 ;
        RECT 381.790 400.000 382.100 400.180 ;
        RECT 381.960 393.030 382.100 400.000 ;
        RECT 381.900 392.710 382.160 393.030 ;
        RECT 444.920 392.710 445.180 393.030 ;
        RECT 444.980 387.590 445.120 392.710 ;
        RECT 444.920 387.270 445.180 387.590 ;
        RECT 479.420 386.590 479.680 386.910 ;
        RECT 479.480 20.390 479.620 386.590 ;
        RECT 479.420 20.070 479.680 20.390 ;
        RECT 499.660 20.070 499.920 20.390 ;
        RECT 499.720 16.990 499.860 20.070 ;
        RECT 499.660 16.670 499.920 16.990 ;
        RECT 593.960 16.670 594.220 16.990 ;
        RECT 594.020 2.400 594.160 16.670 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 427.960 387.700 468.120 387.840 ;
        RECT 387.390 387.500 387.710 387.560 ;
        RECT 427.960 387.500 428.100 387.700 ;
        RECT 387.390 387.360 428.100 387.500 ;
        RECT 467.980 387.500 468.120 387.700 ;
        RECT 486.290 387.500 486.610 387.560 ;
        RECT 467.980 387.360 486.610 387.500 ;
        RECT 387.390 387.300 387.710 387.360 ;
        RECT 486.290 387.300 486.610 387.360 ;
        RECT 486.290 14.520 486.610 14.580 ;
        RECT 611.410 14.520 611.730 14.580 ;
        RECT 486.290 14.380 611.730 14.520 ;
        RECT 486.290 14.320 486.610 14.380 ;
        RECT 611.410 14.320 611.730 14.380 ;
      LAYER via ;
        RECT 387.420 387.300 387.680 387.560 ;
        RECT 486.320 387.300 486.580 387.560 ;
        RECT 486.320 14.320 486.580 14.580 ;
        RECT 611.440 14.320 611.700 14.580 ;
      LAYER met2 ;
        RECT 387.310 400.180 387.590 404.000 ;
        RECT 387.310 400.000 387.620 400.180 ;
        RECT 387.480 387.590 387.620 400.000 ;
        RECT 387.420 387.270 387.680 387.590 ;
        RECT 486.320 387.270 486.580 387.590 ;
        RECT 486.380 14.610 486.520 387.270 ;
        RECT 486.320 14.290 486.580 14.610 ;
        RECT 611.440 14.290 611.700 14.610 ;
        RECT 611.500 2.400 611.640 14.290 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 109.090 16.900 109.410 16.960 ;
        RECT 229.150 16.900 229.470 16.960 ;
        RECT 109.090 16.760 229.470 16.900 ;
        RECT 109.090 16.700 109.410 16.760 ;
        RECT 229.150 16.700 229.470 16.760 ;
      LAYER via ;
        RECT 109.120 16.700 109.380 16.960 ;
        RECT 229.180 16.700 229.440 16.960 ;
      LAYER met2 ;
        RECT 233.210 400.250 233.490 404.000 ;
        RECT 232.000 400.110 233.490 400.250 ;
        RECT 232.000 324.370 232.140 400.110 ;
        RECT 233.210 400.000 233.490 400.110 ;
        RECT 229.240 324.230 232.140 324.370 ;
        RECT 229.240 16.990 229.380 324.230 ;
        RECT 109.120 16.670 109.380 16.990 ;
        RECT 229.180 16.670 229.440 16.990 ;
        RECT 109.180 2.400 109.320 16.670 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 132.550 24.040 132.870 24.100 ;
        RECT 235.590 24.040 235.910 24.100 ;
        RECT 132.550 23.900 235.910 24.040 ;
        RECT 132.550 23.840 132.870 23.900 ;
        RECT 235.590 23.840 235.910 23.900 ;
      LAYER via ;
        RECT 132.580 23.840 132.840 24.100 ;
        RECT 235.620 23.840 235.880 24.100 ;
      LAYER met2 ;
        RECT 240.110 400.250 240.390 404.000 ;
        RECT 238.900 400.110 240.390 400.250 ;
        RECT 238.900 386.650 239.040 400.110 ;
        RECT 240.110 400.000 240.390 400.110 ;
        RECT 235.680 386.510 239.040 386.650 ;
        RECT 235.680 24.130 235.820 386.510 ;
        RECT 132.580 23.810 132.840 24.130 ;
        RECT 235.620 23.810 235.880 24.130 ;
        RECT 132.640 2.400 132.780 23.810 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 150.490 24.380 150.810 24.440 ;
        RECT 242.490 24.380 242.810 24.440 ;
        RECT 150.490 24.240 242.810 24.380 ;
        RECT 150.490 24.180 150.810 24.240 ;
        RECT 242.490 24.180 242.810 24.240 ;
      LAYER via ;
        RECT 150.520 24.180 150.780 24.440 ;
        RECT 242.520 24.180 242.780 24.440 ;
      LAYER met2 ;
        RECT 245.630 400.250 245.910 404.000 ;
        RECT 244.420 400.110 245.910 400.250 ;
        RECT 244.420 384.610 244.560 400.110 ;
        RECT 245.630 400.000 245.910 400.110 ;
        RECT 242.580 384.470 244.560 384.610 ;
        RECT 242.580 24.470 242.720 384.470 ;
        RECT 150.520 24.150 150.780 24.470 ;
        RECT 242.520 24.150 242.780 24.470 ;
        RECT 150.580 2.400 150.720 24.150 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 167.970 24.720 168.290 24.780 ;
        RECT 249.850 24.720 250.170 24.780 ;
        RECT 167.970 24.580 250.170 24.720 ;
        RECT 167.970 24.520 168.290 24.580 ;
        RECT 249.850 24.520 250.170 24.580 ;
      LAYER via ;
        RECT 168.000 24.520 168.260 24.780 ;
        RECT 249.880 24.520 250.140 24.780 ;
      LAYER met2 ;
        RECT 251.150 400.250 251.430 404.000 ;
        RECT 249.940 400.110 251.430 400.250 ;
        RECT 249.940 24.810 250.080 400.110 ;
        RECT 251.150 400.000 251.430 400.110 ;
        RECT 168.000 24.490 168.260 24.810 ;
        RECT 249.880 24.490 250.140 24.810 ;
        RECT 168.060 2.400 168.200 24.490 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 179.470 393.280 179.790 393.340 ;
        RECT 256.750 393.280 257.070 393.340 ;
        RECT 179.470 393.140 257.070 393.280 ;
        RECT 179.470 393.080 179.790 393.140 ;
        RECT 256.750 393.080 257.070 393.140 ;
      LAYER via ;
        RECT 179.500 393.080 179.760 393.340 ;
        RECT 256.780 393.080 257.040 393.340 ;
      LAYER met2 ;
        RECT 256.670 400.180 256.950 404.000 ;
        RECT 256.670 400.000 256.980 400.180 ;
        RECT 256.840 393.370 256.980 400.000 ;
        RECT 179.500 393.050 179.760 393.370 ;
        RECT 256.780 393.050 257.040 393.370 ;
        RECT 179.560 82.870 179.700 393.050 ;
        RECT 179.560 82.730 183.840 82.870 ;
        RECT 183.700 1.770 183.840 82.730 ;
        RECT 185.790 1.770 186.350 2.400 ;
        RECT 183.700 1.630 186.350 1.770 ;
        RECT 185.790 -4.800 186.350 1.630 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 203.390 15.200 203.710 15.260 ;
        RECT 203.390 15.060 227.770 15.200 ;
        RECT 203.390 15.000 203.710 15.060 ;
        RECT 227.630 14.860 227.770 15.060 ;
        RECT 262.730 14.860 263.050 14.920 ;
        RECT 227.630 14.720 263.050 14.860 ;
        RECT 262.730 14.660 263.050 14.720 ;
      LAYER via ;
        RECT 203.420 15.000 203.680 15.260 ;
        RECT 262.760 14.660 263.020 14.920 ;
      LAYER met2 ;
        RECT 262.190 400.250 262.470 404.000 ;
        RECT 262.190 400.110 262.960 400.250 ;
        RECT 262.190 400.000 262.470 400.110 ;
        RECT 203.420 14.970 203.680 15.290 ;
        RECT 203.480 2.400 203.620 14.970 ;
        RECT 262.820 14.950 262.960 400.110 ;
        RECT 262.760 14.630 263.020 14.950 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 221.330 17.240 221.650 17.300 ;
        RECT 263.190 17.240 263.510 17.300 ;
        RECT 221.330 17.100 263.510 17.240 ;
        RECT 221.330 17.040 221.650 17.100 ;
        RECT 263.190 17.040 263.510 17.100 ;
      LAYER via ;
        RECT 221.360 17.040 221.620 17.300 ;
        RECT 263.220 17.040 263.480 17.300 ;
      LAYER met2 ;
        RECT 267.250 400.250 267.530 404.000 ;
        RECT 266.500 400.110 267.530 400.250 ;
        RECT 266.500 386.650 266.640 400.110 ;
        RECT 267.250 400.000 267.530 400.110 ;
        RECT 263.280 386.510 266.640 386.650 ;
        RECT 263.280 17.330 263.420 386.510 ;
        RECT 221.360 17.010 221.620 17.330 ;
        RECT 263.220 17.010 263.480 17.330 ;
        RECT 221.420 2.400 221.560 17.010 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.870 389.880 14.190 389.940 ;
        RECT 205.690 389.880 206.010 389.940 ;
        RECT 13.870 389.740 206.010 389.880 ;
        RECT 13.870 389.680 14.190 389.740 ;
        RECT 205.690 389.680 206.010 389.740 ;
      LAYER via ;
        RECT 13.900 389.680 14.160 389.940 ;
        RECT 205.720 389.680 205.980 389.940 ;
      LAYER met2 ;
        RECT 205.610 400.180 205.890 404.000 ;
        RECT 205.610 400.000 205.920 400.180 ;
        RECT 205.780 389.970 205.920 400.000 ;
        RECT 13.900 389.650 14.160 389.970 ;
        RECT 205.720 389.650 205.980 389.970 ;
        RECT 13.960 82.870 14.100 389.650 ;
        RECT 13.960 82.730 18.240 82.870 ;
        RECT 18.100 1.770 18.240 82.730 ;
        RECT 20.190 1.770 20.750 2.400 ;
        RECT 18.100 1.630 20.750 1.770 ;
        RECT 20.190 -4.800 20.750 1.630 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 207.990 386.480 208.310 386.540 ;
        RECT 211.670 386.480 211.990 386.540 ;
        RECT 207.990 386.340 211.990 386.480 ;
        RECT 207.990 386.280 208.310 386.340 ;
        RECT 211.670 386.280 211.990 386.340 ;
        RECT 43.770 18.260 44.090 18.320 ;
        RECT 207.990 18.260 208.310 18.320 ;
        RECT 43.770 18.120 208.310 18.260 ;
        RECT 43.770 18.060 44.090 18.120 ;
        RECT 207.990 18.060 208.310 18.120 ;
      LAYER via ;
        RECT 208.020 386.280 208.280 386.540 ;
        RECT 211.700 386.280 211.960 386.540 ;
        RECT 43.800 18.060 44.060 18.320 ;
        RECT 208.020 18.060 208.280 18.320 ;
      LAYER met2 ;
        RECT 212.970 400.250 213.250 404.000 ;
        RECT 211.760 400.110 213.250 400.250 ;
        RECT 211.760 386.570 211.900 400.110 ;
        RECT 212.970 400.000 213.250 400.110 ;
        RECT 208.020 386.250 208.280 386.570 ;
        RECT 211.700 386.250 211.960 386.570 ;
        RECT 208.080 18.350 208.220 386.250 ;
        RECT 43.800 18.030 44.060 18.350 ;
        RECT 208.020 18.030 208.280 18.350 ;
        RECT 43.860 2.400 44.000 18.030 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 258.590 387.160 258.910 387.220 ;
        RECT 274.690 387.160 275.010 387.220 ;
        RECT 258.590 387.020 275.010 387.160 ;
        RECT 258.590 386.960 258.910 387.020 ;
        RECT 274.690 386.960 275.010 387.020 ;
        RECT 244.790 17.580 245.110 17.640 ;
        RECT 258.590 17.580 258.910 17.640 ;
        RECT 244.790 17.440 258.910 17.580 ;
        RECT 244.790 17.380 245.110 17.440 ;
        RECT 258.590 17.380 258.910 17.440 ;
      LAYER via ;
        RECT 258.620 386.960 258.880 387.220 ;
        RECT 274.720 386.960 274.980 387.220 ;
        RECT 244.820 17.380 245.080 17.640 ;
        RECT 258.620 17.380 258.880 17.640 ;
      LAYER met2 ;
        RECT 274.610 400.180 274.890 404.000 ;
        RECT 274.610 400.000 274.920 400.180 ;
        RECT 274.780 387.250 274.920 400.000 ;
        RECT 258.620 386.930 258.880 387.250 ;
        RECT 274.720 386.930 274.980 387.250 ;
        RECT 258.680 17.670 258.820 386.930 ;
        RECT 244.820 17.350 245.080 17.670 ;
        RECT 258.620 17.350 258.880 17.670 ;
        RECT 244.880 2.400 245.020 17.350 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 266.870 389.880 267.190 389.940 ;
        RECT 280.210 389.880 280.530 389.940 ;
        RECT 266.870 389.740 280.530 389.880 ;
        RECT 266.870 389.680 267.190 389.740 ;
        RECT 280.210 389.680 280.530 389.740 ;
        RECT 266.870 386.480 267.190 386.540 ;
        RECT 264.200 386.340 267.190 386.480 ;
        RECT 264.200 386.200 264.340 386.340 ;
        RECT 266.870 386.280 267.190 386.340 ;
        RECT 264.110 385.940 264.430 386.200 ;
      LAYER via ;
        RECT 266.900 389.680 267.160 389.940 ;
        RECT 280.240 389.680 280.500 389.940 ;
        RECT 266.900 386.280 267.160 386.540 ;
        RECT 264.140 385.940 264.400 386.200 ;
      LAYER met2 ;
        RECT 280.130 400.180 280.410 404.000 ;
        RECT 280.130 400.000 280.440 400.180 ;
        RECT 280.300 389.970 280.440 400.000 ;
        RECT 266.900 389.650 267.160 389.970 ;
        RECT 280.240 389.650 280.500 389.970 ;
        RECT 266.960 386.570 267.100 389.650 ;
        RECT 266.900 386.250 267.160 386.570 ;
        RECT 264.140 385.910 264.400 386.230 ;
        RECT 262.610 1.770 263.170 2.400 ;
        RECT 264.200 1.770 264.340 385.910 ;
        RECT 262.610 1.630 264.340 1.770 ;
        RECT 262.610 -4.800 263.170 1.630 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 280.210 16.560 280.530 16.620 ;
        RECT 284.350 16.560 284.670 16.620 ;
        RECT 280.210 16.420 284.670 16.560 ;
        RECT 280.210 16.360 280.530 16.420 ;
        RECT 284.350 16.360 284.670 16.420 ;
      LAYER via ;
        RECT 280.240 16.360 280.500 16.620 ;
        RECT 284.380 16.360 284.640 16.620 ;
      LAYER met2 ;
        RECT 285.650 400.250 285.930 404.000 ;
        RECT 284.440 400.110 285.930 400.250 ;
        RECT 284.440 324.370 284.580 400.110 ;
        RECT 285.650 400.000 285.930 400.110 ;
        RECT 283.980 324.230 284.580 324.370 ;
        RECT 283.980 82.870 284.120 324.230 ;
        RECT 283.980 82.730 284.580 82.870 ;
        RECT 284.440 16.650 284.580 82.730 ;
        RECT 280.240 16.330 280.500 16.650 ;
        RECT 284.380 16.330 284.640 16.650 ;
        RECT 280.300 2.400 280.440 16.330 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 291.250 17.920 291.570 17.980 ;
        RECT 298.150 17.920 298.470 17.980 ;
        RECT 291.250 17.780 298.470 17.920 ;
        RECT 291.250 17.720 291.570 17.780 ;
        RECT 298.150 17.720 298.470 17.780 ;
      LAYER via ;
        RECT 291.280 17.720 291.540 17.980 ;
        RECT 298.180 17.720 298.440 17.980 ;
      LAYER met2 ;
        RECT 291.170 400.180 291.450 404.000 ;
        RECT 291.170 400.000 291.480 400.180 ;
        RECT 291.340 18.010 291.480 400.000 ;
        RECT 291.280 17.690 291.540 18.010 ;
        RECT 298.180 17.690 298.440 18.010 ;
        RECT 298.240 2.400 298.380 17.690 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 296.770 16.560 297.090 16.620 ;
        RECT 316.090 16.560 316.410 16.620 ;
        RECT 296.770 16.420 316.410 16.560 ;
        RECT 296.770 16.360 297.090 16.420 ;
        RECT 316.090 16.360 316.410 16.420 ;
      LAYER via ;
        RECT 296.800 16.360 297.060 16.620 ;
        RECT 316.120 16.360 316.380 16.620 ;
      LAYER met2 ;
        RECT 296.690 400.180 296.970 404.000 ;
        RECT 296.690 400.000 297.000 400.180 ;
        RECT 296.860 16.650 297.000 400.000 ;
        RECT 296.800 16.330 297.060 16.650 ;
        RECT 316.120 16.330 316.380 16.650 ;
        RECT 316.180 2.400 316.320 16.330 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 301.830 387.500 302.150 387.560 ;
        RECT 301.830 387.360 303.670 387.500 ;
        RECT 301.830 387.300 302.150 387.360 ;
        RECT 303.530 387.160 303.670 387.360 ;
        RECT 327.590 387.160 327.910 387.220 ;
        RECT 303.530 387.020 327.910 387.160 ;
        RECT 327.590 386.960 327.910 387.020 ;
        RECT 327.590 20.640 327.910 20.700 ;
        RECT 333.570 20.640 333.890 20.700 ;
        RECT 327.590 20.500 333.890 20.640 ;
        RECT 327.590 20.440 327.910 20.500 ;
        RECT 333.570 20.440 333.890 20.500 ;
      LAYER via ;
        RECT 301.860 387.300 302.120 387.560 ;
        RECT 327.620 386.960 327.880 387.220 ;
        RECT 327.620 20.440 327.880 20.700 ;
        RECT 333.600 20.440 333.860 20.700 ;
      LAYER met2 ;
        RECT 301.750 400.180 302.030 404.000 ;
        RECT 301.750 400.000 302.060 400.180 ;
        RECT 301.920 387.590 302.060 400.000 ;
        RECT 301.860 387.270 302.120 387.590 ;
        RECT 327.620 386.930 327.880 387.250 ;
        RECT 327.680 20.730 327.820 386.930 ;
        RECT 327.620 20.410 327.880 20.730 ;
        RECT 333.600 20.410 333.860 20.730 ;
        RECT 333.660 2.400 333.800 20.410 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.130 313.720 304.450 313.780 ;
        RECT 305.050 313.720 305.370 313.780 ;
        RECT 304.130 313.580 305.370 313.720 ;
        RECT 304.130 313.520 304.450 313.580 ;
        RECT 305.050 313.520 305.370 313.580 ;
        RECT 304.130 19.280 304.450 19.340 ;
        RECT 351.510 19.280 351.830 19.340 ;
        RECT 304.130 19.140 351.830 19.280 ;
        RECT 304.130 19.080 304.450 19.140 ;
        RECT 351.510 19.080 351.830 19.140 ;
      LAYER via ;
        RECT 304.160 313.520 304.420 313.780 ;
        RECT 305.080 313.520 305.340 313.780 ;
        RECT 304.160 19.080 304.420 19.340 ;
        RECT 351.540 19.080 351.800 19.340 ;
      LAYER met2 ;
        RECT 307.270 400.250 307.550 404.000 ;
        RECT 306.060 400.110 307.550 400.250 ;
        RECT 306.060 351.970 306.200 400.110 ;
        RECT 307.270 400.000 307.550 400.110 ;
        RECT 305.140 351.830 306.200 351.970 ;
        RECT 305.140 313.810 305.280 351.830 ;
        RECT 304.160 313.490 304.420 313.810 ;
        RECT 305.080 313.490 305.340 313.810 ;
        RECT 304.220 19.370 304.360 313.490 ;
        RECT 304.160 19.050 304.420 19.370 ;
        RECT 351.540 19.050 351.800 19.370 ;
        RECT 351.600 2.400 351.740 19.050 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 311.490 14.860 311.810 14.920 ;
        RECT 368.990 14.860 369.310 14.920 ;
        RECT 311.490 14.720 369.310 14.860 ;
        RECT 311.490 14.660 311.810 14.720 ;
        RECT 368.990 14.660 369.310 14.720 ;
      LAYER via ;
        RECT 311.520 14.660 311.780 14.920 ;
        RECT 369.020 14.660 369.280 14.920 ;
      LAYER met2 ;
        RECT 312.790 400.250 313.070 404.000 ;
        RECT 311.580 400.110 313.070 400.250 ;
        RECT 311.580 14.950 311.720 400.110 ;
        RECT 312.790 400.000 313.070 400.110 ;
        RECT 311.520 14.630 311.780 14.950 ;
        RECT 369.020 14.630 369.280 14.950 ;
        RECT 369.080 2.400 369.220 14.630 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 318.390 15.200 318.710 15.260 ;
        RECT 386.930 15.200 387.250 15.260 ;
        RECT 318.390 15.060 387.250 15.200 ;
        RECT 318.390 15.000 318.710 15.060 ;
        RECT 386.930 15.000 387.250 15.060 ;
      LAYER via ;
        RECT 318.420 15.000 318.680 15.260 ;
        RECT 386.960 15.000 387.220 15.260 ;
      LAYER met2 ;
        RECT 318.310 400.180 318.590 404.000 ;
        RECT 318.310 400.000 318.620 400.180 ;
        RECT 318.480 15.290 318.620 400.000 ;
        RECT 318.420 14.970 318.680 15.290 ;
        RECT 386.960 14.970 387.220 15.290 ;
        RECT 387.020 2.400 387.160 14.970 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.470 375.940 317.790 376.000 ;
        RECT 322.530 375.940 322.850 376.000 ;
        RECT 317.470 375.800 322.850 375.940 ;
        RECT 317.470 375.740 317.790 375.800 ;
        RECT 322.530 375.740 322.850 375.800 ;
        RECT 317.470 19.960 317.790 20.020 ;
        RECT 404.410 19.960 404.730 20.020 ;
        RECT 317.470 19.820 404.730 19.960 ;
        RECT 317.470 19.760 317.790 19.820 ;
        RECT 404.410 19.760 404.730 19.820 ;
      LAYER via ;
        RECT 317.500 375.740 317.760 376.000 ;
        RECT 322.560 375.740 322.820 376.000 ;
        RECT 317.500 19.760 317.760 20.020 ;
        RECT 404.440 19.760 404.700 20.020 ;
      LAYER met2 ;
        RECT 323.830 400.250 324.110 404.000 ;
        RECT 322.620 400.110 324.110 400.250 ;
        RECT 322.620 376.030 322.760 400.110 ;
        RECT 323.830 400.000 324.110 400.110 ;
        RECT 317.500 375.710 317.760 376.030 ;
        RECT 322.560 375.710 322.820 376.030 ;
        RECT 317.560 20.050 317.700 375.710 ;
        RECT 317.500 19.730 317.760 20.050 ;
        RECT 404.440 19.730 404.700 20.050 ;
        RECT 404.500 2.400 404.640 19.730 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.170 390.560 62.490 390.620 ;
        RECT 220.410 390.560 220.730 390.620 ;
        RECT 62.170 390.420 220.730 390.560 ;
        RECT 62.170 390.360 62.490 390.420 ;
        RECT 220.410 390.360 220.730 390.420 ;
      LAYER via ;
        RECT 62.200 390.360 62.460 390.620 ;
        RECT 220.440 390.360 220.700 390.620 ;
      LAYER met2 ;
        RECT 220.330 400.180 220.610 404.000 ;
        RECT 220.330 400.000 220.640 400.180 ;
        RECT 220.500 390.650 220.640 400.000 ;
        RECT 62.200 390.330 62.460 390.650 ;
        RECT 220.440 390.330 220.700 390.650 ;
        RECT 62.260 82.870 62.400 390.330 ;
        RECT 62.260 82.730 67.920 82.870 ;
        RECT 67.780 2.400 67.920 82.730 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.830 376.280 325.150 376.340 ;
        RECT 328.050 376.280 328.370 376.340 ;
        RECT 324.830 376.140 328.370 376.280 ;
        RECT 324.830 376.080 325.150 376.140 ;
        RECT 328.050 376.080 328.370 376.140 ;
        RECT 324.830 17.920 325.150 17.980 ;
        RECT 324.830 17.780 358.180 17.920 ;
        RECT 324.830 17.720 325.150 17.780 ;
        RECT 358.040 17.580 358.180 17.780 ;
        RECT 358.040 17.440 369.680 17.580 ;
        RECT 369.540 16.900 369.680 17.440 ;
        RECT 422.350 16.900 422.670 16.960 ;
        RECT 369.540 16.760 422.670 16.900 ;
        RECT 422.350 16.700 422.670 16.760 ;
      LAYER via ;
        RECT 324.860 376.080 325.120 376.340 ;
        RECT 328.080 376.080 328.340 376.340 ;
        RECT 324.860 17.720 325.120 17.980 ;
        RECT 422.380 16.700 422.640 16.960 ;
      LAYER met2 ;
        RECT 329.350 400.250 329.630 404.000 ;
        RECT 328.140 400.110 329.630 400.250 ;
        RECT 328.140 376.370 328.280 400.110 ;
        RECT 329.350 400.000 329.630 400.110 ;
        RECT 324.860 376.050 325.120 376.370 ;
        RECT 328.080 376.050 328.340 376.370 ;
        RECT 324.920 18.010 325.060 376.050 ;
        RECT 324.860 17.690 325.120 18.010 ;
        RECT 422.380 16.670 422.640 16.990 ;
        RECT 422.440 2.400 422.580 16.670 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 376.280 331.590 376.340 ;
        RECT 333.570 376.280 333.890 376.340 ;
        RECT 331.270 376.140 333.890 376.280 ;
        RECT 331.270 376.080 331.590 376.140 ;
        RECT 333.570 376.080 333.890 376.140 ;
        RECT 331.270 16.220 331.590 16.280 ;
        RECT 439.830 16.220 440.150 16.280 ;
        RECT 331.270 16.080 440.150 16.220 ;
        RECT 331.270 16.020 331.590 16.080 ;
        RECT 439.830 16.020 440.150 16.080 ;
      LAYER via ;
        RECT 331.300 376.080 331.560 376.340 ;
        RECT 333.600 376.080 333.860 376.340 ;
        RECT 331.300 16.020 331.560 16.280 ;
        RECT 439.860 16.020 440.120 16.280 ;
      LAYER met2 ;
        RECT 334.410 400.250 334.690 404.000 ;
        RECT 333.660 400.110 334.690 400.250 ;
        RECT 333.660 376.370 333.800 400.110 ;
        RECT 334.410 400.000 334.690 400.110 ;
        RECT 331.300 376.050 331.560 376.370 ;
        RECT 333.600 376.050 333.860 376.370 ;
        RECT 331.360 16.310 331.500 376.050 ;
        RECT 331.300 15.990 331.560 16.310 ;
        RECT 439.860 15.990 440.120 16.310 ;
        RECT 439.920 2.400 440.060 15.990 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 338.170 376.280 338.490 376.340 ;
        RECT 339.090 376.280 339.410 376.340 ;
        RECT 338.170 376.140 339.410 376.280 ;
        RECT 338.170 376.080 338.490 376.140 ;
        RECT 339.090 376.080 339.410 376.140 ;
        RECT 338.170 20.640 338.490 20.700 ;
        RECT 457.770 20.640 458.090 20.700 ;
        RECT 338.170 20.500 458.090 20.640 ;
        RECT 338.170 20.440 338.490 20.500 ;
        RECT 457.770 20.440 458.090 20.500 ;
      LAYER via ;
        RECT 338.200 376.080 338.460 376.340 ;
        RECT 339.120 376.080 339.380 376.340 ;
        RECT 338.200 20.440 338.460 20.700 ;
        RECT 457.800 20.440 458.060 20.700 ;
      LAYER met2 ;
        RECT 339.930 400.250 340.210 404.000 ;
        RECT 339.180 400.110 340.210 400.250 ;
        RECT 339.180 376.370 339.320 400.110 ;
        RECT 339.930 400.000 340.210 400.110 ;
        RECT 338.200 376.050 338.460 376.370 ;
        RECT 339.120 376.050 339.380 376.370 ;
        RECT 338.260 20.730 338.400 376.050 ;
        RECT 338.200 20.410 338.460 20.730 ;
        RECT 457.800 20.410 458.060 20.730 ;
        RECT 457.860 2.400 458.000 20.410 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.070 20.300 345.390 20.360 ;
        RECT 475.710 20.300 476.030 20.360 ;
        RECT 345.070 20.160 476.030 20.300 ;
        RECT 345.070 20.100 345.390 20.160 ;
        RECT 475.710 20.100 476.030 20.160 ;
      LAYER via ;
        RECT 345.100 20.100 345.360 20.360 ;
        RECT 475.740 20.100 476.000 20.360 ;
      LAYER met2 ;
        RECT 345.450 400.250 345.730 404.000 ;
        RECT 345.160 400.110 345.730 400.250 ;
        RECT 345.160 20.390 345.300 400.110 ;
        RECT 345.450 400.000 345.730 400.110 ;
        RECT 345.100 20.070 345.360 20.390 ;
        RECT 475.740 20.070 476.000 20.390 ;
        RECT 475.800 2.400 475.940 20.070 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.770 392.260 458.090 392.320 ;
        RECT 396.680 392.120 458.090 392.260 ;
        RECT 351.050 391.920 351.370 391.980 ;
        RECT 396.680 391.920 396.820 392.120 ;
        RECT 457.770 392.060 458.090 392.120 ;
        RECT 351.050 391.780 396.820 391.920 ;
        RECT 351.050 391.720 351.370 391.780 ;
        RECT 458.690 16.220 459.010 16.280 ;
        RECT 493.190 16.220 493.510 16.280 ;
        RECT 458.690 16.080 493.510 16.220 ;
        RECT 458.690 16.020 459.010 16.080 ;
        RECT 493.190 16.020 493.510 16.080 ;
      LAYER via ;
        RECT 351.080 391.720 351.340 391.980 ;
        RECT 457.800 392.060 458.060 392.320 ;
        RECT 458.720 16.020 458.980 16.280 ;
        RECT 493.220 16.020 493.480 16.280 ;
      LAYER met2 ;
        RECT 350.970 400.180 351.250 404.000 ;
        RECT 350.970 400.000 351.280 400.180 ;
        RECT 351.140 392.010 351.280 400.000 ;
        RECT 457.800 392.030 458.060 392.350 ;
        RECT 351.080 391.690 351.340 392.010 ;
        RECT 457.860 377.130 458.000 392.030 ;
        RECT 457.860 376.990 458.920 377.130 ;
        RECT 458.780 16.310 458.920 376.990 ;
        RECT 458.720 15.990 458.980 16.310 ;
        RECT 493.220 15.990 493.480 16.310 ;
        RECT 493.280 2.400 493.420 15.990 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.890 19.620 353.210 19.680 ;
        RECT 511.130 19.620 511.450 19.680 ;
        RECT 352.890 19.480 511.450 19.620 ;
        RECT 352.890 19.420 353.210 19.480 ;
        RECT 511.130 19.420 511.450 19.480 ;
      LAYER via ;
        RECT 352.920 19.420 353.180 19.680 ;
        RECT 511.160 19.420 511.420 19.680 ;
      LAYER met2 ;
        RECT 356.490 400.250 356.770 404.000 ;
        RECT 355.280 400.110 356.770 400.250 ;
        RECT 355.280 324.370 355.420 400.110 ;
        RECT 356.490 400.000 356.770 400.110 ;
        RECT 352.980 324.230 355.420 324.370 ;
        RECT 352.980 19.710 353.120 324.230 ;
        RECT 352.920 19.390 353.180 19.710 ;
        RECT 511.160 19.390 511.420 19.710 ;
        RECT 511.220 2.400 511.360 19.390 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 362.090 391.580 362.410 391.640 ;
        RECT 493.190 391.580 493.510 391.640 ;
        RECT 362.090 391.440 493.510 391.580 ;
        RECT 362.090 391.380 362.410 391.440 ;
        RECT 493.190 391.380 493.510 391.440 ;
        RECT 528.610 16.220 528.930 16.280 ;
        RECT 493.740 16.080 528.930 16.220 ;
        RECT 492.730 15.880 493.050 15.940 ;
        RECT 493.740 15.880 493.880 16.080 ;
        RECT 528.610 16.020 528.930 16.080 ;
        RECT 492.730 15.740 493.880 15.880 ;
        RECT 492.730 15.680 493.050 15.740 ;
      LAYER via ;
        RECT 362.120 391.380 362.380 391.640 ;
        RECT 493.220 391.380 493.480 391.640 ;
        RECT 492.760 15.680 493.020 15.940 ;
        RECT 528.640 16.020 528.900 16.280 ;
      LAYER met2 ;
        RECT 362.010 400.180 362.290 404.000 ;
        RECT 362.010 400.000 362.320 400.180 ;
        RECT 362.180 391.670 362.320 400.000 ;
        RECT 362.120 391.350 362.380 391.670 ;
        RECT 493.220 391.350 493.480 391.670 ;
        RECT 493.280 34.570 493.420 391.350 ;
        RECT 492.820 34.430 493.420 34.570 ;
        RECT 492.820 15.970 492.960 34.430 ;
        RECT 528.640 15.990 528.900 16.310 ;
        RECT 492.760 15.650 493.020 15.970 ;
        RECT 528.700 2.400 528.840 15.990 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 365.770 18.600 366.090 18.660 ;
        RECT 546.550 18.600 546.870 18.660 ;
        RECT 365.770 18.460 546.870 18.600 ;
        RECT 365.770 18.400 366.090 18.460 ;
        RECT 546.550 18.400 546.870 18.460 ;
      LAYER via ;
        RECT 365.800 18.400 366.060 18.660 ;
        RECT 546.580 18.400 546.840 18.660 ;
      LAYER met2 ;
        RECT 367.070 400.250 367.350 404.000 ;
        RECT 366.320 400.110 367.350 400.250 ;
        RECT 366.320 386.480 366.460 400.110 ;
        RECT 367.070 400.000 367.350 400.110 ;
        RECT 365.860 386.340 366.460 386.480 ;
        RECT 365.860 18.690 366.000 386.340 ;
        RECT 365.800 18.370 366.060 18.690 ;
        RECT 546.580 18.370 546.840 18.690 ;
        RECT 546.640 2.400 546.780 18.370 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 390.560 372.990 390.620 ;
        RECT 472.490 390.560 472.810 390.620 ;
        RECT 372.670 390.420 472.810 390.560 ;
        RECT 372.670 390.360 372.990 390.420 ;
        RECT 472.490 390.360 472.810 390.420 ;
        RECT 472.490 389.200 472.810 389.260 ;
        RECT 515.730 389.200 516.050 389.260 ;
        RECT 472.490 389.060 516.050 389.200 ;
        RECT 472.490 389.000 472.810 389.060 ;
        RECT 515.730 389.000 516.050 389.060 ;
        RECT 514.810 14.860 515.130 14.920 ;
        RECT 564.030 14.860 564.350 14.920 ;
        RECT 514.810 14.720 564.350 14.860 ;
        RECT 514.810 14.660 515.130 14.720 ;
        RECT 564.030 14.660 564.350 14.720 ;
      LAYER via ;
        RECT 372.700 390.360 372.960 390.620 ;
        RECT 472.520 390.360 472.780 390.620 ;
        RECT 472.520 389.000 472.780 389.260 ;
        RECT 515.760 389.000 516.020 389.260 ;
        RECT 514.840 14.660 515.100 14.920 ;
        RECT 564.060 14.660 564.320 14.920 ;
      LAYER met2 ;
        RECT 372.590 400.180 372.870 404.000 ;
        RECT 372.590 400.000 372.900 400.180 ;
        RECT 372.760 390.650 372.900 400.000 ;
        RECT 372.700 390.330 372.960 390.650 ;
        RECT 472.520 390.330 472.780 390.650 ;
        RECT 472.580 389.290 472.720 390.330 ;
        RECT 472.520 388.970 472.780 389.290 ;
        RECT 515.760 388.970 516.020 389.290 ;
        RECT 515.820 324.370 515.960 388.970 ;
        RECT 514.900 324.230 515.960 324.370 ;
        RECT 514.900 14.950 515.040 324.230 ;
        RECT 514.840 14.630 515.100 14.950 ;
        RECT 564.060 14.630 564.320 14.950 ;
        RECT 564.120 2.400 564.260 14.630 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 372.670 386.480 372.990 386.540 ;
        RECT 376.810 386.480 377.130 386.540 ;
        RECT 372.670 386.340 377.130 386.480 ;
        RECT 372.670 386.280 372.990 386.340 ;
        RECT 376.810 386.280 377.130 386.340 ;
        RECT 372.670 17.240 372.990 17.300 ;
        RECT 581.970 17.240 582.290 17.300 ;
        RECT 372.670 17.100 582.290 17.240 ;
        RECT 372.670 17.040 372.990 17.100 ;
        RECT 581.970 17.040 582.290 17.100 ;
      LAYER via ;
        RECT 372.700 386.280 372.960 386.540 ;
        RECT 376.840 386.280 377.100 386.540 ;
        RECT 372.700 17.040 372.960 17.300 ;
        RECT 582.000 17.040 582.260 17.300 ;
      LAYER met2 ;
        RECT 378.110 400.250 378.390 404.000 ;
        RECT 376.900 400.110 378.390 400.250 ;
        RECT 376.900 386.570 377.040 400.110 ;
        RECT 378.110 400.000 378.390 400.110 ;
        RECT 372.700 386.250 372.960 386.570 ;
        RECT 376.840 386.250 377.100 386.570 ;
        RECT 372.760 17.330 372.900 386.250 ;
        RECT 372.700 17.010 372.960 17.330 ;
        RECT 582.000 17.010 582.260 17.330 ;
        RECT 582.060 2.400 582.200 17.010 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 91.150 19.960 91.470 20.020 ;
        RECT 227.770 19.960 228.090 20.020 ;
        RECT 91.150 19.820 228.090 19.960 ;
        RECT 91.150 19.760 91.470 19.820 ;
        RECT 227.770 19.760 228.090 19.820 ;
      LAYER via ;
        RECT 91.180 19.760 91.440 20.020 ;
        RECT 227.800 19.760 228.060 20.020 ;
      LAYER met2 ;
        RECT 227.690 400.180 227.970 404.000 ;
        RECT 227.690 400.000 228.000 400.180 ;
        RECT 227.860 20.050 228.000 400.000 ;
        RECT 91.180 19.730 91.440 20.050 ;
        RECT 227.800 19.730 228.060 20.050 ;
        RECT 91.240 2.400 91.380 19.730 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 513.890 388.180 514.210 388.240 ;
        RECT 420.830 388.040 514.210 388.180 ;
        RECT 383.710 387.840 384.030 387.900 ;
        RECT 420.830 387.840 420.970 388.040 ;
        RECT 513.890 387.980 514.210 388.040 ;
        RECT 383.710 387.700 420.970 387.840 ;
        RECT 383.710 387.640 384.030 387.700 ;
        RECT 513.890 20.300 514.210 20.360 ;
        RECT 517.110 20.300 517.430 20.360 ;
        RECT 513.890 20.160 517.430 20.300 ;
        RECT 513.890 20.100 514.210 20.160 ;
        RECT 517.110 20.100 517.430 20.160 ;
        RECT 517.110 18.940 517.430 19.000 ;
        RECT 599.450 18.940 599.770 19.000 ;
        RECT 517.110 18.800 599.770 18.940 ;
        RECT 517.110 18.740 517.430 18.800 ;
        RECT 599.450 18.740 599.770 18.800 ;
      LAYER via ;
        RECT 383.740 387.640 384.000 387.900 ;
        RECT 513.920 387.980 514.180 388.240 ;
        RECT 513.920 20.100 514.180 20.360 ;
        RECT 517.140 20.100 517.400 20.360 ;
        RECT 517.140 18.740 517.400 19.000 ;
        RECT 599.480 18.740 599.740 19.000 ;
      LAYER met2 ;
        RECT 383.630 400.180 383.910 404.000 ;
        RECT 383.630 400.000 383.940 400.180 ;
        RECT 383.800 387.930 383.940 400.000 ;
        RECT 513.920 387.950 514.180 388.270 ;
        RECT 383.740 387.610 384.000 387.930 ;
        RECT 513.980 20.390 514.120 387.950 ;
        RECT 513.920 20.070 514.180 20.390 ;
        RECT 517.140 20.070 517.400 20.390 ;
        RECT 517.200 19.030 517.340 20.070 ;
        RECT 517.140 18.710 517.400 19.030 ;
        RECT 599.480 18.710 599.740 19.030 ;
        RECT 599.540 2.400 599.680 18.710 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 617.390 19.280 617.710 19.340 ;
        RECT 396.680 19.140 617.710 19.280 ;
        RECT 386.470 18.940 386.790 19.000 ;
        RECT 396.680 18.940 396.820 19.140 ;
        RECT 617.390 19.080 617.710 19.140 ;
        RECT 386.470 18.800 396.820 18.940 ;
        RECT 386.470 18.740 386.790 18.800 ;
      LAYER via ;
        RECT 386.500 18.740 386.760 19.000 ;
        RECT 617.420 19.080 617.680 19.340 ;
      LAYER met2 ;
        RECT 389.150 400.250 389.430 404.000 ;
        RECT 387.940 400.110 389.430 400.250 ;
        RECT 387.940 386.470 388.080 400.110 ;
        RECT 389.150 400.000 389.430 400.110 ;
        RECT 386.560 386.330 388.080 386.470 ;
        RECT 386.560 19.030 386.700 386.330 ;
        RECT 617.420 19.050 617.680 19.370 ;
        RECT 386.500 18.710 386.760 19.030 ;
        RECT 617.480 2.400 617.620 19.050 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 110.470 391.240 110.790 391.300 ;
        RECT 234.670 391.240 234.990 391.300 ;
        RECT 110.470 391.100 234.990 391.240 ;
        RECT 110.470 391.040 110.790 391.100 ;
        RECT 234.670 391.040 234.990 391.100 ;
      LAYER via ;
        RECT 110.500 391.040 110.760 391.300 ;
        RECT 234.700 391.040 234.960 391.300 ;
      LAYER met2 ;
        RECT 234.590 400.180 234.870 404.000 ;
        RECT 234.590 400.000 234.900 400.180 ;
        RECT 234.760 391.330 234.900 400.000 ;
        RECT 110.500 391.010 110.760 391.330 ;
        RECT 234.700 391.010 234.960 391.330 ;
        RECT 110.560 82.870 110.700 391.010 ;
        RECT 110.560 82.730 113.000 82.870 ;
        RECT 112.860 1.770 113.000 82.730 ;
        RECT 114.950 1.770 115.510 2.400 ;
        RECT 112.860 1.630 115.510 1.770 ;
        RECT 114.950 -4.800 115.510 1.630 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 241.570 372.880 241.890 372.940 ;
        RECT 242.950 372.880 243.270 372.940 ;
        RECT 241.570 372.740 243.270 372.880 ;
        RECT 241.570 372.680 241.890 372.740 ;
        RECT 242.950 372.680 243.270 372.740 ;
        RECT 138.530 16.220 138.850 16.280 ;
        RECT 138.530 16.080 233.060 16.220 ;
        RECT 138.530 16.020 138.850 16.080 ;
        RECT 232.920 15.880 233.060 16.080 ;
        RECT 242.950 15.880 243.270 15.940 ;
        RECT 232.920 15.740 243.270 15.880 ;
        RECT 242.950 15.680 243.270 15.740 ;
      LAYER via ;
        RECT 241.600 372.680 241.860 372.940 ;
        RECT 242.980 372.680 243.240 372.940 ;
        RECT 138.560 16.020 138.820 16.280 ;
        RECT 242.980 15.680 243.240 15.940 ;
      LAYER met2 ;
        RECT 241.950 400.250 242.230 404.000 ;
        RECT 241.660 400.110 242.230 400.250 ;
        RECT 241.660 372.970 241.800 400.110 ;
        RECT 241.950 400.000 242.230 400.110 ;
        RECT 241.600 372.650 241.860 372.970 ;
        RECT 242.980 372.650 243.240 372.970 ;
        RECT 138.560 15.990 138.820 16.310 ;
        RECT 138.620 2.400 138.760 15.990 ;
        RECT 243.040 15.970 243.180 372.650 ;
        RECT 242.980 15.650 243.240 15.970 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 151.870 392.940 152.190 393.000 ;
        RECT 247.550 392.940 247.870 393.000 ;
        RECT 151.870 392.800 247.870 392.940 ;
        RECT 151.870 392.740 152.190 392.800 ;
        RECT 247.550 392.740 247.870 392.800 ;
      LAYER via ;
        RECT 151.900 392.740 152.160 393.000 ;
        RECT 247.580 392.740 247.840 393.000 ;
      LAYER met2 ;
        RECT 247.470 400.180 247.750 404.000 ;
        RECT 247.470 400.000 247.780 400.180 ;
        RECT 247.640 393.030 247.780 400.000 ;
        RECT 151.900 392.710 152.160 393.030 ;
        RECT 247.580 392.710 247.840 393.030 ;
        RECT 151.960 82.870 152.100 392.710 ;
        RECT 151.960 82.730 154.400 82.870 ;
        RECT 154.260 1.770 154.400 82.730 ;
        RECT 156.350 1.770 156.910 2.400 ;
        RECT 154.260 1.630 156.910 1.770 ;
        RECT 156.350 -4.800 156.910 1.630 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.930 386.480 249.250 386.540 ;
        RECT 251.690 386.480 252.010 386.540 ;
        RECT 248.930 386.340 252.010 386.480 ;
        RECT 248.930 386.280 249.250 386.340 ;
        RECT 251.690 386.280 252.010 386.340 ;
        RECT 173.950 15.880 174.270 15.940 ;
        RECT 173.950 15.740 232.600 15.880 ;
        RECT 173.950 15.680 174.270 15.740 ;
        RECT 232.460 15.540 232.600 15.740 ;
        RECT 248.930 15.540 249.250 15.600 ;
        RECT 232.460 15.400 249.250 15.540 ;
        RECT 248.930 15.340 249.250 15.400 ;
      LAYER via ;
        RECT 248.960 386.280 249.220 386.540 ;
        RECT 251.720 386.280 251.980 386.540 ;
        RECT 173.980 15.680 174.240 15.940 ;
        RECT 248.960 15.340 249.220 15.600 ;
      LAYER met2 ;
        RECT 252.990 400.250 253.270 404.000 ;
        RECT 251.780 400.110 253.270 400.250 ;
        RECT 251.780 386.570 251.920 400.110 ;
        RECT 252.990 400.000 253.270 400.110 ;
        RECT 248.960 386.250 249.220 386.570 ;
        RECT 251.720 386.250 251.980 386.570 ;
        RECT 173.980 15.650 174.240 15.970 ;
        RECT 174.040 2.400 174.180 15.650 ;
        RECT 249.020 15.630 249.160 386.250 ;
        RECT 248.960 15.310 249.220 15.630 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 186.370 389.540 186.690 389.600 ;
        RECT 258.590 389.540 258.910 389.600 ;
        RECT 186.370 389.400 258.910 389.540 ;
        RECT 186.370 389.340 186.690 389.400 ;
        RECT 258.590 389.340 258.910 389.400 ;
      LAYER via ;
        RECT 186.400 389.340 186.660 389.600 ;
        RECT 258.620 389.340 258.880 389.600 ;
      LAYER met2 ;
        RECT 258.510 400.180 258.790 404.000 ;
        RECT 258.510 400.000 258.820 400.180 ;
        RECT 258.680 389.630 258.820 400.000 ;
        RECT 186.400 389.310 186.660 389.630 ;
        RECT 258.620 389.310 258.880 389.630 ;
        RECT 186.460 82.870 186.600 389.310 ;
        RECT 186.460 82.730 192.120 82.870 ;
        RECT 191.980 2.400 192.120 82.730 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 239.270 387.840 239.590 387.900 ;
        RECT 264.110 387.840 264.430 387.900 ;
        RECT 239.270 387.700 264.430 387.840 ;
        RECT 239.270 387.640 239.590 387.700 ;
        RECT 264.110 387.640 264.430 387.700 ;
        RECT 209.370 14.520 209.690 14.580 ;
        RECT 237.890 14.520 238.210 14.580 ;
        RECT 209.370 14.380 238.210 14.520 ;
        RECT 209.370 14.320 209.690 14.380 ;
        RECT 237.890 14.320 238.210 14.380 ;
      LAYER via ;
        RECT 239.300 387.640 239.560 387.900 ;
        RECT 264.140 387.640 264.400 387.900 ;
        RECT 209.400 14.320 209.660 14.580 ;
        RECT 237.920 14.320 238.180 14.580 ;
      LAYER met2 ;
        RECT 264.030 400.180 264.310 404.000 ;
        RECT 264.030 400.000 264.340 400.180 ;
        RECT 264.200 387.930 264.340 400.000 ;
        RECT 239.300 387.610 239.560 387.930 ;
        RECT 264.140 387.610 264.400 387.930 ;
        RECT 239.360 324.370 239.500 387.610 ;
        RECT 237.980 324.230 239.500 324.370 ;
        RECT 237.980 14.610 238.120 324.230 ;
        RECT 209.400 14.290 209.660 14.610 ;
        RECT 237.920 14.290 238.180 14.610 ;
        RECT 209.460 2.400 209.600 14.290 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 269.170 390.220 269.490 390.280 ;
        RECT 266.500 390.080 269.490 390.220 ;
        RECT 220.870 389.880 221.190 389.940 ;
        RECT 266.500 389.880 266.640 390.080 ;
        RECT 269.170 390.020 269.490 390.080 ;
        RECT 220.870 389.740 266.640 389.880 ;
        RECT 220.870 389.680 221.190 389.740 ;
      LAYER via ;
        RECT 220.900 389.680 221.160 389.940 ;
        RECT 269.200 390.020 269.460 390.280 ;
      LAYER met2 ;
        RECT 269.090 400.180 269.370 404.000 ;
        RECT 269.090 400.000 269.400 400.180 ;
        RECT 269.260 390.310 269.400 400.000 ;
        RECT 269.200 389.990 269.460 390.310 ;
        RECT 220.900 389.650 221.160 389.970 ;
        RECT 220.960 18.090 221.100 389.650 ;
        RECT 220.960 17.950 223.860 18.090 ;
        RECT 223.720 2.450 223.860 17.950 ;
        RECT 223.720 2.310 225.240 2.450 ;
        RECT 225.100 1.770 225.240 2.310 ;
        RECT 227.190 1.770 227.750 2.400 ;
        RECT 225.100 1.630 227.750 1.770 ;
        RECT 227.190 -4.800 227.750 1.630 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 49.750 18.600 50.070 18.660 ;
        RECT 214.430 18.600 214.750 18.660 ;
        RECT 49.750 18.460 214.750 18.600 ;
        RECT 49.750 18.400 50.070 18.460 ;
        RECT 214.430 18.400 214.750 18.460 ;
      LAYER via ;
        RECT 49.780 18.400 50.040 18.660 ;
        RECT 214.460 18.400 214.720 18.660 ;
      LAYER met2 ;
        RECT 214.810 400.250 215.090 404.000 ;
        RECT 214.520 400.110 215.090 400.250 ;
        RECT 214.520 18.690 214.660 400.110 ;
        RECT 214.810 400.000 215.090 400.110 ;
        RECT 49.780 18.370 50.040 18.690 ;
        RECT 214.460 18.370 214.720 18.690 ;
        RECT 49.840 2.400 49.980 18.370 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 248.470 391.580 248.790 391.640 ;
        RECT 276.530 391.580 276.850 391.640 ;
        RECT 248.470 391.440 276.850 391.580 ;
        RECT 248.470 391.380 248.790 391.440 ;
        RECT 276.530 391.380 276.850 391.440 ;
      LAYER via ;
        RECT 248.500 391.380 248.760 391.640 ;
        RECT 276.560 391.380 276.820 391.640 ;
      LAYER met2 ;
        RECT 276.450 400.180 276.730 404.000 ;
        RECT 276.450 400.000 276.760 400.180 ;
        RECT 276.620 391.670 276.760 400.000 ;
        RECT 248.500 391.350 248.760 391.670 ;
        RECT 276.560 391.350 276.820 391.670 ;
        RECT 248.560 14.690 248.700 391.350 ;
        RECT 248.560 14.550 251.000 14.690 ;
        RECT 250.860 2.400 251.000 14.550 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 272.390 389.540 272.710 389.600 ;
        RECT 282.050 389.540 282.370 389.600 ;
        RECT 272.390 389.400 282.370 389.540 ;
        RECT 272.390 389.340 272.710 389.400 ;
        RECT 282.050 389.340 282.370 389.400 ;
        RECT 268.710 16.560 269.030 16.620 ;
        RECT 272.390 16.560 272.710 16.620 ;
        RECT 268.710 16.420 272.710 16.560 ;
        RECT 268.710 16.360 269.030 16.420 ;
        RECT 272.390 16.360 272.710 16.420 ;
      LAYER via ;
        RECT 272.420 389.340 272.680 389.600 ;
        RECT 282.080 389.340 282.340 389.600 ;
        RECT 268.740 16.360 269.000 16.620 ;
        RECT 272.420 16.360 272.680 16.620 ;
      LAYER met2 ;
        RECT 281.970 400.180 282.250 404.000 ;
        RECT 281.970 400.000 282.280 400.180 ;
        RECT 282.140 389.630 282.280 400.000 ;
        RECT 272.420 389.310 272.680 389.630 ;
        RECT 282.080 389.310 282.340 389.630 ;
        RECT 272.480 16.650 272.620 389.310 ;
        RECT 268.740 16.330 269.000 16.650 ;
        RECT 272.420 16.330 272.680 16.650 ;
        RECT 268.800 2.400 268.940 16.330 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 282.970 386.480 283.290 386.540 ;
        RECT 286.190 386.480 286.510 386.540 ;
        RECT 282.970 386.340 286.510 386.480 ;
        RECT 282.970 386.280 283.290 386.340 ;
        RECT 286.190 386.280 286.510 386.340 ;
      LAYER via ;
        RECT 283.000 386.280 283.260 386.540 ;
        RECT 286.220 386.280 286.480 386.540 ;
      LAYER met2 ;
        RECT 287.490 400.250 287.770 404.000 ;
        RECT 286.280 400.110 287.770 400.250 ;
        RECT 286.280 386.570 286.420 400.110 ;
        RECT 287.490 400.000 287.770 400.110 ;
        RECT 283.000 386.250 283.260 386.570 ;
        RECT 286.220 386.250 286.480 386.570 ;
        RECT 283.060 1.770 283.200 386.250 ;
        RECT 286.070 1.770 286.630 2.400 ;
        RECT 283.060 1.630 286.630 1.770 ;
        RECT 286.070 -4.800 286.630 1.630 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 290.790 386.480 291.110 386.540 ;
        RECT 291.710 386.480 292.030 386.540 ;
        RECT 290.790 386.340 292.030 386.480 ;
        RECT 290.790 386.280 291.110 386.340 ;
        RECT 291.710 386.280 292.030 386.340 ;
        RECT 290.790 18.260 291.110 18.320 ;
        RECT 304.130 18.260 304.450 18.320 ;
        RECT 290.790 18.120 304.450 18.260 ;
        RECT 290.790 18.060 291.110 18.120 ;
        RECT 304.130 18.060 304.450 18.120 ;
      LAYER via ;
        RECT 290.820 386.280 291.080 386.540 ;
        RECT 291.740 386.280 292.000 386.540 ;
        RECT 290.820 18.060 291.080 18.320 ;
        RECT 304.160 18.060 304.420 18.320 ;
      LAYER met2 ;
        RECT 293.010 400.250 293.290 404.000 ;
        RECT 291.800 400.110 293.290 400.250 ;
        RECT 291.800 386.570 291.940 400.110 ;
        RECT 293.010 400.000 293.290 400.110 ;
        RECT 290.820 386.250 291.080 386.570 ;
        RECT 291.740 386.250 292.000 386.570 ;
        RECT 290.880 18.350 291.020 386.250 ;
        RECT 290.820 18.030 291.080 18.350 ;
        RECT 304.160 18.030 304.420 18.350 ;
        RECT 304.220 2.400 304.360 18.030 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 297.230 15.540 297.550 15.600 ;
        RECT 321.610 15.540 321.930 15.600 ;
        RECT 297.230 15.400 321.930 15.540 ;
        RECT 297.230 15.340 297.550 15.400 ;
        RECT 321.610 15.340 321.930 15.400 ;
      LAYER via ;
        RECT 297.260 15.340 297.520 15.600 ;
        RECT 321.640 15.340 321.900 15.600 ;
      LAYER met2 ;
        RECT 298.530 400.250 298.810 404.000 ;
        RECT 297.320 400.110 298.810 400.250 ;
        RECT 297.320 15.630 297.460 400.110 ;
        RECT 298.530 400.000 298.810 400.110 ;
        RECT 297.260 15.310 297.520 15.630 ;
        RECT 321.640 15.310 321.900 15.630 ;
        RECT 321.700 2.400 321.840 15.310 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 304.590 20.300 304.910 20.360 ;
        RECT 339.550 20.300 339.870 20.360 ;
        RECT 304.590 20.160 339.870 20.300 ;
        RECT 304.590 20.100 304.910 20.160 ;
        RECT 339.550 20.100 339.870 20.160 ;
      LAYER via ;
        RECT 304.620 20.100 304.880 20.360 ;
        RECT 339.580 20.100 339.840 20.360 ;
      LAYER met2 ;
        RECT 303.590 400.250 303.870 404.000 ;
        RECT 303.590 400.110 304.820 400.250 ;
        RECT 303.590 400.000 303.870 400.110 ;
        RECT 304.680 338.170 304.820 400.110 ;
        RECT 304.220 338.030 304.820 338.170 ;
        RECT 304.220 314.570 304.360 338.030 ;
        RECT 304.220 314.430 304.820 314.570 ;
        RECT 304.680 20.390 304.820 314.430 ;
        RECT 304.620 20.070 304.880 20.390 ;
        RECT 339.580 20.070 339.840 20.390 ;
        RECT 339.640 2.400 339.780 20.070 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 309.190 390.900 309.510 390.960 ;
        RECT 341.390 390.900 341.710 390.960 ;
        RECT 309.190 390.760 341.710 390.900 ;
        RECT 309.190 390.700 309.510 390.760 ;
        RECT 341.390 390.700 341.710 390.760 ;
        RECT 341.390 17.580 341.710 17.640 ;
        RECT 357.490 17.580 357.810 17.640 ;
        RECT 341.390 17.440 357.810 17.580 ;
        RECT 341.390 17.380 341.710 17.440 ;
        RECT 357.490 17.380 357.810 17.440 ;
      LAYER via ;
        RECT 309.220 390.700 309.480 390.960 ;
        RECT 341.420 390.700 341.680 390.960 ;
        RECT 341.420 17.380 341.680 17.640 ;
        RECT 357.520 17.380 357.780 17.640 ;
      LAYER met2 ;
        RECT 309.110 400.180 309.390 404.000 ;
        RECT 309.110 400.000 309.420 400.180 ;
        RECT 309.280 390.990 309.420 400.000 ;
        RECT 309.220 390.670 309.480 390.990 ;
        RECT 341.420 390.670 341.680 390.990 ;
        RECT 341.480 17.670 341.620 390.670 ;
        RECT 341.420 17.350 341.680 17.670 ;
        RECT 357.520 17.350 357.780 17.670 ;
        RECT 357.580 2.400 357.720 17.350 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.570 387.500 310.890 387.560 ;
        RECT 313.330 387.500 313.650 387.560 ;
        RECT 310.570 387.360 313.650 387.500 ;
        RECT 310.570 387.300 310.890 387.360 ;
        RECT 313.330 387.300 313.650 387.360 ;
        RECT 310.570 18.940 310.890 19.000 ;
        RECT 374.970 18.940 375.290 19.000 ;
        RECT 310.570 18.800 375.290 18.940 ;
        RECT 310.570 18.740 310.890 18.800 ;
        RECT 374.970 18.740 375.290 18.800 ;
      LAYER via ;
        RECT 310.600 387.300 310.860 387.560 ;
        RECT 313.360 387.300 313.620 387.560 ;
        RECT 310.600 18.740 310.860 19.000 ;
        RECT 375.000 18.740 375.260 19.000 ;
      LAYER met2 ;
        RECT 314.630 400.250 314.910 404.000 ;
        RECT 313.420 400.110 314.910 400.250 ;
        RECT 313.420 387.590 313.560 400.110 ;
        RECT 314.630 400.000 314.910 400.110 ;
        RECT 310.600 387.270 310.860 387.590 ;
        RECT 313.360 387.270 313.620 387.590 ;
        RECT 310.660 19.030 310.800 387.270 ;
        RECT 310.600 18.710 310.860 19.030 ;
        RECT 375.000 18.710 375.260 19.030 ;
        RECT 375.060 2.400 375.200 18.710 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 317.930 376.280 318.250 376.340 ;
        RECT 318.850 376.280 319.170 376.340 ;
        RECT 317.930 376.140 319.170 376.280 ;
        RECT 317.930 376.080 318.250 376.140 ;
        RECT 318.850 376.080 319.170 376.140 ;
        RECT 317.930 15.880 318.250 15.940 ;
        RECT 392.910 15.880 393.230 15.940 ;
        RECT 317.930 15.740 393.230 15.880 ;
        RECT 317.930 15.680 318.250 15.740 ;
        RECT 392.910 15.680 393.230 15.740 ;
      LAYER via ;
        RECT 317.960 376.080 318.220 376.340 ;
        RECT 318.880 376.080 319.140 376.340 ;
        RECT 317.960 15.680 318.220 15.940 ;
        RECT 392.940 15.680 393.200 15.940 ;
      LAYER met2 ;
        RECT 320.150 400.250 320.430 404.000 ;
        RECT 318.940 400.110 320.430 400.250 ;
        RECT 318.940 376.370 319.080 400.110 ;
        RECT 320.150 400.000 320.430 400.110 ;
        RECT 317.960 376.050 318.220 376.370 ;
        RECT 318.880 376.050 319.140 376.370 ;
        RECT 318.020 15.970 318.160 376.050 ;
        RECT 317.960 15.650 318.220 15.970 ;
        RECT 392.940 15.650 393.200 15.970 ;
        RECT 393.000 2.400 393.140 15.650 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 324.370 16.560 324.690 16.620 ;
        RECT 410.390 16.560 410.710 16.620 ;
        RECT 324.370 16.420 410.710 16.560 ;
        RECT 324.370 16.360 324.690 16.420 ;
        RECT 410.390 16.360 410.710 16.420 ;
      LAYER via ;
        RECT 324.400 16.360 324.660 16.620 ;
        RECT 410.420 16.360 410.680 16.620 ;
      LAYER met2 ;
        RECT 325.670 400.250 325.950 404.000 ;
        RECT 324.460 400.110 325.950 400.250 ;
        RECT 324.460 16.650 324.600 400.110 ;
        RECT 325.670 400.000 325.950 400.110 ;
        RECT 324.400 16.330 324.660 16.650 ;
        RECT 410.420 16.330 410.680 16.650 ;
        RECT 410.480 2.400 410.620 16.330 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 69.070 390.900 69.390 390.960 ;
        RECT 220.870 390.900 221.190 390.960 ;
        RECT 69.070 390.760 221.190 390.900 ;
        RECT 69.070 390.700 69.390 390.760 ;
        RECT 220.870 390.700 221.190 390.760 ;
      LAYER via ;
        RECT 69.100 390.700 69.360 390.960 ;
        RECT 220.900 390.700 221.160 390.960 ;
      LAYER met2 ;
        RECT 222.170 400.250 222.450 404.000 ;
        RECT 220.960 400.110 222.450 400.250 ;
        RECT 220.960 390.990 221.100 400.110 ;
        RECT 222.170 400.000 222.450 400.110 ;
        RECT 69.100 390.670 69.360 390.990 ;
        RECT 220.900 390.670 221.160 390.990 ;
        RECT 69.160 82.870 69.300 390.670 ;
        RECT 69.160 82.730 71.600 82.870 ;
        RECT 71.460 1.770 71.600 82.730 ;
        RECT 73.550 1.770 74.110 2.400 ;
        RECT 71.460 1.630 74.110 1.770 ;
        RECT 73.550 -4.800 74.110 1.630 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 331.270 393.280 331.590 393.340 ;
        RECT 417.290 393.280 417.610 393.340 ;
        RECT 331.270 393.140 417.610 393.280 ;
        RECT 331.270 393.080 331.590 393.140 ;
        RECT 417.290 393.080 417.610 393.140 ;
        RECT 417.290 15.880 417.610 15.940 ;
        RECT 428.330 15.880 428.650 15.940 ;
        RECT 417.290 15.740 428.650 15.880 ;
        RECT 417.290 15.680 417.610 15.740 ;
        RECT 428.330 15.680 428.650 15.740 ;
      LAYER via ;
        RECT 331.300 393.080 331.560 393.340 ;
        RECT 417.320 393.080 417.580 393.340 ;
        RECT 417.320 15.680 417.580 15.940 ;
        RECT 428.360 15.680 428.620 15.940 ;
      LAYER met2 ;
        RECT 331.190 400.180 331.470 404.000 ;
        RECT 331.190 400.000 331.500 400.180 ;
        RECT 331.360 393.370 331.500 400.000 ;
        RECT 331.300 393.050 331.560 393.370 ;
        RECT 417.320 393.050 417.580 393.370 ;
        RECT 417.380 15.970 417.520 393.050 ;
        RECT 417.320 15.650 417.580 15.970 ;
        RECT 428.360 15.650 428.620 15.970 ;
        RECT 428.420 2.400 428.560 15.650 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 336.330 388.860 336.650 388.920 ;
        RECT 389.690 388.860 390.010 388.920 ;
        RECT 336.330 388.720 390.010 388.860 ;
        RECT 336.330 388.660 336.650 388.720 ;
        RECT 389.690 388.660 390.010 388.720 ;
        RECT 389.690 15.200 390.010 15.260 ;
        RECT 445.810 15.200 446.130 15.260 ;
        RECT 389.690 15.060 446.130 15.200 ;
        RECT 389.690 15.000 390.010 15.060 ;
        RECT 445.810 15.000 446.130 15.060 ;
      LAYER via ;
        RECT 336.360 388.660 336.620 388.920 ;
        RECT 389.720 388.660 389.980 388.920 ;
        RECT 389.720 15.000 389.980 15.260 ;
        RECT 445.840 15.000 446.100 15.260 ;
      LAYER met2 ;
        RECT 336.250 400.180 336.530 404.000 ;
        RECT 336.250 400.000 336.560 400.180 ;
        RECT 336.420 388.950 336.560 400.000 ;
        RECT 336.360 388.630 336.620 388.950 ;
        RECT 389.720 388.630 389.980 388.950 ;
        RECT 389.780 15.290 389.920 388.630 ;
        RECT 389.720 14.970 389.980 15.290 ;
        RECT 445.840 14.970 446.100 15.290 ;
        RECT 445.900 2.400 446.040 14.970 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 397.510 391.920 397.830 391.980 ;
        RECT 459.150 391.920 459.470 391.980 ;
        RECT 397.510 391.780 459.470 391.920 ;
        RECT 397.510 391.720 397.830 391.780 ;
        RECT 459.150 391.720 459.470 391.780 ;
        RECT 341.850 389.200 342.170 389.260 ;
        RECT 397.510 389.200 397.830 389.260 ;
        RECT 341.850 389.060 397.830 389.200 ;
        RECT 341.850 389.000 342.170 389.060 ;
        RECT 397.510 389.000 397.830 389.060 ;
        RECT 459.150 16.560 459.470 16.620 ;
        RECT 463.750 16.560 464.070 16.620 ;
        RECT 459.150 16.420 464.070 16.560 ;
        RECT 459.150 16.360 459.470 16.420 ;
        RECT 463.750 16.360 464.070 16.420 ;
      LAYER via ;
        RECT 397.540 391.720 397.800 391.980 ;
        RECT 459.180 391.720 459.440 391.980 ;
        RECT 341.880 389.000 342.140 389.260 ;
        RECT 397.540 389.000 397.800 389.260 ;
        RECT 459.180 16.360 459.440 16.620 ;
        RECT 463.780 16.360 464.040 16.620 ;
      LAYER met2 ;
        RECT 341.770 400.180 342.050 404.000 ;
        RECT 341.770 400.000 342.080 400.180 ;
        RECT 341.940 389.290 342.080 400.000 ;
        RECT 397.540 391.690 397.800 392.010 ;
        RECT 459.180 391.690 459.440 392.010 ;
        RECT 397.600 389.290 397.740 391.690 ;
        RECT 341.880 388.970 342.140 389.290 ;
        RECT 397.540 388.970 397.800 389.290 ;
        RECT 459.240 16.650 459.380 391.690 ;
        RECT 459.180 16.330 459.440 16.650 ;
        RECT 463.780 16.330 464.040 16.650 ;
        RECT 463.840 2.400 463.980 16.330 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 345.530 24.040 345.850 24.100 ;
        RECT 481.230 24.040 481.550 24.100 ;
        RECT 345.530 23.900 481.550 24.040 ;
        RECT 345.530 23.840 345.850 23.900 ;
        RECT 481.230 23.840 481.550 23.900 ;
      LAYER via ;
        RECT 345.560 23.840 345.820 24.100 ;
        RECT 481.260 23.840 481.520 24.100 ;
      LAYER met2 ;
        RECT 347.290 400.250 347.570 404.000 ;
        RECT 346.080 400.110 347.570 400.250 ;
        RECT 346.080 303.670 346.220 400.110 ;
        RECT 347.290 400.000 347.570 400.110 ;
        RECT 345.620 303.530 346.220 303.670 ;
        RECT 345.620 24.130 345.760 303.530 ;
        RECT 345.560 23.810 345.820 24.130 ;
        RECT 481.260 23.810 481.520 24.130 ;
        RECT 481.320 2.400 481.460 23.810 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 352.890 390.900 353.210 390.960 ;
        RECT 493.650 390.900 493.970 390.960 ;
        RECT 352.890 390.760 493.970 390.900 ;
        RECT 352.890 390.700 353.210 390.760 ;
        RECT 493.650 390.700 493.970 390.760 ;
        RECT 493.650 16.900 493.970 16.960 ;
        RECT 499.170 16.900 499.490 16.960 ;
        RECT 493.650 16.760 499.490 16.900 ;
        RECT 493.650 16.700 493.970 16.760 ;
        RECT 499.170 16.700 499.490 16.760 ;
      LAYER via ;
        RECT 352.920 390.700 353.180 390.960 ;
        RECT 493.680 390.700 493.940 390.960 ;
        RECT 493.680 16.700 493.940 16.960 ;
        RECT 499.200 16.700 499.460 16.960 ;
      LAYER met2 ;
        RECT 352.810 400.180 353.090 404.000 ;
        RECT 352.810 400.000 353.120 400.180 ;
        RECT 352.980 390.990 353.120 400.000 ;
        RECT 352.920 390.670 353.180 390.990 ;
        RECT 493.680 390.670 493.940 390.990 ;
        RECT 493.740 16.990 493.880 390.670 ;
        RECT 493.680 16.670 493.940 16.990 ;
        RECT 499.200 16.670 499.460 16.990 ;
        RECT 499.260 2.400 499.400 16.670 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 351.970 386.480 352.290 386.540 ;
        RECT 357.030 386.480 357.350 386.540 ;
        RECT 351.970 386.340 357.350 386.480 ;
        RECT 351.970 386.280 352.290 386.340 ;
        RECT 357.030 386.280 357.350 386.340 ;
        RECT 351.970 19.280 352.290 19.340 ;
        RECT 396.130 19.280 396.450 19.340 ;
        RECT 351.970 19.140 396.450 19.280 ;
        RECT 351.970 19.080 352.290 19.140 ;
        RECT 396.130 19.080 396.450 19.140 ;
        RECT 397.050 18.940 397.370 19.000 ;
        RECT 516.650 18.940 516.970 19.000 ;
        RECT 397.050 18.800 516.970 18.940 ;
        RECT 397.050 18.740 397.370 18.800 ;
        RECT 516.650 18.740 516.970 18.800 ;
      LAYER via ;
        RECT 352.000 386.280 352.260 386.540 ;
        RECT 357.060 386.280 357.320 386.540 ;
        RECT 352.000 19.080 352.260 19.340 ;
        RECT 396.160 19.080 396.420 19.340 ;
        RECT 397.080 18.740 397.340 19.000 ;
        RECT 516.680 18.740 516.940 19.000 ;
      LAYER met2 ;
        RECT 358.330 400.250 358.610 404.000 ;
        RECT 357.120 400.110 358.610 400.250 ;
        RECT 357.120 386.570 357.260 400.110 ;
        RECT 358.330 400.000 358.610 400.110 ;
        RECT 352.000 386.250 352.260 386.570 ;
        RECT 357.060 386.250 357.320 386.570 ;
        RECT 352.060 19.370 352.200 386.250 ;
        RECT 352.000 19.050 352.260 19.370 ;
        RECT 396.160 19.050 396.420 19.370 ;
        RECT 396.220 18.770 396.360 19.050 ;
        RECT 397.080 18.770 397.340 19.030 ;
        RECT 396.220 18.710 397.340 18.770 ;
        RECT 516.680 18.710 516.940 19.030 ;
        RECT 396.220 18.630 397.280 18.710 ;
        RECT 516.740 2.400 516.880 18.710 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 363.930 389.880 364.250 389.940 ;
        RECT 515.270 389.880 515.590 389.940 ;
        RECT 363.930 389.740 515.590 389.880 ;
        RECT 363.930 389.680 364.250 389.740 ;
        RECT 515.270 389.680 515.590 389.740 ;
        RECT 514.350 15.880 514.670 15.940 ;
        RECT 534.590 15.880 534.910 15.940 ;
        RECT 514.350 15.740 534.910 15.880 ;
        RECT 514.350 15.680 514.670 15.740 ;
        RECT 534.590 15.680 534.910 15.740 ;
      LAYER via ;
        RECT 363.960 389.680 364.220 389.940 ;
        RECT 515.300 389.680 515.560 389.940 ;
        RECT 514.380 15.680 514.640 15.940 ;
        RECT 534.620 15.680 534.880 15.940 ;
      LAYER met2 ;
        RECT 363.850 400.180 364.130 404.000 ;
        RECT 363.850 400.000 364.160 400.180 ;
        RECT 364.020 389.970 364.160 400.000 ;
        RECT 363.960 389.650 364.220 389.970 ;
        RECT 515.300 389.650 515.560 389.970 ;
        RECT 515.360 385.290 515.500 389.650 ;
        RECT 514.440 385.150 515.500 385.290 ;
        RECT 514.440 15.970 514.580 385.150 ;
        RECT 514.380 15.650 514.640 15.970 ;
        RECT 534.620 15.650 534.880 15.970 ;
        RECT 534.680 2.400 534.820 15.650 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 366.230 17.920 366.550 17.980 ;
        RECT 552.530 17.920 552.850 17.980 ;
        RECT 366.230 17.780 552.850 17.920 ;
        RECT 366.230 17.720 366.550 17.780 ;
        RECT 552.530 17.720 552.850 17.780 ;
      LAYER via ;
        RECT 366.260 17.720 366.520 17.980 ;
        RECT 552.560 17.720 552.820 17.980 ;
      LAYER met2 ;
        RECT 368.910 400.250 369.190 404.000 ;
        RECT 367.700 400.110 369.190 400.250 ;
        RECT 367.700 324.370 367.840 400.110 ;
        RECT 368.910 400.000 369.190 400.110 ;
        RECT 366.320 324.230 367.840 324.370 ;
        RECT 366.320 18.010 366.460 324.230 ;
        RECT 366.260 17.690 366.520 18.010 ;
        RECT 552.560 17.690 552.820 18.010 ;
        RECT 552.620 2.400 552.760 17.690 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 374.510 390.220 374.830 390.280 ;
        RECT 472.030 390.220 472.350 390.280 ;
        RECT 374.510 390.080 472.350 390.220 ;
        RECT 374.510 390.020 374.830 390.080 ;
        RECT 472.030 390.020 472.350 390.080 ;
        RECT 472.030 387.840 472.350 387.900 ;
        RECT 520.790 387.840 521.110 387.900 ;
        RECT 472.030 387.700 521.110 387.840 ;
        RECT 472.030 387.640 472.350 387.700 ;
        RECT 520.790 387.640 521.110 387.700 ;
        RECT 520.790 15.200 521.110 15.260 ;
        RECT 570.010 15.200 570.330 15.260 ;
        RECT 520.790 15.060 570.330 15.200 ;
        RECT 520.790 15.000 521.110 15.060 ;
        RECT 570.010 15.000 570.330 15.060 ;
      LAYER via ;
        RECT 374.540 390.020 374.800 390.280 ;
        RECT 472.060 390.020 472.320 390.280 ;
        RECT 472.060 387.640 472.320 387.900 ;
        RECT 520.820 387.640 521.080 387.900 ;
        RECT 520.820 15.000 521.080 15.260 ;
        RECT 570.040 15.000 570.300 15.260 ;
      LAYER met2 ;
        RECT 374.430 400.180 374.710 404.000 ;
        RECT 374.430 400.000 374.740 400.180 ;
        RECT 374.600 390.310 374.740 400.000 ;
        RECT 374.540 389.990 374.800 390.310 ;
        RECT 472.060 389.990 472.320 390.310 ;
        RECT 472.120 387.930 472.260 389.990 ;
        RECT 472.060 387.610 472.320 387.930 ;
        RECT 520.820 387.610 521.080 387.930 ;
        RECT 520.880 15.290 521.020 387.610 ;
        RECT 520.820 14.970 521.080 15.290 ;
        RECT 570.040 14.970 570.300 15.290 ;
        RECT 570.100 2.400 570.240 14.970 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 380.030 22.680 380.350 22.740 ;
        RECT 523.090 22.680 523.410 22.740 ;
        RECT 380.030 22.540 523.410 22.680 ;
        RECT 380.030 22.480 380.350 22.540 ;
        RECT 523.090 22.480 523.410 22.540 ;
        RECT 523.090 19.620 523.410 19.680 ;
        RECT 587.950 19.620 588.270 19.680 ;
        RECT 523.090 19.480 588.270 19.620 ;
        RECT 523.090 19.420 523.410 19.480 ;
        RECT 587.950 19.420 588.270 19.480 ;
      LAYER via ;
        RECT 380.060 22.480 380.320 22.740 ;
        RECT 523.120 22.480 523.380 22.740 ;
        RECT 523.120 19.420 523.380 19.680 ;
        RECT 587.980 19.420 588.240 19.680 ;
      LAYER met2 ;
        RECT 379.950 400.180 380.230 404.000 ;
        RECT 379.950 400.000 380.260 400.180 ;
        RECT 380.120 22.770 380.260 400.000 ;
        RECT 380.060 22.450 380.320 22.770 ;
        RECT 523.120 22.450 523.380 22.770 ;
        RECT 523.180 19.710 523.320 22.450 ;
        RECT 523.120 19.390 523.380 19.710 ;
        RECT 587.980 19.390 588.240 19.710 ;
        RECT 588.040 2.400 588.180 19.390 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 97.130 20.300 97.450 20.360 ;
        RECT 228.690 20.300 229.010 20.360 ;
        RECT 97.130 20.160 229.010 20.300 ;
        RECT 97.130 20.100 97.450 20.160 ;
        RECT 228.690 20.100 229.010 20.160 ;
      LAYER via ;
        RECT 97.160 20.100 97.420 20.360 ;
        RECT 228.720 20.100 228.980 20.360 ;
      LAYER met2 ;
        RECT 229.530 400.250 229.810 404.000 ;
        RECT 228.780 400.110 229.810 400.250 ;
        RECT 228.780 20.390 228.920 400.110 ;
        RECT 229.530 400.000 229.810 400.110 ;
        RECT 97.160 20.070 97.420 20.390 ;
        RECT 228.720 20.070 228.980 20.390 ;
        RECT 97.220 2.400 97.360 20.070 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 527.690 15.540 528.010 15.600 ;
        RECT 605.430 15.540 605.750 15.600 ;
        RECT 527.690 15.400 605.750 15.540 ;
        RECT 527.690 15.340 528.010 15.400 ;
        RECT 605.430 15.340 605.750 15.400 ;
      LAYER via ;
        RECT 527.720 15.340 527.980 15.600 ;
        RECT 605.460 15.340 605.720 15.600 ;
      LAYER met2 ;
        RECT 385.470 400.180 385.750 404.000 ;
        RECT 385.470 400.000 385.780 400.180 ;
        RECT 385.640 390.165 385.780 400.000 ;
        RECT 385.570 389.795 385.850 390.165 ;
        RECT 527.710 389.795 527.990 390.165 ;
        RECT 527.780 15.630 527.920 389.795 ;
        RECT 527.720 15.310 527.980 15.630 ;
        RECT 605.460 15.310 605.720 15.630 ;
        RECT 605.520 2.400 605.660 15.310 ;
        RECT 605.310 -4.800 605.870 2.400 ;
      LAYER via2 ;
        RECT 385.570 389.840 385.850 390.120 ;
        RECT 527.710 389.840 527.990 390.120 ;
      LAYER met3 ;
        RECT 385.545 390.130 385.875 390.145 ;
        RECT 527.685 390.130 528.015 390.145 ;
        RECT 385.545 389.830 528.015 390.130 ;
        RECT 385.545 389.815 385.875 389.830 ;
        RECT 527.685 389.815 528.015 389.830 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 535.050 15.880 535.370 15.940 ;
        RECT 623.370 15.880 623.690 15.940 ;
        RECT 535.050 15.740 623.690 15.880 ;
        RECT 535.050 15.680 535.370 15.740 ;
        RECT 623.370 15.680 623.690 15.740 ;
      LAYER via ;
        RECT 535.080 15.680 535.340 15.940 ;
        RECT 623.400 15.680 623.660 15.940 ;
      LAYER met2 ;
        RECT 390.990 400.180 391.270 404.000 ;
        RECT 390.990 400.000 391.300 400.180 ;
        RECT 391.160 389.485 391.300 400.000 ;
        RECT 391.090 389.115 391.370 389.485 ;
        RECT 534.150 389.115 534.430 389.485 ;
        RECT 534.220 372.670 534.360 389.115 ;
        RECT 534.220 372.530 534.820 372.670 ;
        RECT 534.680 82.870 534.820 372.530 ;
        RECT 534.680 82.730 535.280 82.870 ;
        RECT 535.140 15.970 535.280 82.730 ;
        RECT 535.080 15.650 535.340 15.970 ;
        RECT 623.400 15.650 623.660 15.970 ;
        RECT 623.460 2.400 623.600 15.650 ;
        RECT 623.250 -4.800 623.810 2.400 ;
      LAYER via2 ;
        RECT 391.090 389.160 391.370 389.440 ;
        RECT 534.150 389.160 534.430 389.440 ;
      LAYER met3 ;
        RECT 391.065 389.450 391.395 389.465 ;
        RECT 534.125 389.450 534.455 389.465 ;
        RECT 391.065 389.150 534.455 389.450 ;
        RECT 391.065 389.135 391.395 389.150 ;
        RECT 534.125 389.135 534.455 389.150 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 117.370 391.920 117.690 391.980 ;
        RECT 236.510 391.920 236.830 391.980 ;
        RECT 117.370 391.780 236.830 391.920 ;
        RECT 117.370 391.720 117.690 391.780 ;
        RECT 236.510 391.720 236.830 391.780 ;
      LAYER via ;
        RECT 117.400 391.720 117.660 391.980 ;
        RECT 236.540 391.720 236.800 391.980 ;
      LAYER met2 ;
        RECT 236.430 400.180 236.710 404.000 ;
        RECT 236.430 400.000 236.740 400.180 ;
        RECT 236.600 392.010 236.740 400.000 ;
        RECT 117.400 391.690 117.660 392.010 ;
        RECT 236.540 391.690 236.800 392.010 ;
        RECT 117.460 82.870 117.600 391.690 ;
        RECT 117.460 82.730 121.280 82.870 ;
        RECT 121.140 2.400 121.280 82.730 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 144.510 16.560 144.830 16.620 ;
        RECT 242.030 16.560 242.350 16.620 ;
        RECT 144.510 16.420 242.350 16.560 ;
        RECT 144.510 16.360 144.830 16.420 ;
        RECT 242.030 16.360 242.350 16.420 ;
      LAYER via ;
        RECT 144.540 16.360 144.800 16.620 ;
        RECT 242.060 16.360 242.320 16.620 ;
      LAYER met2 ;
        RECT 243.790 400.250 244.070 404.000 ;
        RECT 242.580 400.110 244.070 400.250 ;
        RECT 242.580 386.650 242.720 400.110 ;
        RECT 243.790 400.000 244.070 400.110 ;
        RECT 242.120 386.510 242.720 386.650 ;
        RECT 242.120 16.650 242.260 386.510 ;
        RECT 144.540 16.330 144.800 16.650 ;
        RECT 242.060 16.330 242.320 16.650 ;
        RECT 144.600 2.400 144.740 16.330 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.770 392.260 159.090 392.320 ;
        RECT 249.390 392.260 249.710 392.320 ;
        RECT 158.770 392.120 249.710 392.260 ;
        RECT 158.770 392.060 159.090 392.120 ;
        RECT 249.390 392.060 249.710 392.120 ;
      LAYER via ;
        RECT 158.800 392.060 159.060 392.320 ;
        RECT 249.420 392.060 249.680 392.320 ;
      LAYER met2 ;
        RECT 249.310 400.180 249.590 404.000 ;
        RECT 249.310 400.000 249.620 400.180 ;
        RECT 249.480 392.350 249.620 400.000 ;
        RECT 158.800 392.030 159.060 392.350 ;
        RECT 249.420 392.030 249.680 392.350 ;
        RECT 158.860 82.870 159.000 392.030 ;
        RECT 158.860 82.730 159.920 82.870 ;
        RECT 159.780 1.770 159.920 82.730 ;
        RECT 161.870 1.770 162.430 2.400 ;
        RECT 159.780 1.630 162.430 1.770 ;
        RECT 161.870 -4.800 162.430 1.630 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 249.390 386.140 249.710 386.200 ;
        RECT 253.530 386.140 253.850 386.200 ;
        RECT 249.390 386.000 253.850 386.140 ;
        RECT 249.390 385.940 249.710 386.000 ;
        RECT 253.530 385.940 253.850 386.000 ;
        RECT 231.910 17.920 232.230 17.980 ;
        RECT 249.390 17.920 249.710 17.980 ;
        RECT 231.910 17.780 249.710 17.920 ;
        RECT 231.910 17.720 232.230 17.780 ;
        RECT 249.390 17.720 249.710 17.780 ;
        RECT 179.930 15.540 180.250 15.600 ;
        RECT 231.910 15.540 232.230 15.600 ;
        RECT 179.930 15.400 232.230 15.540 ;
        RECT 179.930 15.340 180.250 15.400 ;
        RECT 231.910 15.340 232.230 15.400 ;
      LAYER via ;
        RECT 249.420 385.940 249.680 386.200 ;
        RECT 253.560 385.940 253.820 386.200 ;
        RECT 231.940 17.720 232.200 17.980 ;
        RECT 249.420 17.720 249.680 17.980 ;
        RECT 179.960 15.340 180.220 15.600 ;
        RECT 231.940 15.340 232.200 15.600 ;
      LAYER met2 ;
        RECT 254.830 400.250 255.110 404.000 ;
        RECT 253.620 400.110 255.110 400.250 ;
        RECT 253.620 386.230 253.760 400.110 ;
        RECT 254.830 400.000 255.110 400.110 ;
        RECT 249.420 385.910 249.680 386.230 ;
        RECT 253.560 385.910 253.820 386.230 ;
        RECT 249.480 18.010 249.620 385.910 ;
        RECT 231.940 17.690 232.200 18.010 ;
        RECT 249.420 17.690 249.680 18.010 ;
        RECT 232.000 15.630 232.140 17.690 ;
        RECT 179.960 15.310 180.220 15.630 ;
        RECT 231.940 15.310 232.200 15.630 ;
        RECT 180.020 2.400 180.160 15.310 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 193.270 388.860 193.590 388.920 ;
        RECT 260.430 388.860 260.750 388.920 ;
        RECT 193.270 388.720 260.750 388.860 ;
        RECT 193.270 388.660 193.590 388.720 ;
        RECT 260.430 388.660 260.750 388.720 ;
      LAYER via ;
        RECT 193.300 388.660 193.560 388.920 ;
        RECT 260.460 388.660 260.720 388.920 ;
      LAYER met2 ;
        RECT 260.350 400.180 260.630 404.000 ;
        RECT 260.350 400.000 260.660 400.180 ;
        RECT 260.520 388.950 260.660 400.000 ;
        RECT 193.300 388.630 193.560 388.950 ;
        RECT 260.460 388.630 260.720 388.950 ;
        RECT 193.360 82.870 193.500 388.630 ;
        RECT 193.360 82.730 195.800 82.870 ;
        RECT 195.660 1.770 195.800 82.730 ;
        RECT 197.750 1.770 198.310 2.400 ;
        RECT 195.660 1.630 198.310 1.770 ;
        RECT 197.750 -4.800 198.310 1.630 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 224.090 390.220 224.410 390.280 ;
        RECT 265.950 390.220 266.270 390.280 ;
        RECT 224.090 390.080 266.270 390.220 ;
        RECT 224.090 390.020 224.410 390.080 ;
        RECT 265.950 390.020 266.270 390.080 ;
        RECT 215.350 17.580 215.670 17.640 ;
        RECT 224.090 17.580 224.410 17.640 ;
        RECT 215.350 17.440 224.410 17.580 ;
        RECT 215.350 17.380 215.670 17.440 ;
        RECT 224.090 17.380 224.410 17.440 ;
      LAYER via ;
        RECT 224.120 390.020 224.380 390.280 ;
        RECT 265.980 390.020 266.240 390.280 ;
        RECT 215.380 17.380 215.640 17.640 ;
        RECT 224.120 17.380 224.380 17.640 ;
      LAYER met2 ;
        RECT 265.870 400.180 266.150 404.000 ;
        RECT 265.870 400.000 266.180 400.180 ;
        RECT 266.040 390.310 266.180 400.000 ;
        RECT 224.120 389.990 224.380 390.310 ;
        RECT 265.980 389.990 266.240 390.310 ;
        RECT 224.180 17.670 224.320 389.990 ;
        RECT 215.380 17.350 215.640 17.670 ;
        RECT 224.120 17.350 224.380 17.670 ;
        RECT 215.440 2.400 215.580 17.350 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 252.150 387.500 252.470 387.560 ;
        RECT 271.010 387.500 271.330 387.560 ;
        RECT 252.150 387.360 271.330 387.500 ;
        RECT 252.150 387.300 252.470 387.360 ;
        RECT 271.010 387.300 271.330 387.360 ;
        RECT 233.290 16.220 233.610 16.280 ;
        RECT 251.690 16.220 252.010 16.280 ;
        RECT 233.290 16.080 252.010 16.220 ;
        RECT 233.290 16.020 233.610 16.080 ;
        RECT 251.690 16.020 252.010 16.080 ;
      LAYER via ;
        RECT 252.180 387.300 252.440 387.560 ;
        RECT 271.040 387.300 271.300 387.560 ;
        RECT 233.320 16.020 233.580 16.280 ;
        RECT 251.720 16.020 251.980 16.280 ;
      LAYER met2 ;
        RECT 270.930 400.180 271.210 404.000 ;
        RECT 270.930 400.000 271.240 400.180 ;
        RECT 271.100 387.590 271.240 400.000 ;
        RECT 252.180 387.270 252.440 387.590 ;
        RECT 271.040 387.270 271.300 387.590 ;
        RECT 252.240 324.370 252.380 387.270 ;
        RECT 251.780 324.230 252.380 324.370 ;
        RECT 251.780 16.310 251.920 324.230 ;
        RECT 233.320 15.990 233.580 16.310 ;
        RECT 251.720 15.990 251.980 16.310 ;
        RECT 233.380 2.400 233.520 15.990 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 55.730 18.940 56.050 19.000 ;
        RECT 214.890 18.940 215.210 19.000 ;
        RECT 55.730 18.800 215.210 18.940 ;
        RECT 55.730 18.740 56.050 18.800 ;
        RECT 214.890 18.740 215.210 18.800 ;
      LAYER via ;
        RECT 55.760 18.740 56.020 19.000 ;
        RECT 214.920 18.740 215.180 19.000 ;
      LAYER met2 ;
        RECT 216.650 400.250 216.930 404.000 ;
        RECT 215.440 400.110 216.930 400.250 ;
        RECT 215.440 382.570 215.580 400.110 ;
        RECT 216.650 400.000 216.930 400.110 ;
        RECT 214.980 382.430 215.580 382.570 ;
        RECT 214.980 19.030 215.120 382.430 ;
        RECT 55.760 18.710 56.020 19.030 ;
        RECT 214.920 18.710 215.180 19.030 ;
        RECT 55.820 2.400 55.960 18.710 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 75.970 391.580 76.290 391.640 ;
        RECT 224.090 391.580 224.410 391.640 ;
        RECT 75.970 391.440 224.410 391.580 ;
        RECT 75.970 391.380 76.290 391.440 ;
        RECT 224.090 391.380 224.410 391.440 ;
      LAYER via ;
        RECT 76.000 391.380 76.260 391.640 ;
        RECT 224.120 391.380 224.380 391.640 ;
      LAYER met2 ;
        RECT 224.010 400.180 224.290 404.000 ;
        RECT 224.010 400.000 224.320 400.180 ;
        RECT 224.180 391.670 224.320 400.000 ;
        RECT 76.000 391.350 76.260 391.670 ;
        RECT 224.120 391.350 224.380 391.670 ;
        RECT 76.060 82.870 76.200 391.350 ;
        RECT 76.060 82.730 79.880 82.870 ;
        RECT 79.740 2.400 79.880 82.730 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.230 386.480 228.550 386.540 ;
        RECT 230.070 386.480 230.390 386.540 ;
        RECT 228.230 386.340 230.390 386.480 ;
        RECT 228.230 386.280 228.550 386.340 ;
        RECT 230.070 386.280 230.390 386.340 ;
        RECT 103.110 20.640 103.430 20.700 ;
        RECT 228.230 20.640 228.550 20.700 ;
        RECT 103.110 20.500 228.550 20.640 ;
        RECT 103.110 20.440 103.430 20.500 ;
        RECT 228.230 20.440 228.550 20.500 ;
      LAYER via ;
        RECT 228.260 386.280 228.520 386.540 ;
        RECT 230.100 386.280 230.360 386.540 ;
        RECT 103.140 20.440 103.400 20.700 ;
        RECT 228.260 20.440 228.520 20.700 ;
      LAYER met2 ;
        RECT 231.370 400.250 231.650 404.000 ;
        RECT 230.160 400.110 231.650 400.250 ;
        RECT 230.160 386.570 230.300 400.110 ;
        RECT 231.370 400.000 231.650 400.110 ;
        RECT 228.260 386.250 228.520 386.570 ;
        RECT 230.100 386.250 230.360 386.570 ;
        RECT 228.320 20.730 228.460 386.250 ;
        RECT 103.140 20.410 103.400 20.730 ;
        RECT 228.260 20.410 228.520 20.730 ;
        RECT 103.200 2.400 103.340 20.410 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 124.270 392.600 124.590 392.660 ;
        RECT 238.350 392.600 238.670 392.660 ;
        RECT 124.270 392.460 238.670 392.600 ;
        RECT 124.270 392.400 124.590 392.460 ;
        RECT 238.350 392.400 238.670 392.460 ;
      LAYER via ;
        RECT 124.300 392.400 124.560 392.660 ;
        RECT 238.380 392.400 238.640 392.660 ;
      LAYER met2 ;
        RECT 238.270 400.180 238.550 404.000 ;
        RECT 238.270 400.000 238.580 400.180 ;
        RECT 238.440 392.690 238.580 400.000 ;
        RECT 124.300 392.370 124.560 392.690 ;
        RECT 238.380 392.370 238.640 392.690 ;
        RECT 124.360 82.870 124.500 392.370 ;
        RECT 124.360 82.730 126.800 82.870 ;
        RECT 126.660 2.400 126.800 82.730 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 207.530 17.240 207.850 17.300 ;
        RECT 26.290 17.100 207.850 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 207.530 17.040 207.850 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 207.560 17.040 207.820 17.300 ;
      LAYER met2 ;
        RECT 207.450 400.180 207.730 404.000 ;
        RECT 207.450 400.000 207.760 400.180 ;
        RECT 207.620 17.330 207.760 400.000 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 207.560 17.010 207.820 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.670 390.220 27.990 390.280 ;
        RECT 209.370 390.220 209.690 390.280 ;
        RECT 27.670 390.080 209.690 390.220 ;
        RECT 27.670 390.020 27.990 390.080 ;
        RECT 209.370 390.020 209.690 390.080 ;
      LAYER via ;
        RECT 27.700 390.020 27.960 390.280 ;
        RECT 209.400 390.020 209.660 390.280 ;
      LAYER met2 ;
        RECT 209.290 400.180 209.570 404.000 ;
        RECT 209.290 400.000 209.600 400.180 ;
        RECT 209.460 390.310 209.600 400.000 ;
        RECT 27.700 389.990 27.960 390.310 ;
        RECT 209.400 389.990 209.660 390.310 ;
        RECT 27.760 82.870 27.900 389.990 ;
        RECT 27.760 82.730 30.200 82.870 ;
        RECT 30.060 1.770 30.200 82.730 ;
        RECT 32.150 1.770 32.710 2.400 ;
        RECT 30.060 1.630 32.710 1.770 ;
        RECT 32.150 -4.800 32.710 1.630 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 205.520 410.795 1094.240 987.605 ;
      LAYER met1 ;
        RECT 203.750 410.640 1094.240 991.900 ;
      LAYER met2 ;
        RECT 204.330 995.720 210.850 996.770 ;
        RECT 211.690 995.720 218.210 996.770 ;
        RECT 219.050 995.720 225.570 996.770 ;
        RECT 226.410 995.720 232.930 996.770 ;
        RECT 233.770 995.720 240.290 996.770 ;
        RECT 241.130 995.720 248.110 996.770 ;
        RECT 248.950 995.720 255.470 996.770 ;
        RECT 256.310 995.720 262.830 996.770 ;
        RECT 263.670 995.720 270.190 996.770 ;
        RECT 271.030 995.720 277.550 996.770 ;
        RECT 278.390 995.720 284.910 996.770 ;
        RECT 285.750 995.720 292.730 996.770 ;
        RECT 293.570 995.720 300.090 996.770 ;
        RECT 300.930 995.720 307.450 996.770 ;
        RECT 308.290 995.720 314.810 996.770 ;
        RECT 315.650 995.720 322.170 996.770 ;
        RECT 323.010 995.720 329.530 996.770 ;
        RECT 330.370 995.720 337.350 996.770 ;
        RECT 338.190 995.720 344.710 996.770 ;
        RECT 345.550 995.720 352.070 996.770 ;
        RECT 352.910 995.720 359.430 996.770 ;
        RECT 360.270 995.720 366.790 996.770 ;
        RECT 367.630 995.720 374.150 996.770 ;
        RECT 374.990 995.720 381.970 996.770 ;
        RECT 382.810 995.720 389.330 996.770 ;
        RECT 390.170 995.720 396.690 996.770 ;
        RECT 397.530 995.720 404.050 996.770 ;
        RECT 404.890 995.720 411.410 996.770 ;
        RECT 412.250 995.720 419.230 996.770 ;
        RECT 420.070 995.720 426.590 996.770 ;
        RECT 427.430 995.720 433.950 996.770 ;
        RECT 434.790 995.720 441.310 996.770 ;
        RECT 442.150 995.720 448.670 996.770 ;
        RECT 449.510 995.720 456.030 996.770 ;
        RECT 456.870 995.720 463.850 996.770 ;
        RECT 464.690 995.720 471.210 996.770 ;
        RECT 472.050 995.720 478.570 996.770 ;
        RECT 479.410 995.720 485.930 996.770 ;
        RECT 486.770 995.720 493.290 996.770 ;
        RECT 494.130 995.720 500.650 996.770 ;
        RECT 501.490 995.720 508.470 996.770 ;
        RECT 509.310 995.720 515.830 996.770 ;
        RECT 516.670 995.720 523.190 996.770 ;
        RECT 524.030 995.720 530.550 996.770 ;
        RECT 531.390 995.720 537.910 996.770 ;
        RECT 538.750 995.720 545.270 996.770 ;
        RECT 546.110 995.720 553.090 996.770 ;
        RECT 553.930 995.720 560.450 996.770 ;
        RECT 561.290 995.720 567.810 996.770 ;
        RECT 568.650 995.720 575.170 996.770 ;
        RECT 576.010 995.720 582.530 996.770 ;
        RECT 583.370 995.720 590.350 996.770 ;
        RECT 591.190 995.720 597.710 996.770 ;
        RECT 598.550 995.720 605.070 996.770 ;
        RECT 605.910 995.720 612.430 996.770 ;
        RECT 613.270 995.720 619.790 996.770 ;
        RECT 620.630 995.720 627.150 996.770 ;
        RECT 627.990 995.720 634.970 996.770 ;
        RECT 635.810 995.720 642.330 996.770 ;
        RECT 643.170 995.720 649.690 996.770 ;
        RECT 650.530 995.720 657.050 996.770 ;
        RECT 657.890 995.720 664.410 996.770 ;
        RECT 665.250 995.720 671.770 996.770 ;
        RECT 672.610 995.720 679.590 996.770 ;
        RECT 680.430 995.720 686.950 996.770 ;
        RECT 687.790 995.720 694.310 996.770 ;
        RECT 695.150 995.720 701.670 996.770 ;
        RECT 702.510 995.720 709.030 996.770 ;
        RECT 709.870 995.720 716.390 996.770 ;
        RECT 717.230 995.720 724.210 996.770 ;
        RECT 725.050 995.720 731.570 996.770 ;
        RECT 732.410 995.720 738.930 996.770 ;
        RECT 739.770 995.720 746.290 996.770 ;
        RECT 747.130 995.720 753.650 996.770 ;
        RECT 754.490 995.720 761.470 996.770 ;
        RECT 762.310 995.720 768.830 996.770 ;
        RECT 769.670 995.720 776.190 996.770 ;
        RECT 777.030 995.720 783.550 996.770 ;
        RECT 784.390 995.720 790.910 996.770 ;
        RECT 791.750 995.720 798.270 996.770 ;
        RECT 799.110 995.720 806.090 996.770 ;
        RECT 806.930 995.720 813.450 996.770 ;
        RECT 814.290 995.720 820.810 996.770 ;
        RECT 821.650 995.720 828.170 996.770 ;
        RECT 829.010 995.720 835.530 996.770 ;
        RECT 836.370 995.720 842.890 996.770 ;
        RECT 843.730 995.720 850.710 996.770 ;
        RECT 851.550 995.720 858.070 996.770 ;
        RECT 858.910 995.720 865.430 996.770 ;
        RECT 866.270 995.720 872.790 996.770 ;
        RECT 873.630 995.720 880.150 996.770 ;
        RECT 880.990 995.720 887.510 996.770 ;
        RECT 888.350 995.720 895.330 996.770 ;
        RECT 896.170 995.720 902.690 996.770 ;
        RECT 903.530 995.720 910.050 996.770 ;
        RECT 910.890 995.720 917.410 996.770 ;
        RECT 918.250 995.720 924.770 996.770 ;
        RECT 925.610 995.720 932.590 996.770 ;
        RECT 933.430 995.720 939.950 996.770 ;
        RECT 940.790 995.720 947.310 996.770 ;
        RECT 948.150 995.720 954.670 996.770 ;
        RECT 955.510 995.720 962.030 996.770 ;
        RECT 962.870 995.720 969.390 996.770 ;
        RECT 970.230 995.720 977.210 996.770 ;
        RECT 978.050 995.720 984.570 996.770 ;
        RECT 985.410 995.720 991.930 996.770 ;
        RECT 992.770 995.720 999.290 996.770 ;
        RECT 1000.130 995.720 1006.650 996.770 ;
        RECT 1007.490 995.720 1014.010 996.770 ;
        RECT 1014.850 995.720 1021.830 996.770 ;
        RECT 1022.670 995.720 1029.190 996.770 ;
        RECT 1030.030 995.720 1036.550 996.770 ;
        RECT 1037.390 995.720 1043.910 996.770 ;
        RECT 1044.750 995.720 1051.270 996.770 ;
        RECT 1052.110 995.720 1058.630 996.770 ;
        RECT 1059.470 995.720 1066.450 996.770 ;
        RECT 1067.290 995.720 1073.810 996.770 ;
        RECT 1074.650 995.720 1081.170 996.770 ;
        RECT 1082.010 995.720 1088.530 996.770 ;
        RECT 1089.370 995.720 1091.840 996.770 ;
        RECT 203.780 404.280 1091.840 995.720 ;
      LAYER met2 ;
        RECT 200.550 400.000 200.830 404.000 ;
      LAYER met2 ;
        RECT 204.330 403.670 205.330 404.280 ;
        RECT 206.170 403.670 207.170 404.280 ;
        RECT 208.010 403.670 209.010 404.280 ;
        RECT 209.850 403.670 210.850 404.280 ;
        RECT 211.690 403.670 212.690 404.280 ;
        RECT 213.530 403.670 214.530 404.280 ;
        RECT 215.370 403.670 216.370 404.280 ;
        RECT 217.210 403.670 218.210 404.280 ;
        RECT 219.050 403.670 220.050 404.280 ;
        RECT 220.890 403.670 221.890 404.280 ;
        RECT 222.730 403.670 223.730 404.280 ;
        RECT 224.570 403.670 225.570 404.280 ;
        RECT 226.410 403.670 227.410 404.280 ;
        RECT 228.250 403.670 229.250 404.280 ;
        RECT 230.090 403.670 231.090 404.280 ;
        RECT 231.930 403.670 232.930 404.280 ;
        RECT 233.770 403.670 234.310 404.280 ;
        RECT 235.150 403.670 236.150 404.280 ;
        RECT 236.990 403.670 237.990 404.280 ;
        RECT 238.830 403.670 239.830 404.280 ;
        RECT 240.670 403.670 241.670 404.280 ;
        RECT 242.510 403.670 243.510 404.280 ;
        RECT 244.350 403.670 245.350 404.280 ;
        RECT 246.190 403.670 247.190 404.280 ;
        RECT 248.030 403.670 249.030 404.280 ;
        RECT 249.870 403.670 250.870 404.280 ;
        RECT 251.710 403.670 252.710 404.280 ;
        RECT 253.550 403.670 254.550 404.280 ;
        RECT 255.390 403.670 256.390 404.280 ;
        RECT 257.230 403.670 258.230 404.280 ;
        RECT 259.070 403.670 260.070 404.280 ;
        RECT 260.910 403.670 261.910 404.280 ;
        RECT 262.750 403.670 263.750 404.280 ;
        RECT 264.590 403.670 265.590 404.280 ;
        RECT 266.430 403.670 266.970 404.280 ;
        RECT 267.810 403.670 268.810 404.280 ;
        RECT 269.650 403.670 270.650 404.280 ;
        RECT 271.490 403.670 272.490 404.280 ;
        RECT 273.330 403.670 274.330 404.280 ;
        RECT 275.170 403.670 276.170 404.280 ;
        RECT 277.010 403.670 278.010 404.280 ;
        RECT 278.850 403.670 279.850 404.280 ;
        RECT 280.690 403.670 281.690 404.280 ;
        RECT 282.530 403.670 283.530 404.280 ;
        RECT 284.370 403.670 285.370 404.280 ;
        RECT 286.210 403.670 287.210 404.280 ;
        RECT 288.050 403.670 289.050 404.280 ;
        RECT 289.890 403.670 290.890 404.280 ;
        RECT 291.730 403.670 292.730 404.280 ;
        RECT 293.570 403.670 294.570 404.280 ;
        RECT 295.410 403.670 296.410 404.280 ;
        RECT 297.250 403.670 298.250 404.280 ;
        RECT 299.090 403.670 300.090 404.280 ;
        RECT 300.930 403.670 301.470 404.280 ;
        RECT 302.310 403.670 303.310 404.280 ;
        RECT 304.150 403.670 305.150 404.280 ;
        RECT 305.990 403.670 306.990 404.280 ;
        RECT 307.830 403.670 308.830 404.280 ;
        RECT 309.670 403.670 310.670 404.280 ;
        RECT 311.510 403.670 312.510 404.280 ;
        RECT 313.350 403.670 314.350 404.280 ;
        RECT 315.190 403.670 316.190 404.280 ;
        RECT 317.030 403.670 318.030 404.280 ;
        RECT 318.870 403.670 319.870 404.280 ;
        RECT 320.710 403.670 321.710 404.280 ;
        RECT 322.550 403.670 323.550 404.280 ;
        RECT 324.390 403.670 325.390 404.280 ;
        RECT 326.230 403.670 327.230 404.280 ;
        RECT 328.070 403.670 329.070 404.280 ;
        RECT 329.910 403.670 330.910 404.280 ;
        RECT 331.750 403.670 332.750 404.280 ;
        RECT 333.590 403.670 334.130 404.280 ;
        RECT 334.970 403.670 335.970 404.280 ;
        RECT 336.810 403.670 337.810 404.280 ;
        RECT 338.650 403.670 339.650 404.280 ;
        RECT 340.490 403.670 341.490 404.280 ;
        RECT 342.330 403.670 343.330 404.280 ;
        RECT 344.170 403.670 345.170 404.280 ;
        RECT 346.010 403.670 347.010 404.280 ;
        RECT 347.850 403.670 348.850 404.280 ;
        RECT 349.690 403.670 350.690 404.280 ;
        RECT 351.530 403.670 352.530 404.280 ;
        RECT 353.370 403.670 354.370 404.280 ;
        RECT 355.210 403.670 356.210 404.280 ;
        RECT 357.050 403.670 358.050 404.280 ;
        RECT 358.890 403.670 359.890 404.280 ;
        RECT 360.730 403.670 361.730 404.280 ;
        RECT 362.570 403.670 363.570 404.280 ;
        RECT 364.410 403.670 365.410 404.280 ;
        RECT 366.250 403.670 366.790 404.280 ;
        RECT 367.630 403.670 368.630 404.280 ;
        RECT 369.470 403.670 370.470 404.280 ;
        RECT 371.310 403.670 372.310 404.280 ;
        RECT 373.150 403.670 374.150 404.280 ;
        RECT 374.990 403.670 375.990 404.280 ;
        RECT 376.830 403.670 377.830 404.280 ;
        RECT 378.670 403.670 379.670 404.280 ;
        RECT 380.510 403.670 381.510 404.280 ;
        RECT 382.350 403.670 383.350 404.280 ;
        RECT 384.190 403.670 385.190 404.280 ;
        RECT 386.030 403.670 387.030 404.280 ;
        RECT 387.870 403.670 388.870 404.280 ;
        RECT 389.710 403.670 390.710 404.280 ;
        RECT 391.550 403.670 392.550 404.280 ;
        RECT 393.390 403.670 394.390 404.280 ;
        RECT 395.230 403.670 396.230 404.280 ;
        RECT 397.070 403.670 398.070 404.280 ;
        RECT 398.910 403.670 399.910 404.280 ;
        RECT 400.750 403.670 401.290 404.280 ;
        RECT 402.130 403.670 403.130 404.280 ;
        RECT 403.970 403.670 404.970 404.280 ;
        RECT 405.810 403.670 406.810 404.280 ;
        RECT 407.650 403.670 408.650 404.280 ;
        RECT 409.490 403.670 410.490 404.280 ;
        RECT 411.330 403.670 412.330 404.280 ;
        RECT 413.170 403.670 414.170 404.280 ;
        RECT 415.010 403.670 416.010 404.280 ;
        RECT 416.850 403.670 417.850 404.280 ;
        RECT 418.690 403.670 419.690 404.280 ;
        RECT 420.530 403.670 421.530 404.280 ;
        RECT 422.370 403.670 423.370 404.280 ;
        RECT 424.210 403.670 425.210 404.280 ;
        RECT 426.050 403.670 427.050 404.280 ;
        RECT 427.890 403.670 428.890 404.280 ;
        RECT 429.730 403.670 430.730 404.280 ;
        RECT 431.570 403.670 432.570 404.280 ;
        RECT 433.410 403.670 433.950 404.280 ;
        RECT 434.790 403.670 435.790 404.280 ;
        RECT 436.630 403.670 437.630 404.280 ;
        RECT 438.470 403.670 439.470 404.280 ;
        RECT 440.310 403.670 441.310 404.280 ;
        RECT 442.150 403.670 443.150 404.280 ;
        RECT 443.990 403.670 444.990 404.280 ;
        RECT 445.830 403.670 446.830 404.280 ;
        RECT 447.670 403.670 448.670 404.280 ;
        RECT 449.510 403.670 450.510 404.280 ;
        RECT 451.350 403.670 452.350 404.280 ;
        RECT 453.190 403.670 454.190 404.280 ;
        RECT 455.030 403.670 456.030 404.280 ;
        RECT 456.870 403.670 457.870 404.280 ;
        RECT 458.710 403.670 459.710 404.280 ;
        RECT 460.550 403.670 461.550 404.280 ;
        RECT 462.390 403.670 463.390 404.280 ;
        RECT 464.230 403.670 465.230 404.280 ;
        RECT 466.070 403.670 466.610 404.280 ;
        RECT 467.450 403.670 468.450 404.280 ;
        RECT 469.290 403.670 470.290 404.280 ;
        RECT 471.130 403.670 472.130 404.280 ;
        RECT 472.970 403.670 473.970 404.280 ;
        RECT 474.810 403.670 475.810 404.280 ;
        RECT 476.650 403.670 477.650 404.280 ;
        RECT 478.490 403.670 479.490 404.280 ;
        RECT 480.330 403.670 481.330 404.280 ;
        RECT 482.170 403.670 483.170 404.280 ;
        RECT 484.010 403.670 485.010 404.280 ;
        RECT 485.850 403.670 486.850 404.280 ;
        RECT 487.690 403.670 488.690 404.280 ;
        RECT 489.530 403.670 490.530 404.280 ;
        RECT 491.370 403.670 492.370 404.280 ;
        RECT 493.210 403.670 494.210 404.280 ;
        RECT 495.050 403.670 496.050 404.280 ;
        RECT 496.890 403.670 497.890 404.280 ;
        RECT 498.730 403.670 499.730 404.280 ;
        RECT 500.570 403.670 501.110 404.280 ;
        RECT 501.950 403.670 502.950 404.280 ;
        RECT 503.790 403.670 504.790 404.280 ;
        RECT 505.630 403.670 506.630 404.280 ;
        RECT 507.470 403.670 508.470 404.280 ;
        RECT 509.310 403.670 510.310 404.280 ;
        RECT 511.150 403.670 512.150 404.280 ;
        RECT 512.990 403.670 513.990 404.280 ;
        RECT 514.830 403.670 515.830 404.280 ;
        RECT 516.670 403.670 517.670 404.280 ;
        RECT 518.510 403.670 519.510 404.280 ;
        RECT 520.350 403.670 521.350 404.280 ;
        RECT 522.190 403.670 523.190 404.280 ;
        RECT 524.030 403.670 525.030 404.280 ;
        RECT 525.870 403.670 526.870 404.280 ;
        RECT 527.710 403.670 528.710 404.280 ;
        RECT 529.550 403.670 530.550 404.280 ;
        RECT 531.390 403.670 532.390 404.280 ;
        RECT 533.230 403.670 533.770 404.280 ;
        RECT 534.610 403.670 535.610 404.280 ;
        RECT 536.450 403.670 537.450 404.280 ;
        RECT 538.290 403.670 539.290 404.280 ;
        RECT 540.130 403.670 541.130 404.280 ;
        RECT 541.970 403.670 542.970 404.280 ;
        RECT 543.810 403.670 544.810 404.280 ;
        RECT 545.650 403.670 546.650 404.280 ;
        RECT 547.490 403.670 548.490 404.280 ;
        RECT 549.330 403.670 550.330 404.280 ;
        RECT 551.170 403.670 552.170 404.280 ;
        RECT 553.010 403.670 554.010 404.280 ;
        RECT 554.850 403.670 555.850 404.280 ;
        RECT 556.690 403.670 557.690 404.280 ;
        RECT 558.530 403.670 559.530 404.280 ;
        RECT 560.370 403.670 561.370 404.280 ;
        RECT 562.210 403.670 563.210 404.280 ;
        RECT 564.050 403.670 565.050 404.280 ;
        RECT 565.890 403.670 566.890 404.280 ;
        RECT 567.730 403.670 568.270 404.280 ;
        RECT 569.110 403.670 570.110 404.280 ;
        RECT 570.950 403.670 571.950 404.280 ;
        RECT 572.790 403.670 573.790 404.280 ;
        RECT 574.630 403.670 575.630 404.280 ;
        RECT 576.470 403.670 577.470 404.280 ;
        RECT 578.310 403.670 579.310 404.280 ;
        RECT 580.150 403.670 581.150 404.280 ;
        RECT 581.990 403.670 582.990 404.280 ;
        RECT 583.830 403.670 584.830 404.280 ;
        RECT 585.670 403.670 586.670 404.280 ;
        RECT 587.510 403.670 588.510 404.280 ;
        RECT 589.350 403.670 590.350 404.280 ;
        RECT 591.190 403.670 592.190 404.280 ;
        RECT 593.030 403.670 594.030 404.280 ;
        RECT 594.870 403.670 595.870 404.280 ;
        RECT 596.710 403.670 597.710 404.280 ;
        RECT 598.550 403.670 599.550 404.280 ;
        RECT 600.390 403.670 600.930 404.280 ;
        RECT 601.770 403.670 602.770 404.280 ;
        RECT 603.610 403.670 604.610 404.280 ;
        RECT 605.450 403.670 606.450 404.280 ;
        RECT 607.290 403.670 608.290 404.280 ;
        RECT 609.130 403.670 610.130 404.280 ;
        RECT 610.970 403.670 611.970 404.280 ;
        RECT 612.810 403.670 613.810 404.280 ;
        RECT 614.650 403.670 615.650 404.280 ;
        RECT 616.490 403.670 617.490 404.280 ;
        RECT 618.330 403.670 619.330 404.280 ;
        RECT 620.170 403.670 621.170 404.280 ;
        RECT 622.010 403.670 623.010 404.280 ;
        RECT 623.850 403.670 624.850 404.280 ;
        RECT 625.690 403.670 626.690 404.280 ;
        RECT 627.530 403.670 628.530 404.280 ;
        RECT 629.370 403.670 630.370 404.280 ;
        RECT 631.210 403.670 632.210 404.280 ;
        RECT 633.050 403.670 633.590 404.280 ;
        RECT 634.430 403.670 635.430 404.280 ;
        RECT 636.270 403.670 637.270 404.280 ;
        RECT 638.110 403.670 639.110 404.280 ;
        RECT 639.950 403.670 640.950 404.280 ;
        RECT 641.790 403.670 642.790 404.280 ;
        RECT 643.630 403.670 644.630 404.280 ;
        RECT 645.470 403.670 646.470 404.280 ;
        RECT 647.310 403.670 648.310 404.280 ;
        RECT 649.150 403.670 650.150 404.280 ;
        RECT 650.990 403.670 651.990 404.280 ;
        RECT 652.830 403.670 653.830 404.280 ;
        RECT 654.670 403.670 655.670 404.280 ;
        RECT 656.510 403.670 657.510 404.280 ;
        RECT 658.350 403.670 659.350 404.280 ;
        RECT 660.190 403.670 661.190 404.280 ;
        RECT 662.030 403.670 663.030 404.280 ;
        RECT 663.870 403.670 664.870 404.280 ;
        RECT 665.710 403.670 666.710 404.280 ;
        RECT 667.550 403.670 668.090 404.280 ;
        RECT 668.930 403.670 669.930 404.280 ;
        RECT 670.770 403.670 671.770 404.280 ;
        RECT 672.610 403.670 673.610 404.280 ;
        RECT 674.450 403.670 675.450 404.280 ;
        RECT 676.290 403.670 677.290 404.280 ;
        RECT 678.130 403.670 679.130 404.280 ;
        RECT 679.970 403.670 680.970 404.280 ;
        RECT 681.810 403.670 682.810 404.280 ;
        RECT 683.650 403.670 684.650 404.280 ;
        RECT 685.490 403.670 686.490 404.280 ;
        RECT 687.330 403.670 688.330 404.280 ;
        RECT 689.170 403.670 690.170 404.280 ;
        RECT 691.010 403.670 692.010 404.280 ;
        RECT 692.850 403.670 693.850 404.280 ;
        RECT 694.690 403.670 695.690 404.280 ;
        RECT 696.530 403.670 697.530 404.280 ;
        RECT 698.370 403.670 699.370 404.280 ;
        RECT 700.210 403.670 700.750 404.280 ;
        RECT 701.590 403.670 702.590 404.280 ;
        RECT 703.430 403.670 704.430 404.280 ;
        RECT 705.270 403.670 706.270 404.280 ;
        RECT 707.110 403.670 708.110 404.280 ;
        RECT 708.950 403.670 709.950 404.280 ;
        RECT 710.790 403.670 711.790 404.280 ;
        RECT 712.630 403.670 713.630 404.280 ;
        RECT 714.470 403.670 715.470 404.280 ;
        RECT 716.310 403.670 717.310 404.280 ;
        RECT 718.150 403.670 719.150 404.280 ;
        RECT 719.990 403.670 720.990 404.280 ;
        RECT 721.830 403.670 722.830 404.280 ;
        RECT 723.670 403.670 724.670 404.280 ;
        RECT 725.510 403.670 726.510 404.280 ;
        RECT 727.350 403.670 728.350 404.280 ;
        RECT 729.190 403.670 730.190 404.280 ;
        RECT 731.030 403.670 732.030 404.280 ;
        RECT 732.870 403.670 733.410 404.280 ;
        RECT 734.250 403.670 735.250 404.280 ;
        RECT 736.090 403.670 737.090 404.280 ;
        RECT 737.930 403.670 738.930 404.280 ;
        RECT 739.770 403.670 740.770 404.280 ;
        RECT 741.610 403.670 742.610 404.280 ;
        RECT 743.450 403.670 744.450 404.280 ;
        RECT 745.290 403.670 746.290 404.280 ;
        RECT 747.130 403.670 748.130 404.280 ;
        RECT 748.970 403.670 749.970 404.280 ;
        RECT 750.810 403.670 751.810 404.280 ;
        RECT 752.650 403.670 753.650 404.280 ;
        RECT 754.490 403.670 755.490 404.280 ;
        RECT 756.330 403.670 757.330 404.280 ;
        RECT 758.170 403.670 759.170 404.280 ;
        RECT 760.010 403.670 761.010 404.280 ;
        RECT 761.850 403.670 762.850 404.280 ;
        RECT 763.690 403.670 764.690 404.280 ;
        RECT 765.530 403.670 766.530 404.280 ;
        RECT 767.370 403.670 767.910 404.280 ;
        RECT 768.750 403.670 769.750 404.280 ;
        RECT 770.590 403.670 771.590 404.280 ;
        RECT 772.430 403.670 773.430 404.280 ;
        RECT 774.270 403.670 775.270 404.280 ;
        RECT 776.110 403.670 777.110 404.280 ;
        RECT 777.950 403.670 778.950 404.280 ;
        RECT 779.790 403.670 780.790 404.280 ;
        RECT 781.630 403.670 782.630 404.280 ;
        RECT 783.470 403.670 784.470 404.280 ;
        RECT 785.310 403.670 786.310 404.280 ;
        RECT 787.150 403.670 788.150 404.280 ;
        RECT 788.990 403.670 789.990 404.280 ;
        RECT 790.830 403.670 791.830 404.280 ;
        RECT 792.670 403.670 793.670 404.280 ;
        RECT 794.510 403.670 795.510 404.280 ;
        RECT 796.350 403.670 797.350 404.280 ;
        RECT 798.190 403.670 799.190 404.280 ;
        RECT 800.030 403.670 800.570 404.280 ;
        RECT 801.410 403.670 802.410 404.280 ;
        RECT 803.250 403.670 804.250 404.280 ;
        RECT 805.090 403.670 806.090 404.280 ;
        RECT 806.930 403.670 807.930 404.280 ;
        RECT 808.770 403.670 809.770 404.280 ;
        RECT 810.610 403.670 811.610 404.280 ;
        RECT 812.450 403.670 813.450 404.280 ;
        RECT 814.290 403.670 815.290 404.280 ;
        RECT 816.130 403.670 817.130 404.280 ;
        RECT 817.970 403.670 818.970 404.280 ;
        RECT 819.810 403.670 820.810 404.280 ;
        RECT 821.650 403.670 822.650 404.280 ;
        RECT 823.490 403.670 824.490 404.280 ;
        RECT 825.330 403.670 826.330 404.280 ;
        RECT 827.170 403.670 828.170 404.280 ;
        RECT 829.010 403.670 830.010 404.280 ;
        RECT 830.850 403.670 831.850 404.280 ;
        RECT 832.690 403.670 833.690 404.280 ;
        RECT 834.530 403.670 835.070 404.280 ;
        RECT 835.910 403.670 836.910 404.280 ;
        RECT 837.750 403.670 838.750 404.280 ;
        RECT 839.590 403.670 840.590 404.280 ;
        RECT 841.430 403.670 842.430 404.280 ;
        RECT 843.270 403.670 844.270 404.280 ;
        RECT 845.110 403.670 846.110 404.280 ;
        RECT 846.950 403.670 847.950 404.280 ;
        RECT 848.790 403.670 849.790 404.280 ;
        RECT 850.630 403.670 851.630 404.280 ;
        RECT 852.470 403.670 853.470 404.280 ;
        RECT 854.310 403.670 855.310 404.280 ;
        RECT 856.150 403.670 857.150 404.280 ;
        RECT 857.990 403.670 858.990 404.280 ;
        RECT 859.830 403.670 860.830 404.280 ;
        RECT 861.670 403.670 862.670 404.280 ;
        RECT 863.510 403.670 864.510 404.280 ;
        RECT 865.350 403.670 866.350 404.280 ;
        RECT 867.190 403.670 867.730 404.280 ;
        RECT 868.570 403.670 869.570 404.280 ;
        RECT 870.410 403.670 871.410 404.280 ;
        RECT 872.250 403.670 873.250 404.280 ;
        RECT 874.090 403.670 875.090 404.280 ;
        RECT 875.930 403.670 876.930 404.280 ;
        RECT 877.770 403.670 878.770 404.280 ;
        RECT 879.610 403.670 880.610 404.280 ;
        RECT 881.450 403.670 882.450 404.280 ;
        RECT 883.290 403.670 884.290 404.280 ;
        RECT 885.130 403.670 886.130 404.280 ;
        RECT 886.970 403.670 887.970 404.280 ;
        RECT 888.810 403.670 889.810 404.280 ;
        RECT 890.650 403.670 891.650 404.280 ;
        RECT 892.490 403.670 893.490 404.280 ;
        RECT 894.330 403.670 895.330 404.280 ;
        RECT 896.170 403.670 897.170 404.280 ;
        RECT 898.010 403.670 899.010 404.280 ;
        RECT 899.850 403.670 900.390 404.280 ;
        RECT 901.230 403.670 902.230 404.280 ;
        RECT 903.070 403.670 904.070 404.280 ;
        RECT 904.910 403.670 905.910 404.280 ;
        RECT 906.750 403.670 907.750 404.280 ;
        RECT 908.590 403.670 909.590 404.280 ;
        RECT 910.430 403.670 911.430 404.280 ;
        RECT 912.270 403.670 913.270 404.280 ;
        RECT 914.110 403.670 915.110 404.280 ;
        RECT 915.950 403.670 916.950 404.280 ;
        RECT 917.790 403.670 918.790 404.280 ;
        RECT 919.630 403.670 920.630 404.280 ;
        RECT 921.470 403.670 922.470 404.280 ;
        RECT 923.310 403.670 924.310 404.280 ;
        RECT 925.150 403.670 926.150 404.280 ;
        RECT 926.990 403.670 927.990 404.280 ;
        RECT 928.830 403.670 929.830 404.280 ;
        RECT 930.670 403.670 931.670 404.280 ;
        RECT 932.510 403.670 933.510 404.280 ;
        RECT 934.350 403.670 934.890 404.280 ;
        RECT 935.730 403.670 936.730 404.280 ;
        RECT 937.570 403.670 938.570 404.280 ;
        RECT 939.410 403.670 940.410 404.280 ;
        RECT 941.250 403.670 942.250 404.280 ;
        RECT 943.090 403.670 944.090 404.280 ;
        RECT 944.930 403.670 945.930 404.280 ;
        RECT 946.770 403.670 947.770 404.280 ;
        RECT 948.610 403.670 949.610 404.280 ;
        RECT 950.450 403.670 951.450 404.280 ;
        RECT 952.290 403.670 953.290 404.280 ;
        RECT 954.130 403.670 955.130 404.280 ;
        RECT 955.970 403.670 956.970 404.280 ;
        RECT 957.810 403.670 958.810 404.280 ;
        RECT 959.650 403.670 960.650 404.280 ;
        RECT 961.490 403.670 962.490 404.280 ;
        RECT 963.330 403.670 964.330 404.280 ;
        RECT 965.170 403.670 966.170 404.280 ;
        RECT 967.010 403.670 967.550 404.280 ;
        RECT 968.390 403.670 969.390 404.280 ;
        RECT 970.230 403.670 971.230 404.280 ;
        RECT 972.070 403.670 973.070 404.280 ;
        RECT 973.910 403.670 974.910 404.280 ;
        RECT 975.750 403.670 976.750 404.280 ;
        RECT 977.590 403.670 978.590 404.280 ;
        RECT 979.430 403.670 980.430 404.280 ;
        RECT 981.270 403.670 982.270 404.280 ;
        RECT 983.110 403.670 984.110 404.280 ;
        RECT 984.950 403.670 985.950 404.280 ;
        RECT 986.790 403.670 987.790 404.280 ;
        RECT 988.630 403.670 989.630 404.280 ;
        RECT 990.470 403.670 991.470 404.280 ;
        RECT 992.310 403.670 993.310 404.280 ;
        RECT 994.150 403.670 995.150 404.280 ;
        RECT 995.990 403.670 996.990 404.280 ;
        RECT 997.830 403.670 998.830 404.280 ;
        RECT 999.670 403.670 1000.210 404.280 ;
        RECT 1001.050 403.670 1002.050 404.280 ;
        RECT 1002.890 403.670 1003.890 404.280 ;
        RECT 1004.730 403.670 1005.730 404.280 ;
        RECT 1006.570 403.670 1007.570 404.280 ;
        RECT 1008.410 403.670 1009.410 404.280 ;
        RECT 1010.250 403.670 1011.250 404.280 ;
        RECT 1012.090 403.670 1013.090 404.280 ;
        RECT 1013.930 403.670 1014.930 404.280 ;
        RECT 1015.770 403.670 1016.770 404.280 ;
        RECT 1017.610 403.670 1018.610 404.280 ;
        RECT 1019.450 403.670 1020.450 404.280 ;
        RECT 1021.290 403.670 1022.290 404.280 ;
        RECT 1023.130 403.670 1024.130 404.280 ;
        RECT 1024.970 403.670 1025.970 404.280 ;
        RECT 1026.810 403.670 1027.810 404.280 ;
        RECT 1028.650 403.670 1029.650 404.280 ;
        RECT 1030.490 403.670 1031.490 404.280 ;
        RECT 1032.330 403.670 1033.330 404.280 ;
        RECT 1034.170 403.670 1034.710 404.280 ;
        RECT 1035.550 403.670 1036.550 404.280 ;
        RECT 1037.390 403.670 1038.390 404.280 ;
        RECT 1039.230 403.670 1040.230 404.280 ;
        RECT 1041.070 403.670 1042.070 404.280 ;
        RECT 1042.910 403.670 1043.910 404.280 ;
        RECT 1044.750 403.670 1045.750 404.280 ;
        RECT 1046.590 403.670 1047.590 404.280 ;
        RECT 1048.430 403.670 1049.430 404.280 ;
        RECT 1050.270 403.670 1051.270 404.280 ;
        RECT 1052.110 403.670 1053.110 404.280 ;
        RECT 1053.950 403.670 1054.950 404.280 ;
        RECT 1055.790 403.670 1056.790 404.280 ;
        RECT 1057.630 403.670 1058.630 404.280 ;
        RECT 1059.470 403.670 1060.470 404.280 ;
        RECT 1061.310 403.670 1062.310 404.280 ;
        RECT 1063.150 403.670 1064.150 404.280 ;
        RECT 1064.990 403.670 1065.990 404.280 ;
        RECT 1066.830 403.670 1067.370 404.280 ;
        RECT 1068.210 403.670 1069.210 404.280 ;
        RECT 1070.050 403.670 1071.050 404.280 ;
        RECT 1071.890 403.670 1072.890 404.280 ;
        RECT 1073.730 403.670 1074.730 404.280 ;
        RECT 1075.570 403.670 1076.570 404.280 ;
        RECT 1077.410 403.670 1078.410 404.280 ;
        RECT 1079.250 403.670 1080.250 404.280 ;
        RECT 1081.090 403.670 1082.090 404.280 ;
        RECT 1082.930 403.670 1083.930 404.280 ;
        RECT 1084.770 403.670 1085.770 404.280 ;
        RECT 1086.610 403.670 1087.610 404.280 ;
        RECT 1088.450 403.670 1089.450 404.280 ;
        RECT 1090.290 403.670 1091.290 404.280 ;
      LAYER met3 ;
        RECT 208.345 979.040 1096.000 990.745 ;
        RECT 208.345 977.640 1095.600 979.040 ;
        RECT 208.345 936.200 1096.000 977.640 ;
        RECT 208.345 934.800 1095.600 936.200 ;
        RECT 208.345 893.360 1096.000 934.800 ;
        RECT 208.345 891.960 1095.600 893.360 ;
        RECT 208.345 850.520 1096.000 891.960 ;
        RECT 208.345 849.120 1095.600 850.520 ;
        RECT 208.345 807.680 1096.000 849.120 ;
        RECT 208.345 806.280 1095.600 807.680 ;
        RECT 208.345 764.840 1096.000 806.280 ;
        RECT 208.345 763.440 1095.600 764.840 ;
        RECT 208.345 722.000 1096.000 763.440 ;
        RECT 208.345 720.600 1095.600 722.000 ;
        RECT 208.345 679.160 1096.000 720.600 ;
        RECT 208.345 677.760 1095.600 679.160 ;
        RECT 208.345 636.320 1096.000 677.760 ;
        RECT 208.345 634.920 1095.600 636.320 ;
        RECT 208.345 593.480 1096.000 634.920 ;
        RECT 208.345 592.080 1095.600 593.480 ;
        RECT 208.345 550.640 1096.000 592.080 ;
        RECT 208.345 549.240 1095.600 550.640 ;
        RECT 208.345 507.800 1096.000 549.240 ;
        RECT 208.345 506.400 1095.600 507.800 ;
        RECT 208.345 464.960 1096.000 506.400 ;
        RECT 208.345 463.560 1095.600 464.960 ;
        RECT 208.345 422.120 1096.000 463.560 ;
        RECT 208.345 420.720 1095.600 422.120 ;
        RECT 208.345 410.715 1096.000 420.720 ;
      LAYER met4 ;
        RECT 537.935 988.160 684.545 990.065 ;
        RECT 537.935 951.655 604.640 988.160 ;
        RECT 607.040 951.655 681.440 988.160 ;
        RECT 683.840 951.655 684.545 988.160 ;
  END
END user_project_wrapper
END LIBRARY

